module picorv32(clk, resetn, trap, mem_valid, mem_instr, mem_ready, mem_addr, mem_wdata, mem_wstrb, mem_rdata, mem_la_read, mem_la_write, mem_la_addr, mem_la_wdata, mem_la_wstrb, pcpi_valid, pcpi_insn, pcpi_rs1, pcpi_rs2, pcpi_wr, pcpi_rd
, pcpi_wait, pcpi_ready, irq, eoi, trace_valid, trace_data);
  wire _00000_;
  wire _00001_;
  wire _00002_;
  wire _00003_;
  wire _00004_;
  wire [31:0] _00005_;
  wire [4:0] _00006_;
  wire [4:0] _00007_;
  wire [4:0] _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  wire _09001_;
  wire _09002_;
  wire _09003_;
  wire _09004_;
  wire _09005_;
  wire _09006_;
  wire _09007_;
  wire _09008_;
  wire _09009_;
  wire _09010_;
  wire _09011_;
  wire _09012_;
  wire _09013_;
  wire _09014_;
  wire _09015_;
  wire _09016_;
  wire _09017_;
  wire _09018_;
  wire _09019_;
  wire _09020_;
  wire _09021_;
  wire _09022_;
  wire _09023_;
  wire _09024_;
  wire _09025_;
  wire _09026_;
  wire _09027_;
  wire _09028_;
  wire _09029_;
  wire _09030_;
  wire _09031_;
  wire _09032_;
  wire _09033_;
  wire _09034_;
  wire _09035_;
  wire _09036_;
  wire _09037_;
  wire _09038_;
  wire _09039_;
  wire _09040_;
  wire _09041_;
  wire _09042_;
  wire _09043_;
  wire _09044_;
  wire _09045_;
  wire _09046_;
  wire _09047_;
  wire _09048_;
  wire _09049_;
  wire _09050_;
  wire _09051_;
  wire _09052_;
  wire _09053_;
  wire _09054_;
  wire _09055_;
  wire _09056_;
  wire _09057_;
  wire _09058_;
  wire _09059_;
  wire _09060_;
  wire _09061_;
  wire _09062_;
  wire _09063_;
  wire _09064_;
  wire _09065_;
  wire _09066_;
  wire _09067_;
  wire _09068_;
  wire _09069_;
  wire _09070_;
  wire _09071_;
  wire _09072_;
  wire _09073_;
  wire _09074_;
  wire _09075_;
  wire _09076_;
  wire _09077_;
  wire _09078_;
  wire _09079_;
  wire _09080_;
  wire _09081_;
  wire _09082_;
  wire _09083_;
  wire _09084_;
  wire _09085_;
  wire _09086_;
  wire _09087_;
  wire _09088_;
  wire _09089_;
  wire _09090_;
  wire _09091_;
  wire _09092_;
  wire _09093_;
  wire _09094_;
  wire _09095_;
  wire _09096_;
  wire _09097_;
  wire _09098_;
  wire _09099_;
  wire _09100_;
  wire _09101_;
  wire _09102_;
  wire _09103_;
  wire _09104_;
  wire _09105_;
  wire _09106_;
  wire _09107_;
  wire _09108_;
  wire _09109_;
  wire _09110_;
  wire _09111_;
  wire _09112_;
  wire _09113_;
  wire _09114_;
  wire _09115_;
  wire _09116_;
  wire _09117_;
  wire _09118_;
  wire _09119_;
  wire _09120_;
  wire _09121_;
  wire _09122_;
  wire _09123_;
  wire _09124_;
  wire _09125_;
  wire _09126_;
  wire _09127_;
  wire _09128_;
  wire _09129_;
  wire _09130_;
  wire _09131_;
  wire _09132_;
  wire _09133_;
  wire _09134_;
  wire _09135_;
  wire _09136_;
  wire _09137_;
  wire _09138_;
  wire _09139_;
  wire _09140_;
  wire _09141_;
  wire _09142_;
  wire _09143_;
  wire _09144_;
  wire _09145_;
  wire _09146_;
  wire _09147_;
  wire _09148_;
  wire _09149_;
  wire _09150_;
  wire _09151_;
  wire _09152_;
  wire _09153_;
  wire _09154_;
  wire _09155_;
  wire _09156_;
  wire _09157_;
  wire _09158_;
  wire _09159_;
  wire _09160_;
  wire _09161_;
  wire _09162_;
  wire _09163_;
  wire _09164_;
  wire _09165_;
  wire _09166_;
  wire _09167_;
  wire _09168_;
  wire _09169_;
  wire _09170_;
  wire _09171_;
  wire _09172_;
  wire _09173_;
  wire _09174_;
  wire _09175_;
  wire _09176_;
  wire _09177_;
  wire _09178_;
  wire _09179_;
  wire _09180_;
  wire _09181_;
  wire _09182_;
  wire _09183_;
  wire _09184_;
  wire _09185_;
  wire _09186_;
  wire _09187_;
  wire _09188_;
  wire _09189_;
  wire _09190_;
  wire _09191_;
  wire _09192_;
  wire _09193_;
  wire _09194_;
  wire _09195_;
  wire _09196_;
  wire _09197_;
  wire _09198_;
  wire _09199_;
  wire _09200_;
  wire _09201_;
  wire _09202_;
  wire _09203_;
  wire _09204_;
  wire _09205_;
  wire _09206_;
  wire _09207_;
  wire _09208_;
  wire _09209_;
  wire _09210_;
  wire _09211_;
  wire _09212_;
  wire _09213_;
  wire _09214_;
  wire _09215_;
  wire _09216_;
  wire _09217_;
  wire _09218_;
  wire _09219_;
  wire _09220_;
  wire _09221_;
  wire _09222_;
  wire _09223_;
  wire _09224_;
  wire _09225_;
  wire _09226_;
  wire _09227_;
  wire _09228_;
  wire _09229_;
  wire _09230_;
  wire _09231_;
  wire _09232_;
  wire _09233_;
  wire _09234_;
  wire _09235_;
  wire _09236_;
  wire _09237_;
  wire _09238_;
  wire _09239_;
  wire _09240_;
  wire _09241_;
  wire _09242_;
  wire _09243_;
  wire _09244_;
  wire _09245_;
  wire _09246_;
  wire _09247_;
  wire _09248_;
  wire _09249_;
  wire _09250_;
  wire _09251_;
  wire _09252_;
  wire _09253_;
  wire _09254_;
  wire _09255_;
  wire _09256_;
  wire _09257_;
  wire _09258_;
  wire _09259_;
  wire _09260_;
  wire _09261_;
  wire _09262_;
  wire _09263_;
  wire _09264_;
  wire _09265_;
  wire _09266_;
  wire _09267_;
  wire _09268_;
  wire _09269_;
  wire _09270_;
  wire _09271_;
  wire _09272_;
  wire _09273_;
  wire _09274_;
  wire _09275_;
  wire _09276_;
  wire _09277_;
  wire _09278_;
  wire _09279_;
  wire _09280_;
  wire _09281_;
  wire _09282_;
  wire _09283_;
  wire _09284_;
  wire _09285_;
  wire _09286_;
  wire _09287_;
  wire _09288_;
  wire _09289_;
  wire _09290_;
  wire _09291_;
  wire _09292_;
  wire _09293_;
  wire _09294_;
  wire _09295_;
  wire _09296_;
  wire _09297_;
  wire _09298_;
  wire _09299_;
  wire _09300_;
  wire _09301_;
  wire _09302_;
  wire _09303_;
  wire _09304_;
  wire _09305_;
  wire _09306_;
  wire _09307_;
  wire _09308_;
  wire _09309_;
  wire _09310_;
  wire _09311_;
  wire _09312_;
  wire _09313_;
  wire _09314_;
  wire _09315_;
  wire _09316_;
  wire _09317_;
  wire _09318_;
  wire _09319_;
  wire _09320_;
  wire _09321_;
  wire _09322_;
  wire _09323_;
  wire _09324_;
  wire _09325_;
  wire _09326_;
  wire _09327_;
  wire _09328_;
  wire _09329_;
  wire _09330_;
  wire _09331_;
  wire _09332_;
  wire _09333_;
  wire _09334_;
  wire _09335_;
  wire _09336_;
  wire _09337_;
  wire _09338_;
  wire _09339_;
  wire _09340_;
  wire _09341_;
  wire _09342_;
  wire _09343_;
  wire _09344_;
  wire _09345_;
  wire _09346_;
  wire _09347_;
  wire _09348_;
  wire _09349_;
  wire _09350_;
  wire _09351_;
  wire _09352_;
  wire _09353_;
  wire _09354_;
  wire _09355_;
  wire _09356_;
  wire _09357_;
  wire _09358_;
  wire _09359_;
  wire _09360_;
  wire _09361_;
  wire _09362_;
  wire _09363_;
  wire _09364_;
  wire _09365_;
  wire _09366_;
  wire _09367_;
  wire _09368_;
  wire _09369_;
  wire _09370_;
  wire _09371_;
  wire _09372_;
  wire _09373_;
  wire _09374_;
  wire _09375_;
  wire _09376_;
  wire _09377_;
  wire _09378_;
  wire _09379_;
  wire _09380_;
  wire _09381_;
  wire _09382_;
  wire _09383_;
  wire _09384_;
  wire _09385_;
  wire _09386_;
  wire _09387_;
  wire _09388_;
  wire _09389_;
  wire _09390_;
  wire _09391_;
  wire _09392_;
  wire _09393_;
  wire _09394_;
  wire _09395_;
  wire _09396_;
  wire _09397_;
  wire _09398_;
  wire _09399_;
  wire _09400_;
  wire _09401_;
  wire _09402_;
  wire _09403_;
  wire _09404_;
  wire _09405_;
  wire _09406_;
  wire _09407_;
  wire _09408_;
  wire _09409_;
  wire _09410_;
  wire _09411_;
  wire _09412_;
  wire _09413_;
  wire _09414_;
  wire _09415_;
  wire _09416_;
  wire _09417_;
  wire _09418_;
  wire _09419_;
  wire _09420_;
  wire _09421_;
  wire _09422_;
  wire _09423_;
  wire _09424_;
  wire _09425_;
  wire _09426_;
  wire _09427_;
  wire _09428_;
  wire _09429_;
  wire _09430_;
  wire _09431_;
  wire _09432_;
  wire _09433_;
  wire _09434_;
  wire _09435_;
  wire _09436_;
  wire _09437_;
  wire _09438_;
  wire _09439_;
  wire _09440_;
  wire _09441_;
  wire _09442_;
  wire _09443_;
  wire _09444_;
  wire _09445_;
  wire _09446_;
  wire _09447_;
  wire _09448_;
  wire _09449_;
  wire _09450_;
  wire _09451_;
  wire _09452_;
  wire _09453_;
  wire _09454_;
  wire _09455_;
  wire _09456_;
  wire _09457_;
  wire _09458_;
  wire _09459_;
  wire _09460_;
  wire _09461_;
  wire _09462_;
  wire _09463_;
  wire _09464_;
  wire _09465_;
  wire _09466_;
  wire _09467_;
  wire _09468_;
  wire _09469_;
  wire _09470_;
  wire _09471_;
  wire _09472_;
  wire _09473_;
  wire _09474_;
  wire _09475_;
  wire _09476_;
  wire _09477_;
  wire _09478_;
  wire _09479_;
  wire _09480_;
  wire _09481_;
  wire _09482_;
  wire _09483_;
  wire _09484_;
  wire _09485_;
  wire _09486_;
  wire _09487_;
  wire _09488_;
  wire _09489_;
  wire _09490_;
  wire _09491_;
  wire _09492_;
  wire _09493_;
  wire _09494_;
  wire _09495_;
  wire _09496_;
  wire _09497_;
  wire _09498_;
  wire _09499_;
  wire _09500_;
  wire _09501_;
  wire _09502_;
  wire _09503_;
  wire _09504_;
  wire _09505_;
  wire _09506_;
  wire _09507_;
  wire _09508_;
  wire _09509_;
  wire _09510_;
  wire _09511_;
  wire _09512_;
  wire _09513_;
  wire _09514_;
  wire _09515_;
  wire _09516_;
  wire _09517_;
  wire _09518_;
  wire _09519_;
  wire _09520_;
  wire _09521_;
  wire _09522_;
  wire _09523_;
  wire _09524_;
  wire _09525_;
  wire _09526_;
  wire _09527_;
  wire _09528_;
  wire _09529_;
  wire _09530_;
  wire _09531_;
  wire _09532_;
  wire _09533_;
  wire _09534_;
  wire _09535_;
  wire _09536_;
  wire _09537_;
  wire _09538_;
  wire _09539_;
  wire _09540_;
  wire _09541_;
  wire _09542_;
  wire _09543_;
  wire _09544_;
  wire _09545_;
  wire _09546_;
  wire _09547_;
  wire _09548_;
  wire _09549_;
  wire _09550_;
  wire _09551_;
  wire _09552_;
  wire _09553_;
  wire _09554_;
  wire _09555_;
  wire _09556_;
  wire _09557_;
  wire _09558_;
  wire _09559_;
  wire _09560_;
  wire _09561_;
  wire _09562_;
  wire _09563_;
  wire _09564_;
  wire _09565_;
  wire _09566_;
  wire _09567_;
  wire _09568_;
  wire _09569_;
  wire _09570_;
  wire _09571_;
  wire _09572_;
  wire _09573_;
  wire _09574_;
  wire _09575_;
  wire _09576_;
  wire _09577_;
  wire _09578_;
  wire _09579_;
  wire _09580_;
  wire _09581_;
  wire _09582_;
  wire _09583_;
  wire _09584_;
  wire _09585_;
  wire _09586_;
  wire _09587_;
  wire _09588_;
  wire _09589_;
  wire _09590_;
  wire _09591_;
  wire _09592_;
  wire _09593_;
  wire _09594_;
  wire _09595_;
  wire _09596_;
  wire _09597_;
  wire _09598_;
  wire _09599_;
  wire _09600_;
  wire _09601_;
  wire _09602_;
  wire _09603_;
  wire _09604_;
  wire _09605_;
  wire _09606_;
  wire _09607_;
  wire _09608_;
  wire _09609_;
  wire _09610_;
  wire _09611_;
  wire _09612_;
  wire _09613_;
  wire _09614_;
  wire _09615_;
  wire _09616_;
  wire _09617_;
  wire _09618_;
  wire _09619_;
  wire _09620_;
  wire _09621_;
  wire _09622_;
  wire _09623_;
  wire _09624_;
  wire _09625_;
  wire _09626_;
  wire _09627_;
  wire _09628_;
  wire _09629_;
  wire _09630_;
  wire _09631_;
  wire _09632_;
  wire _09633_;
  wire _09634_;
  wire _09635_;
  wire _09636_;
  wire _09637_;
  wire _09638_;
  wire _09639_;
  wire _09640_;
  wire _09641_;
  wire _09642_;
  wire _09643_;
  wire _09644_;
  wire _09645_;
  wire _09646_;
  wire _09647_;
  wire _09648_;
  wire _09649_;
  wire _09650_;
  wire _09651_;
  wire _09652_;
  wire _09653_;
  wire _09654_;
  wire _09655_;
  wire _09656_;
  wire _09657_;
  wire _09658_;
  wire _09659_;
  wire _09660_;
  wire _09661_;
  wire _09662_;
  wire _09663_;
  wire _09664_;
  wire _09665_;
  wire _09666_;
  wire _09667_;
  wire _09668_;
  wire _09669_;
  wire _09670_;
  wire _09671_;
  wire _09672_;
  wire _09673_;
  wire _09674_;
  wire _09675_;
  wire _09676_;
  wire _09677_;
  wire _09678_;
  wire _09679_;
  wire _09680_;
  wire _09681_;
  wire _09682_;
  wire _09683_;
  wire _09684_;
  wire _09685_;
  wire _09686_;
  wire _09687_;
  wire _09688_;
  wire _09689_;
  wire _09690_;
  wire _09691_;
  wire _09692_;
  wire _09693_;
  wire _09694_;
  wire _09695_;
  wire _09696_;
  wire _09697_;
  wire _09698_;
  wire _09699_;
  wire _09700_;
  wire _09701_;
  wire _09702_;
  wire _09703_;
  wire _09704_;
  wire _09705_;
  wire _09706_;
  wire _09707_;
  wire _09708_;
  wire _09709_;
  wire _09710_;
  wire _09711_;
  wire _09712_;
  wire _09713_;
  wire _09714_;
  wire _09715_;
  wire _09716_;
  wire _09717_;
  wire _09718_;
  wire _09719_;
  wire _09720_;
  wire _09721_;
  wire _09722_;
  wire _09723_;
  wire _09724_;
  wire _09725_;
  wire _09726_;
  wire _09727_;
  wire _09728_;
  wire _09729_;
  wire _09730_;
  wire _09731_;
  wire _09732_;
  wire _09733_;
  wire _09734_;
  wire _09735_;
  wire _09736_;
  wire _09737_;
  wire _09738_;
  wire _09739_;
  wire _09740_;
  wire _09741_;
  wire _09742_;
  wire _09743_;
  wire _09744_;
  wire _09745_;
  wire _09746_;
  wire _09747_;
  wire _09748_;
  wire _09749_;
  wire _09750_;
  wire _09751_;
  wire _09752_;
  wire _09753_;
  wire _09754_;
  wire _09755_;
  wire _09756_;
  wire _09757_;
  wire _09758_;
  wire _09759_;
  wire _09760_;
  wire _09761_;
  wire _09762_;
  wire _09763_;
  wire _09764_;
  wire _09765_;
  wire _09766_;
  wire _09767_;
  wire _09768_;
  wire _09769_;
  wire _09770_;
  wire _09771_;
  wire _09772_;
  wire _09773_;
  wire _09774_;
  wire _09775_;
  wire _09776_;
  wire _09777_;
  wire _09778_;
  wire _09779_;
  wire _09780_;
  wire _09781_;
  wire _09782_;
  wire _09783_;
  wire _09784_;
  wire _09785_;
  wire _09786_;
  wire _09787_;
  wire _09788_;
  wire _09789_;
  wire _09790_;
  wire _09791_;
  wire _09792_;
  wire _09793_;
  wire _09794_;
  wire _09795_;
  wire _09796_;
  wire _09797_;
  wire _09798_;
  wire _09799_;
  wire _09800_;
  wire _09801_;
  wire _09802_;
  wire _09803_;
  wire _09804_;
  wire _09805_;
  wire _09806_;
  wire _09807_;
  wire _09808_;
  wire _09809_;
  wire _09810_;
  wire _09811_;
  wire _09812_;
  wire _09813_;
  wire _09814_;
  wire _09815_;
  wire _09816_;
  wire _09817_;
  wire _09818_;
  wire _09819_;
  wire _09820_;
  wire _09821_;
  wire _09822_;
  wire _09823_;
  wire _09824_;
  wire _09825_;
  wire _09826_;
  wire _09827_;
  wire _09828_;
  wire _09829_;
  wire _09830_;
  wire _09831_;
  wire _09832_;
  wire _09833_;
  wire _09834_;
  wire _09835_;
  wire _09836_;
  wire _09837_;
  wire _09838_;
  wire _09839_;
  wire _09840_;
  wire _09841_;
  wire _09842_;
  wire _09843_;
  wire _09844_;
  wire _09845_;
  wire _09846_;
  wire _09847_;
  wire _09848_;
  wire _09849_;
  wire _09850_;
  wire _09851_;
  wire _09852_;
  wire _09853_;
  wire _09854_;
  wire _09855_;
  wire _09856_;
  wire _09857_;
  wire _09858_;
  wire _09859_;
  wire _09860_;
  wire _09861_;
  wire _09862_;
  wire _09863_;
  wire _09864_;
  wire _09865_;
  wire _09866_;
  wire _09867_;
  wire _09868_;
  wire _09869_;
  wire _09870_;
  wire _09871_;
  wire _09872_;
  wire _09873_;
  wire _09874_;
  wire _09875_;
  wire _09876_;
  wire _09877_;
  wire _09878_;
  wire _09879_;
  wire _09880_;
  wire _09881_;
  wire _09882_;
  wire _09883_;
  wire _09884_;
  wire _09885_;
  wire _09886_;
  wire _09887_;
  wire _09888_;
  wire _09889_;
  wire _09890_;
  wire _09891_;
  wire _09892_;
  wire _09893_;
  wire _09894_;
  wire _09895_;
  wire _09896_;
  wire _09897_;
  wire _09898_;
  wire _09899_;
  wire _09900_;
  wire _09901_;
  wire _09902_;
  wire _09903_;
  wire _09904_;
  wire _09905_;
  wire _09906_;
  wire _09907_;
  wire _09908_;
  wire _09909_;
  wire _09910_;
  wire _09911_;
  wire _09912_;
  wire _09913_;
  wire _09914_;
  wire _09915_;
  wire _09916_;
  wire _09917_;
  wire _09918_;
  wire _09919_;
  wire _09920_;
  wire _09921_;
  wire _09922_;
  wire _09923_;
  wire _09924_;
  wire _09925_;
  wire _09926_;
  wire _09927_;
  wire _09928_;
  wire _09929_;
  wire _09930_;
  wire _09931_;
  wire _09932_;
  wire _09933_;
  wire _09934_;
  wire _09935_;
  wire _09936_;
  wire _09937_;
  wire _09938_;
  wire _09939_;
  wire _09940_;
  wire _09941_;
  wire _09942_;
  wire _09943_;
  wire _09944_;
  wire _09945_;
  wire _09946_;
  wire _09947_;
  wire _09948_;
  wire _09949_;
  wire _09950_;
  wire _09951_;
  wire _09952_;
  wire _09953_;
  wire _09954_;
  wire _09955_;
  wire _09956_;
  wire _09957_;
  wire _09958_;
  wire _09959_;
  wire _09960_;
  wire _09961_;
  wire _09962_;
  wire _09963_;
  wire _09964_;
  wire _09965_;
  wire _09966_;
  wire _09967_;
  wire _09968_;
  wire _09969_;
  wire _09970_;
  wire _09971_;
  wire _09972_;
  wire _09973_;
  wire _09974_;
  wire _09975_;
  wire _09976_;
  wire _09977_;
  wire _09978_;
  wire _09979_;
  wire _09980_;
  wire _09981_;
  wire _09982_;
  wire _09983_;
  wire _09984_;
  wire _09985_;
  wire _09986_;
  wire _09987_;
  wire _09988_;
  wire _09989_;
  wire _09990_;
  wire _09991_;
  wire _09992_;
  wire _09993_;
  wire _09994_;
  wire _09995_;
  wire _09996_;
  wire _09997_;
  wire _09998_;
  wire _09999_;
  wire _10000_;
  wire _10001_;
  wire _10002_;
  wire _10003_;
  wire _10004_;
  wire _10005_;
  wire _10006_;
  wire _10007_;
  wire _10008_;
  wire _10009_;
  wire _10010_;
  wire _10011_;
  wire _10012_;
  wire _10013_;
  wire _10014_;
  wire _10015_;
  wire _10016_;
  wire _10017_;
  wire _10018_;
  wire _10019_;
  wire _10020_;
  wire _10021_;
  wire _10022_;
  wire _10023_;
  wire _10024_;
  wire _10025_;
  wire _10026_;
  wire _10027_;
  wire _10028_;
  wire _10029_;
  wire _10030_;
  wire _10031_;
  wire _10032_;
  wire _10033_;
  wire _10034_;
  wire _10035_;
  wire _10036_;
  wire _10037_;
  wire _10038_;
  wire _10039_;
  wire _10040_;
  wire _10041_;
  wire _10042_;
  wire _10043_;
  wire _10044_;
  wire _10045_;
  wire _10046_;
  wire _10047_;
  wire _10048_;
  wire _10049_;
  wire _10050_;
  wire _10051_;
  wire _10052_;
  wire _10053_;
  wire _10054_;
  wire _10055_;
  wire _10056_;
  wire _10057_;
  wire _10058_;
  wire _10059_;
  wire _10060_;
  wire _10061_;
  wire _10062_;
  wire _10063_;
  wire _10064_;
  wire _10065_;
  wire _10066_;
  wire _10067_;
  wire _10068_;
  wire _10069_;
  wire _10070_;
  wire _10071_;
  wire _10072_;
  wire _10073_;
  wire _10074_;
  wire _10075_;
  wire _10076_;
  wire _10077_;
  wire _10078_;
  wire _10079_;
  wire _10080_;
  wire _10081_;
  wire _10082_;
  wire _10083_;
  wire _10084_;
  wire _10085_;
  wire _10086_;
  wire _10087_;
  wire _10088_;
  wire _10089_;
  wire _10090_;
  wire _10091_;
  wire _10092_;
  wire _10093_;
  wire _10094_;
  wire _10095_;
  wire _10096_;
  wire _10097_;
  wire _10098_;
  wire _10099_;
  wire _10100_;
  wire _10101_;
  wire _10102_;
  wire _10103_;
  wire _10104_;
  wire _10105_;
  wire _10106_;
  wire _10107_;
  wire _10108_;
  wire _10109_;
  wire _10110_;
  wire _10111_;
  wire _10112_;
  wire _10113_;
  wire _10114_;
  wire _10115_;
  wire _10116_;
  wire _10117_;
  wire _10118_;
  wire _10119_;
  wire _10120_;
  wire _10121_;
  wire _10122_;
  wire _10123_;
  wire _10124_;
  wire _10125_;
  wire _10126_;
  wire _10127_;
  wire _10128_;
  wire _10129_;
  wire _10130_;
  wire _10131_;
  wire _10132_;
  wire _10133_;
  wire _10134_;
  wire _10135_;
  wire _10136_;
  wire _10137_;
  wire _10138_;
  wire _10139_;
  wire _10140_;
  wire _10141_;
  wire _10142_;
  wire _10143_;
  wire _10144_;
  wire _10145_;
  wire _10146_;
  wire _10147_;
  wire _10148_;
  wire _10149_;
  wire _10150_;
  wire _10151_;
  wire _10152_;
  wire _10153_;
  wire _10154_;
  wire _10155_;
  wire _10156_;
  wire _10157_;
  wire _10158_;
  wire _10159_;
  wire _10160_;
  wire _10161_;
  wire _10162_;
  wire _10163_;
  wire _10164_;
  wire _10165_;
  wire _10166_;
  wire _10167_;
  wire _10168_;
  wire _10169_;
  wire _10170_;
  wire _10171_;
  wire _10172_;
  wire _10173_;
  wire _10174_;
  wire _10175_;
  wire _10176_;
  wire _10177_;
  wire _10178_;
  wire _10179_;
  wire _10180_;
  wire _10181_;
  wire _10182_;
  wire _10183_;
  wire _10184_;
  wire _10185_;
  wire _10186_;
  wire _10187_;
  wire _10188_;
  wire _10189_;
  wire _10190_;
  wire _10191_;
  wire _10192_;
  wire _10193_;
  wire _10194_;
  wire _10195_;
  wire _10196_;
  wire _10197_;
  wire _10198_;
  wire _10199_;
  wire _10200_;
  wire _10201_;
  wire _10202_;
  wire _10203_;
  wire _10204_;
  wire _10205_;
  wire _10206_;
  wire _10207_;
  wire _10208_;
  wire _10209_;
  wire _10210_;
  wire _10211_;
  wire _10212_;
  wire _10213_;
  wire _10214_;
  wire _10215_;
  wire _10216_;
  wire _10217_;
  wire _10218_;
  wire _10219_;
  wire _10220_;
  wire _10221_;
  wire _10222_;
  wire _10223_;
  wire _10224_;
  wire _10225_;
  wire _10226_;
  wire _10227_;
  wire _10228_;
  wire _10229_;
  wire _10230_;
  wire _10231_;
  wire _10232_;
  wire _10233_;
  wire _10234_;
  wire _10235_;
  wire _10236_;
  wire _10237_;
  wire _10238_;
  wire _10239_;
  wire _10240_;
  wire _10241_;
  wire _10242_;
  wire _10243_;
  wire _10244_;
  wire _10245_;
  wire _10246_;
  wire _10247_;
  wire _10248_;
  wire _10249_;
  wire _10250_;
  wire _10251_;
  wire _10252_;
  wire _10253_;
  wire _10254_;
  wire _10255_;
  wire _10256_;
  wire _10257_;
  wire _10258_;
  wire _10259_;
  wire _10260_;
  wire _10261_;
  wire _10262_;
  wire _10263_;
  wire _10264_;
  wire _10265_;
  wire _10266_;
  wire _10267_;
  wire _10268_;
  wire _10269_;
  wire _10270_;
  wire _10271_;
  wire _10272_;
  wire _10273_;
  wire _10274_;
  wire _10275_;
  wire _10276_;
  wire _10277_;
  wire _10278_;
  wire _10279_;
  wire _10280_;
  wire _10281_;
  wire _10282_;
  wire _10283_;
  wire _10284_;
  wire _10285_;
  wire _10286_;
  wire _10287_;
  wire _10288_;
  wire _10289_;
  wire _10290_;
  wire _10291_;
  wire _10292_;
  wire _10293_;
  wire _10294_;
  wire _10295_;
  wire _10296_;
  wire _10297_;
  wire _10298_;
  wire _10299_;
  wire _10300_;
  wire _10301_;
  wire _10302_;
  wire _10303_;
  wire _10304_;
  wire _10305_;
  wire _10306_;
  wire _10307_;
  wire _10308_;
  wire _10309_;
  wire _10310_;
  wire _10311_;
  wire _10312_;
  wire _10313_;
  wire _10314_;
  wire _10315_;
  wire _10316_;
  wire _10317_;
  wire _10318_;
  wire _10319_;
  wire _10320_;
  wire _10321_;
  wire _10322_;
  wire _10323_;
  wire _10324_;
  wire _10325_;
  wire _10326_;
  wire _10327_;
  wire _10328_;
  wire _10329_;
  wire _10330_;
  wire _10331_;
  wire _10332_;
  wire _10333_;
  wire _10334_;
  wire _10335_;
  wire _10336_;
  wire _10337_;
  wire _10338_;
  wire _10339_;
  wire _10340_;
  wire _10341_;
  wire _10342_;
  wire _10343_;
  wire _10344_;
  wire _10345_;
  wire _10346_;
  wire _10347_;
  wire _10348_;
  wire _10349_;
  wire _10350_;
  wire _10351_;
  wire _10352_;
  wire _10353_;
  wire _10354_;
  wire _10355_;
  wire _10356_;
  wire _10357_;
  wire _10358_;
  wire _10359_;
  wire _10360_;
  wire _10361_;
  wire _10362_;
  wire _10363_;
  wire _10364_;
  wire _10365_;
  wire _10366_;
  wire _10367_;
  wire _10368_;
  wire _10369_;
  wire _10370_;
  wire _10371_;
  wire _10372_;
  wire _10373_;
  wire _10374_;
  wire _10375_;
  wire _10376_;
  wire _10377_;
  wire _10378_;
  wire _10379_;
  wire _10380_;
  wire _10381_;
  wire _10382_;
  wire _10383_;
  wire _10384_;
  wire _10385_;
  wire _10386_;
  wire _10387_;
  wire _10388_;
  wire _10389_;
  wire _10390_;
  wire _10391_;
  wire _10392_;
  wire _10393_;
  wire _10394_;
  wire _10395_;
  wire _10396_;
  wire _10397_;
  wire _10398_;
  wire _10399_;
  wire _10400_;
  wire _10401_;
  wire _10402_;
  wire _10403_;
  wire _10404_;
  wire _10405_;
  wire _10406_;
  wire _10407_;
  wire _10408_;
  wire _10409_;
  wire _10410_;
  wire _10411_;
  wire _10412_;
  wire _10413_;
  wire _10414_;
  wire _10415_;
  wire _10416_;
  wire _10417_;
  wire _10418_;
  wire _10419_;
  wire _10420_;
  wire _10421_;
  wire _10422_;
  wire _10423_;
  wire _10424_;
  wire _10425_;
  wire _10426_;
  wire _10427_;
  wire _10428_;
  wire _10429_;
  wire _10430_;
  wire _10431_;
  wire _10432_;
  wire _10433_;
  wire _10434_;
  wire _10435_;
  wire _10436_;
  wire _10437_;
  wire _10438_;
  wire _10439_;
  wire _10440_;
  wire _10441_;
  wire _10442_;
  wire _10443_;
  wire _10444_;
  wire _10445_;
  wire _10446_;
  wire _10447_;
  wire _10448_;
  wire _10449_;
  wire _10450_;
  wire _10451_;
  wire _10452_;
  wire _10453_;
  wire _10454_;
  wire _10455_;
  wire _10456_;
  wire _10457_;
  wire _10458_;
  wire _10459_;
  wire _10460_;
  wire _10461_;
  wire _10462_;
  wire _10463_;
  wire _10464_;
  wire _10465_;
  wire _10466_;
  wire _10467_;
  wire _10468_;
  wire _10469_;
  wire _10470_;
  wire _10471_;
  wire _10472_;
  wire _10473_;
  wire _10474_;
  wire _10475_;
  wire _10476_;
  wire _10477_;
  wire _10478_;
  wire _10479_;
  wire _10480_;
  wire _10481_;
  wire _10482_;
  wire _10483_;
  wire _10484_;
  wire _10485_;
  wire _10486_;
  wire _10487_;
  wire _10488_;
  wire _10489_;
  wire _10490_;
  wire _10491_;
  wire _10492_;
  wire _10493_;
  wire _10494_;
  wire _10495_;
  wire _10496_;
  wire _10497_;
  wire _10498_;
  wire _10499_;
  wire _10500_;
  wire _10501_;
  wire _10502_;
  wire _10503_;
  wire _10504_;
  wire _10505_;
  wire _10506_;
  wire _10507_;
  wire _10508_;
  wire _10509_;
  wire _10510_;
  wire _10511_;
  wire _10512_;
  wire _10513_;
  wire _10514_;
  wire _10515_;
  wire _10516_;
  wire _10517_;
  wire _10518_;
  wire _10519_;
  wire _10520_;
  wire _10521_;
  wire _10522_;
  wire _10523_;
  wire _10524_;
  wire _10525_;
  wire _10526_;
  wire _10527_;
  wire _10528_;
  wire _10529_;
  wire _10530_;
  wire _10531_;
  wire _10532_;
  wire _10533_;
  wire _10534_;
  wire _10535_;
  wire _10536_;
  wire _10537_;
  wire _10538_;
  wire _10539_;
  wire _10540_;
  wire _10541_;
  wire _10542_;
  wire _10543_;
  wire _10544_;
  wire _10545_;
  wire _10546_;
  wire _10547_;
  wire _10548_;
  wire _10549_;
  wire _10550_;
  wire _10551_;
  wire _10552_;
  wire _10553_;
  wire _10554_;
  wire _10555_;
  wire _10556_;
  wire _10557_;
  wire _10558_;
  wire _10559_;
  wire _10560_;
  wire _10561_;
  wire _10562_;
  wire _10563_;
  wire _10564_;
  wire _10565_;
  wire _10566_;
  wire _10567_;
  wire _10568_;
  wire _10569_;
  wire _10570_;
  wire _10571_;
  wire _10572_;
  wire _10573_;
  wire _10574_;
  wire _10575_;
  wire _10576_;
  wire _10577_;
  wire _10578_;
  wire _10579_;
  wire _10580_;
  wire _10581_;
  wire _10582_;
  wire _10583_;
  wire _10584_;
  wire _10585_;
  wire _10586_;
  wire _10587_;
  wire _10588_;
  wire _10589_;
  wire _10590_;
  wire _10591_;
  wire _10592_;
  wire _10593_;
  wire _10594_;
  wire _10595_;
  wire _10596_;
  wire _10597_;
  wire _10598_;
  wire _10599_;
  wire _10600_;
  wire _10601_;
  wire _10602_;
  wire _10603_;
  wire _10604_;
  wire _10605_;
  wire _10606_;
  wire _10607_;
  wire _10608_;
  wire _10609_;
  wire _10610_;
  wire _10611_;
  wire _10612_;
  wire _10613_;
  wire _10614_;
  wire _10615_;
  wire _10616_;
  wire _10617_;
  wire _10618_;
  wire _10619_;
  wire _10620_;
  wire _10621_;
  wire _10622_;
  wire _10623_;
  wire _10624_;
  wire _10625_;
  wire _10626_;
  wire _10627_;
  wire _10628_;
  wire _10629_;
  wire _10630_;
  wire _10631_;
  wire _10632_;
  wire _10633_;
  wire _10634_;
  wire _10635_;
  wire _10636_;
  wire _10637_;
  wire _10638_;
  wire _10639_;
  wire _10640_;
  wire _10641_;
  wire _10642_;
  wire _10643_;
  wire _10644_;
  wire _10645_;
  wire _10646_;
  wire _10647_;
  wire _10648_;
  wire _10649_;
  wire _10650_;
  wire _10651_;
  wire _10652_;
  wire _10653_;
  wire _10654_;
  wire _10655_;
  wire _10656_;
  wire _10657_;
  wire _10658_;
  wire _10659_;
  wire _10660_;
  wire _10661_;
  wire _10662_;
  wire _10663_;
  wire _10664_;
  wire _10665_;
  wire _10666_;
  wire _10667_;
  wire _10668_;
  wire _10669_;
  wire _10670_;
  wire _10671_;
  wire _10672_;
  wire _10673_;
  wire _10674_;
  wire _10675_;
  wire _10676_;
  wire _10677_;
  wire _10678_;
  wire _10679_;
  wire _10680_;
  wire _10681_;
  wire _10682_;
  wire _10683_;
  wire _10684_;
  wire _10685_;
  wire _10686_;
  wire _10687_;
  wire _10688_;
  wire _10689_;
  wire _10690_;
  wire _10691_;
  wire _10692_;
  wire _10693_;
  wire _10694_;
  wire _10695_;
  wire _10696_;
  wire _10697_;
  wire _10698_;
  wire _10699_;
  wire _10700_;
  wire _10701_;
  wire _10702_;
  wire _10703_;
  wire _10704_;
  wire _10705_;
  wire _10706_;
  wire _10707_;
  wire _10708_;
  wire _10709_;
  wire _10710_;
  wire _10711_;
  wire _10712_;
  wire _10713_;
  wire _10714_;
  wire _10715_;
  wire _10716_;
  wire _10717_;
  wire _10718_;
  wire _10719_;
  wire _10720_;
  wire _10721_;
  wire _10722_;
  wire _10723_;
  wire _10724_;
  wire _10725_;
  wire _10726_;
  wire _10727_;
  wire _10728_;
  wire _10729_;
  wire _10730_;
  wire _10731_;
  wire _10732_;
  wire _10733_;
  wire _10734_;
  wire _10735_;
  wire _10736_;
  wire _10737_;
  wire _10738_;
  wire _10739_;
  wire _10740_;
  wire _10741_;
  wire _10742_;
  wire _10743_;
  wire _10744_;
  wire _10745_;
  wire _10746_;
  wire _10747_;
  wire _10748_;
  wire _10749_;
  wire _10750_;
  wire _10751_;
  wire _10752_;
  wire _10753_;
  wire _10754_;
  wire _10755_;
  wire _10756_;
  wire _10757_;
  wire _10758_;
  wire _10759_;
  wire _10760_;
  wire _10761_;
  wire _10762_;
  wire _10763_;
  wire _10764_;
  wire _10765_;
  wire _10766_;
  wire _10767_;
  wire _10768_;
  wire _10769_;
  wire _10770_;
  wire _10771_;
  wire _10772_;
  wire _10773_;
  wire _10774_;
  wire _10775_;
  wire _10776_;
  wire _10777_;
  wire _10778_;
  wire _10779_;
  wire _10780_;
  wire _10781_;
  wire _10782_;
  wire _10783_;
  wire _10784_;
  wire _10785_;
  wire _10786_;
  wire _10787_;
  wire _10788_;
  wire _10789_;
  wire _10790_;
  wire _10791_;
  wire _10792_;
  wire _10793_;
  wire _10794_;
  wire _10795_;
  wire _10796_;
  wire _10797_;
  wire _10798_;
  wire _10799_;
  wire _10800_;
  wire _10801_;
  wire _10802_;
  wire _10803_;
  wire _10804_;
  wire _10805_;
  wire _10806_;
  wire _10807_;
  wire _10808_;
  wire _10809_;
  wire _10810_;
  wire _10811_;
  wire _10812_;
  wire _10813_;
  wire _10814_;
  wire _10815_;
  wire _10816_;
  wire _10817_;
  wire _10818_;
  wire _10819_;
  wire _10820_;
  wire _10821_;
  wire _10822_;
  wire _10823_;
  wire _10824_;
  wire _10825_;
  wire _10826_;
  wire _10827_;
  wire _10828_;
  wire _10829_;
  wire _10830_;
  wire _10831_;
  wire _10832_;
  wire _10833_;
  wire _10834_;
  wire _10835_;
  wire _10836_;
  wire _10837_;
  wire _10838_;
  wire _10839_;
  wire _10840_;
  wire _10841_;
  wire _10842_;
  wire _10843_;
  wire _10844_;
  wire _10845_;
  wire _10846_;
  wire _10847_;
  wire _10848_;
  wire _10849_;
  wire _10850_;
  wire _10851_;
  wire _10852_;
  wire _10853_;
  wire _10854_;
  wire _10855_;
  wire _10856_;
  wire _10857_;
  wire _10858_;
  wire _10859_;
  wire _10860_;
  wire _10861_;
  wire _10862_;
  wire _10863_;
  wire _10864_;
  wire _10865_;
  wire _10866_;
  wire _10867_;
  wire _10868_;
  wire _10869_;
  wire _10870_;
  wire _10871_;
  wire _10872_;
  wire _10873_;
  wire _10874_;
  wire _10875_;
  wire _10876_;
  wire _10877_;
  wire _10878_;
  wire _10879_;
  wire _10880_;
  wire _10881_;
  wire _10882_;
  wire _10883_;
  wire _10884_;
  wire _10885_;
  wire _10886_;
  wire _10887_;
  wire _10888_;
  wire _10889_;
  wire _10890_;
  wire _10891_;
  wire _10892_;
  wire _10893_;
  wire _10894_;
  wire _10895_;
  wire _10896_;
  wire _10897_;
  wire _10898_;
  wire _10899_;
  wire _10900_;
  wire _10901_;
  wire _10902_;
  wire _10903_;
  wire _10904_;
  wire _10905_;
  wire _10906_;
  wire _10907_;
  wire _10908_;
  wire _10909_;
  wire _10910_;
  wire _10911_;
  wire _10912_;
  wire _10913_;
  wire _10914_;
  wire _10915_;
  wire _10916_;
  wire _10917_;
  wire _10918_;
  wire _10919_;
  wire _10920_;
  wire _10921_;
  wire _10922_;
  wire _10923_;
  wire _10924_;
  wire _10925_;
  wire _10926_;
  wire _10927_;
  wire _10928_;
  wire _10929_;
  wire _10930_;
  wire _10931_;
  wire _10932_;
  wire _10933_;
  wire _10934_;
  wire _10935_;
  wire _10936_;
  wire _10937_;
  wire _10938_;
  wire _10939_;
  wire _10940_;
  wire _10941_;
  wire _10942_;
  wire _10943_;
  wire _10944_;
  wire _10945_;
  wire _10946_;
  wire _10947_;
  wire _10948_;
  wire _10949_;
  wire _10950_;
  wire _10951_;
  wire _10952_;
  wire _10953_;
  wire _10954_;
  wire _10955_;
  wire _10956_;
  wire _10957_;
  wire _10958_;
  wire _10959_;
  wire _10960_;
  wire _10961_;
  wire _10962_;
  wire _10963_;
  wire _10964_;
  wire _10965_;
  wire _10966_;
  wire _10967_;
  wire _10968_;
  wire _10969_;
  wire _10970_;
  wire _10971_;
  wire _10972_;
  wire _10973_;
  wire _10974_;
  wire _10975_;
  wire _10976_;
  wire _10977_;
  wire _10978_;
  wire _10979_;
  wire _10980_;
  wire _10981_;
  wire _10982_;
  wire _10983_;
  wire _10984_;
  wire _10985_;
  wire _10986_;
  wire _10987_;
  wire _10988_;
  wire _10989_;
  wire _10990_;
  wire _10991_;
  wire _10992_;
  wire _10993_;
  wire _10994_;
  wire _10995_;
  wire _10996_;
  wire _10997_;
  wire _10998_;
  wire _10999_;
  wire _11000_;
  wire _11001_;
  wire _11002_;
  wire _11003_;
  wire _11004_;
  wire _11005_;
  wire _11006_;
  wire _11007_;
  wire _11008_;
  wire _11009_;
  wire _11010_;
  wire _11011_;
  wire _11012_;
  wire _11013_;
  wire _11014_;
  wire _11015_;
  wire _11016_;
  wire _11017_;
  wire _11018_;
  wire _11019_;
  wire _11020_;
  wire _11021_;
  wire _11022_;
  wire _11023_;
  wire _11024_;
  wire _11025_;
  wire _11026_;
  wire _11027_;
  wire _11028_;
  wire _11029_;
  wire _11030_;
  wire _11031_;
  wire _11032_;
  wire _11033_;
  wire _11034_;
  wire _11035_;
  wire _11036_;
  wire _11037_;
  wire _11038_;
  wire _11039_;
  wire _11040_;
  wire _11041_;
  wire _11042_;
  wire _11043_;
  wire _11044_;
  wire _11045_;
  wire _11046_;
  wire _11047_;
  wire _11048_;
  wire _11049_;
  wire _11050_;
  wire _11051_;
  wire _11052_;
  wire _11053_;
  wire _11054_;
  wire _11055_;
  wire _11056_;
  wire _11057_;
  wire _11058_;
  wire _11059_;
  wire _11060_;
  wire _11061_;
  wire _11062_;
  wire _11063_;
  wire _11064_;
  wire _11065_;
  wire _11066_;
  wire _11067_;
  wire _11068_;
  wire _11069_;
  wire _11070_;
  wire _11071_;
  wire _11072_;
  wire _11073_;
  wire _11074_;
  wire _11075_;
  wire _11076_;
  wire _11077_;
  wire _11078_;
  wire _11079_;
  wire _11080_;
  wire _11081_;
  wire _11082_;
  wire _11083_;
  wire _11084_;
  wire _11085_;
  wire _11086_;
  wire _11087_;
  wire _11088_;
  wire _11089_;
  wire _11090_;
  wire _11091_;
  wire _11092_;
  wire _11093_;
  wire _11094_;
  wire _11095_;
  wire _11096_;
  wire _11097_;
  wire _11098_;
  wire _11099_;
  wire _11100_;
  wire _11101_;
  wire _11102_;
  wire _11103_;
  wire _11104_;
  wire _11105_;
  wire _11106_;
  wire _11107_;
  wire _11108_;
  wire _11109_;
  wire _11110_;
  wire _11111_;
  wire _11112_;
  wire _11113_;
  wire _11114_;
  wire _11115_;
  wire _11116_;
  wire _11117_;
  wire _11118_;
  wire _11119_;
  wire _11120_;
  wire _11121_;
  wire _11122_;
  wire _11123_;
  wire _11124_;
  wire _11125_;
  wire _11126_;
  wire _11127_;
  wire _11128_;
  wire _11129_;
  wire _11130_;
  wire _11131_;
  wire _11132_;
  wire _11133_;
  wire _11134_;
  wire _11135_;
  wire _11136_;
  wire _11137_;
  wire _11138_;
  wire _11139_;
  wire _11140_;
  wire _11141_;
  wire _11142_;
  wire _11143_;
  wire _11144_;
  wire _11145_;
  wire _11146_;
  wire _11147_;
  wire _11148_;
  wire _11149_;
  wire _11150_;
  wire _11151_;
  wire _11152_;
  wire _11153_;
  wire _11154_;
  wire _11155_;
  wire _11156_;
  wire _11157_;
  wire _11158_;
  wire _11159_;
  wire _11160_;
  wire _11161_;
  wire _11162_;
  wire _11163_;
  wire _11164_;
  wire _11165_;
  wire _11166_;
  wire _11167_;
  wire _11168_;
  wire _11169_;
  wire _11170_;
  wire _11171_;
  wire _11172_;
  wire _11173_;
  wire _11174_;
  wire _11175_;
  wire _11176_;
  wire _11177_;
  wire _11178_;
  wire _11179_;
  wire _11180_;
  wire _11181_;
  wire _11182_;
  wire _11183_;
  wire _11184_;
  wire _11185_;
  wire _11186_;
  wire _11187_;
  wire _11188_;
  wire _11189_;
  wire _11190_;
  wire _11191_;
  wire _11192_;
  wire _11193_;
  wire _11194_;
  wire _11195_;
  wire _11196_;
  wire _11197_;
  wire _11198_;
  wire _11199_;
  wire _11200_;
  wire _11201_;
  wire _11202_;
  wire _11203_;
  wire _11204_;
  wire _11205_;
  wire _11206_;
  wire _11207_;
  wire _11208_;
  wire _11209_;
  wire _11210_;
  wire _11211_;
  wire _11212_;
  wire _11213_;
  wire _11214_;
  wire _11215_;
  wire _11216_;
  wire _11217_;
  wire _11218_;
  wire _11219_;
  wire _11220_;
  wire _11221_;
  wire _11222_;
  wire _11223_;
  wire _11224_;
  wire _11225_;
  wire _11226_;
  wire _11227_;
  wire _11228_;
  wire _11229_;
  wire _11230_;
  wire _11231_;
  wire _11232_;
  wire _11233_;
  wire _11234_;
  wire _11235_;
  wire _11236_;
  wire _11237_;
  wire _11238_;
  wire _11239_;
  wire _11240_;
  wire _11241_;
  wire _11242_;
  wire _11243_;
  wire _11244_;
  wire _11245_;
  wire _11246_;
  wire _11247_;
  wire _11248_;
  wire _11249_;
  wire _11250_;
  wire _11251_;
  wire _11252_;
  wire _11253_;
  wire _11254_;
  wire _11255_;
  wire _11256_;
  wire _11257_;
  wire _11258_;
  wire _11259_;
  wire _11260_;
  wire _11261_;
  wire _11262_;
  wire _11263_;
  wire _11264_;
  wire _11265_;
  wire _11266_;
  wire _11267_;
  wire _11268_;
  wire _11269_;
  wire _11270_;
  wire _11271_;
  wire _11272_;
  wire _11273_;
  wire _11274_;
  wire _11275_;
  wire _11276_;
  wire _11277_;
  wire _11278_;
  wire _11279_;
  wire _11280_;
  wire _11281_;
  wire _11282_;
  wire _11283_;
  wire _11284_;
  wire _11285_;
  wire _11286_;
  wire _11287_;
  wire _11288_;
  wire _11289_;
  wire _11290_;
  wire _11291_;
  wire _11292_;
  wire _11293_;
  wire _11294_;
  wire _11295_;
  wire _11296_;
  wire _11297_;
  wire _11298_;
  wire _11299_;
  wire _11300_;
  wire _11301_;
  wire _11302_;
  wire _11303_;
  wire _11304_;
  wire _11305_;
  wire _11306_;
  wire _11307_;
  wire _11308_;
  wire _11309_;
  wire _11310_;
  wire _11311_;
  wire _11312_;
  wire _11313_;
  wire _11314_;
  wire _11315_;
  wire _11316_;
  wire _11317_;
  wire _11318_;
  wire _11319_;
  wire _11320_;
  wire _11321_;
  wire _11322_;
  wire _11323_;
  wire _11324_;
  wire _11325_;
  wire _11326_;
  wire _11327_;
  wire _11328_;
  wire _11329_;
  wire _11330_;
  wire _11331_;
  wire _11332_;
  wire _11333_;
  wire _11334_;
  wire _11335_;
  wire _11336_;
  wire _11337_;
  wire _11338_;
  wire _11339_;
  wire _11340_;
  wire _11341_;
  wire _11342_;
  wire _11343_;
  wire _11344_;
  wire _11345_;
  wire _11346_;
  wire _11347_;
  wire _11348_;
  wire _11349_;
  wire _11350_;
  wire _11351_;
  wire _11352_;
  wire _11353_;
  wire _11354_;
  wire _11355_;
  wire _11356_;
  wire _11357_;
  wire _11358_;
  wire _11359_;
  wire _11360_;
  wire _11361_;
  wire _11362_;
  wire _11363_;
  wire _11364_;
  wire _11365_;
  wire _11366_;
  wire _11367_;
  wire _11368_;
  wire _11369_;
  wire _11370_;
  wire _11371_;
  wire _11372_;
  wire _11373_;
  wire _11374_;
  wire _11375_;
  wire _11376_;
  wire _11377_;
  wire _11378_;
  wire _11379_;
  wire _11380_;
  wire _11381_;
  wire _11382_;
  wire _11383_;
  wire _11384_;
  wire _11385_;
  wire _11386_;
  wire _11387_;
  wire _11388_;
  wire _11389_;
  wire _11390_;
  wire _11391_;
  wire _11392_;
  wire _11393_;
  wire _11394_;
  wire _11395_;
  wire _11396_;
  wire _11397_;
  wire _11398_;
  wire _11399_;
  wire _11400_;
  wire _11401_;
  wire _11402_;
  wire _11403_;
  wire _11404_;
  wire _11405_;
  wire _11406_;
  wire _11407_;
  wire _11408_;
  wire _11409_;
  wire _11410_;
  wire _11411_;
  wire _11412_;
  wire _11413_;
  wire _11414_;
  wire _11415_;
  wire _11416_;
  wire _11417_;
  wire _11418_;
  wire _11419_;
  wire _11420_;
  wire _11421_;
  wire _11422_;
  wire _11423_;
  wire _11424_;
  wire _11425_;
  wire _11426_;
  wire _11427_;
  wire _11428_;
  wire _11429_;
  wire _11430_;
  wire _11431_;
  wire _11432_;
  wire _11433_;
  wire _11434_;
  wire _11435_;
  wire _11436_;
  wire _11437_;
  wire _11438_;
  wire _11439_;
  wire _11440_;
  wire _11441_;
  wire _11442_;
  wire _11443_;
  wire _11444_;
  wire _11445_;
  wire _11446_;
  wire _11447_;
  wire _11448_;
  wire _11449_;
  wire _11450_;
  wire _11451_;
  wire _11452_;
  wire _11453_;
  wire _11454_;
  wire _11455_;
  wire _11456_;
  wire _11457_;
  wire _11458_;
  wire _11459_;
  wire _11460_;
  wire _11461_;
  wire _11462_;
  wire _11463_;
  wire _11464_;
  wire _11465_;
  wire _11466_;
  wire _11467_;
  wire _11468_;
  wire _11469_;
  wire _11470_;
  wire _11471_;
  wire _11472_;
  wire _11473_;
  wire _11474_;
  wire _11475_;
  wire _11476_;
  wire _11477_;
  wire _11478_;
  wire _11479_;
  wire _11480_;
  wire _11481_;
  wire _11482_;
  wire _11483_;
  wire _11484_;
  wire _11485_;
  wire _11486_;
  wire _11487_;
  wire _11488_;
  wire _11489_;
  wire _11490_;
  wire _11491_;
  wire _11492_;
  wire _11493_;
  wire _11494_;
  wire _11495_;
  wire _11496_;
  wire _11497_;
  wire _11498_;
  wire _11499_;
  wire _11500_;
  wire _11501_;
  wire _11502_;
  wire _11503_;
  wire _11504_;
  wire _11505_;
  wire _11506_;
  wire _11507_;
  wire _11508_;
  wire _11509_;
  wire _11510_;
  wire _11511_;
  wire _11512_;
  wire _11513_;
  wire _11514_;
  wire _11515_;
  wire _11516_;
  wire _11517_;
  wire _11518_;
  wire _11519_;
  wire _11520_;
  wire _11521_;
  wire _11522_;
  wire _11523_;
  wire _11524_;
  wire _11525_;
  wire _11526_;
  wire _11527_;
  wire _11528_;
  wire _11529_;
  wire _11530_;
  wire _11531_;
  wire _11532_;
  wire _11533_;
  wire _11534_;
  wire _11535_;
  wire _11536_;
  wire _11537_;
  wire _11538_;
  wire _11539_;
  wire _11540_;
  wire _11541_;
  wire _11542_;
  wire _11543_;
  wire _11544_;
  wire _11545_;
  wire _11546_;
  wire _11547_;
  wire _11548_;
  wire _11549_;
  wire _11550_;
  wire _11551_;
  wire _11552_;
  wire _11553_;
  wire _11554_;
  wire _11555_;
  wire _11556_;
  wire _11557_;
  wire _11558_;
  wire _11559_;
  wire _11560_;
  wire _11561_;
  wire _11562_;
  wire _11563_;
  wire _11564_;
  wire _11565_;
  wire _11566_;
  wire _11567_;
  wire _11568_;
  wire _11569_;
  wire _11570_;
  wire _11571_;
  wire _11572_;
  wire _11573_;
  wire _11574_;
  wire _11575_;
  wire _11576_;
  wire _11577_;
  wire _11578_;
  wire _11579_;
  wire _11580_;
  wire _11581_;
  wire _11582_;
  wire _11583_;
  wire _11584_;
  wire _11585_;
  wire _11586_;
  wire _11587_;
  wire _11588_;
  wire _11589_;
  wire _11590_;
  wire _11591_;
  wire _11592_;
  wire _11593_;
  wire _11594_;
  wire _11595_;
  wire _11596_;
  wire _11597_;
  wire _11598_;
  wire _11599_;
  wire _11600_;
  wire _11601_;
  wire _11602_;
  wire _11603_;
  wire _11604_;
  wire _11605_;
  wire _11606_;
  wire _11607_;
  wire _11608_;
  wire _11609_;
  wire _11610_;
  wire _11611_;
  wire _11612_;
  wire _11613_;
  wire _11614_;
  wire _11615_;
  wire _11616_;
  wire _11617_;
  wire _11618_;
  wire _11619_;
  wire _11620_;
  wire _11621_;
  wire _11622_;
  wire _11623_;
  wire _11624_;
  wire _11625_;
  wire _11626_;
  wire _11627_;
  wire _11628_;
  wire _11629_;
  wire _11630_;
  wire _11631_;
  wire _11632_;
  wire _11633_;
  wire _11634_;
  wire _11635_;
  wire _11636_;
  wire _11637_;
  wire _11638_;
  wire _11639_;
  wire _11640_;
  wire _11641_;
  wire _11642_;
  wire _11643_;
  wire _11644_;
  wire _11645_;
  wire _11646_;
  wire _11647_;
  wire _11648_;
  wire _11649_;
  wire _11650_;
  wire _11651_;
  wire _11652_;
  wire _11653_;
  wire _11654_;
  wire _11655_;
  wire _11656_;
  wire _11657_;
  wire _11658_;
  wire _11659_;
  wire _11660_;
  wire _11661_;
  wire _11662_;
  wire _11663_;
  wire _11664_;
  wire _11665_;
  wire _11666_;
  wire _11667_;
  wire _11668_;
  wire _11669_;
  wire _11670_;
  wire _11671_;
  wire _11672_;
  wire _11673_;
  wire _11674_;
  wire _11675_;
  wire _11676_;
  wire _11677_;
  wire _11678_;
  wire _11679_;
  wire _11680_;
  wire _11681_;
  wire _11682_;
  wire _11683_;
  wire _11684_;
  wire _11685_;
  wire _11686_;
  wire _11687_;
  wire _11688_;
  wire _11689_;
  wire _11690_;
  wire _11691_;
  wire _11692_;
  wire _11693_;
  wire _11694_;
  wire _11695_;
  wire _11696_;
  wire _11697_;
  wire _11698_;
  wire _11699_;
  wire _11700_;
  wire _11701_;
  wire _11702_;
  wire _11703_;
  wire _11704_;
  wire _11705_;
  wire _11706_;
  wire _11707_;
  wire _11708_;
  wire _11709_;
  wire _11710_;
  wire _11711_;
  wire _11712_;
  wire _11713_;
  wire _11714_;
  wire _11715_;
  wire _11716_;
  wire _11717_;
  wire _11718_;
  wire _11719_;
  wire _11720_;
  wire _11721_;
  wire _11722_;
  wire _11723_;
  wire _11724_;
  wire _11725_;
  wire _11726_;
  wire _11727_;
  wire _11728_;
  wire _11729_;
  wire _11730_;
  wire _11731_;
  wire _11732_;
  wire _11733_;
  wire _11734_;
  wire _11735_;
  wire _11736_;
  wire _11737_;
  wire _11738_;
  wire _11739_;
  wire _11740_;
  wire _11741_;
  wire _11742_;
  wire _11743_;
  wire _11744_;
  wire _11745_;
  wire _11746_;
  wire _11747_;
  wire _11748_;
  wire _11749_;
  wire _11750_;
  wire _11751_;
  wire _11752_;
  wire _11753_;
  wire _11754_;
  wire _11755_;
  wire _11756_;
  wire _11757_;
  wire _11758_;
  wire _11759_;
  wire _11760_;
  wire _11761_;
  wire _11762_;
  wire _11763_;
  wire _11764_;
  wire _11765_;
  wire _11766_;
  wire _11767_;
  wire _11768_;
  wire _11769_;
  wire _11770_;
  wire _11771_;
  wire _11772_;
  wire _11773_;
  wire _11774_;
  wire _11775_;
  wire _11776_;
  wire _11777_;
  wire _11778_;
  wire _11779_;
  wire _11780_;
  wire _11781_;
  wire _11782_;
  wire _11783_;
  wire _11784_;
  wire _11785_;
  wire _11786_;
  wire _11787_;
  wire _11788_;
  wire _11789_;
  wire _11790_;
  wire _11791_;
  wire _11792_;
  wire _11793_;
  wire _11794_;
  wire _11795_;
  wire _11796_;
  wire _11797_;
  wire _11798_;
  wire _11799_;
  wire _11800_;
  wire _11801_;
  wire _11802_;
  wire _11803_;
  wire _11804_;
  wire _11805_;
  wire _11806_;
  wire _11807_;
  wire _11808_;
  wire _11809_;
  wire _11810_;
  wire _11811_;
  wire _11812_;
  wire _11813_;
  wire _11814_;
  wire _11815_;
  wire _11816_;
  wire _11817_;
  wire _11818_;
  wire _11819_;
  wire _11820_;
  wire _11821_;
  wire _11822_;
  wire _11823_;
  wire _11824_;
  wire _11825_;
  wire _11826_;
  wire _11827_;
  wire _11828_;
  wire _11829_;
  wire _11830_;
  wire _11831_;
  wire _11832_;
  wire _11833_;
  wire _11834_;
  wire _11835_;
  wire _11836_;
  wire _11837_;
  wire _11838_;
  wire _11839_;
  wire _11840_;
  wire _11841_;
  wire _11842_;
  wire _11843_;
  wire _11844_;
  wire _11845_;
  wire _11846_;
  wire _11847_;
  wire _11848_;
  wire _11849_;
  wire _11850_;
  wire _11851_;
  wire _11852_;
  wire _11853_;
  wire _11854_;
  wire _11855_;
  wire _11856_;
  wire _11857_;
  wire _11858_;
  wire _11859_;
  wire _11860_;
  wire _11861_;
  wire _11862_;
  wire _11863_;
  wire _11864_;
  wire _11865_;
  wire _11866_;
  wire _11867_;
  wire _11868_;
  wire _11869_;
  wire _11870_;
  wire _11871_;
  wire _11872_;
  wire _11873_;
  wire _11874_;
  wire _11875_;
  wire _11876_;
  wire _11877_;
  wire _11878_;
  wire _11879_;
  wire _11880_;
  wire _11881_;
  wire _11882_;
  wire _11883_;
  wire _11884_;
  wire _11885_;
  wire _11886_;
  wire _11887_;
  wire _11888_;
  wire _11889_;
  wire _11890_;
  wire _11891_;
  wire _11892_;
  wire _11893_;
  wire _11894_;
  wire _11895_;
  wire _11896_;
  wire _11897_;
  wire _11898_;
  wire _11899_;
  wire _11900_;
  wire _11901_;
  wire _11902_;
  wire _11903_;
  wire _11904_;
  wire _11905_;
  wire _11906_;
  wire _11907_;
  wire _11908_;
  wire _11909_;
  wire _11910_;
  wire _11911_;
  wire _11912_;
  wire _11913_;
  wire _11914_;
  wire _11915_;
  wire _11916_;
  wire _11917_;
  wire _11918_;
  wire _11919_;
  wire _11920_;
  wire _11921_;
  wire _11922_;
  wire _11923_;
  wire _11924_;
  wire _11925_;
  wire _11926_;
  wire _11927_;
  wire _11928_;
  wire _11929_;
  wire _11930_;
  wire _11931_;
  wire _11932_;
  wire _11933_;
  wire _11934_;
  wire _11935_;
  wire _11936_;
  wire _11937_;
  wire _11938_;
  wire _11939_;
  wire _11940_;
  wire _11941_;
  wire _11942_;
  wire _11943_;
  wire _11944_;
  wire _11945_;
  wire _11946_;
  wire _11947_;
  wire _11948_;
  wire _11949_;
  wire _11950_;
  wire _11951_;
  wire _11952_;
  wire _11953_;
  wire _11954_;
  wire _11955_;
  wire _11956_;
  wire _11957_;
  wire _11958_;
  wire _11959_;
  wire _11960_;
  wire _11961_;
  wire _11962_;
  wire _11963_;
  wire _11964_;
  wire _11965_;
  wire _11966_;
  wire _11967_;
  wire _11968_;
  wire _11969_;
  wire _11970_;
  wire _11971_;
  wire _11972_;
  wire _11973_;
  wire _11974_;
  wire _11975_;
  wire _11976_;
  wire _11977_;
  wire _11978_;
  wire _11979_;
  wire _11980_;
  wire _11981_;
  wire _11982_;
  wire _11983_;
  wire _11984_;
  wire _11985_;
  wire _11986_;
  wire _11987_;
  wire _11988_;
  wire _11989_;
  wire _11990_;
  wire _11991_;
  wire _11992_;
  wire _11993_;
  wire _11994_;
  wire _11995_;
  wire _11996_;
  wire _11997_;
  wire _11998_;
  wire _11999_;
  wire _12000_;
  wire _12001_;
  wire _12002_;
  wire _12003_;
  wire _12004_;
  wire _12005_;
  wire _12006_;
  wire _12007_;
  wire _12008_;
  wire _12009_;
  wire _12010_;
  wire _12011_;
  wire _12012_;
  wire _12013_;
  wire _12014_;
  wire _12015_;
  wire _12016_;
  wire _12017_;
  wire _12018_;
  wire _12019_;
  wire _12020_;
  wire _12021_;
  wire _12022_;
  wire _12023_;
  wire _12024_;
  wire _12025_;
  wire _12026_;
  wire _12027_;
  wire _12028_;
  wire _12029_;
  wire _12030_;
  wire _12031_;
  wire _12032_;
  wire _12033_;
  wire _12034_;
  wire _12035_;
  wire _12036_;
  wire _12037_;
  wire _12038_;
  wire _12039_;
  wire _12040_;
  wire _12041_;
  wire _12042_;
  wire _12043_;
  wire _12044_;
  wire _12045_;
  wire _12046_;
  wire _12047_;
  wire _12048_;
  wire _12049_;
  wire _12050_;
  wire _12051_;
  wire _12052_;
  wire _12053_;
  wire _12054_;
  wire _12055_;
  wire _12056_;
  wire _12057_;
  wire _12058_;
  wire _12059_;
  wire _12060_;
  wire _12061_;
  wire _12062_;
  wire _12063_;
  wire _12064_;
  wire _12065_;
  wire _12066_;
  wire _12067_;
  wire _12068_;
  wire _12069_;
  wire _12070_;
  wire _12071_;
  wire _12072_;
  wire _12073_;
  wire _12074_;
  wire _12075_;
  wire _12076_;
  wire _12077_;
  wire _12078_;
  wire _12079_;
  wire _12080_;
  wire _12081_;
  wire _12082_;
  wire _12083_;
  wire _12084_;
  wire _12085_;
  wire _12086_;
  wire _12087_;
  wire _12088_;
  wire _12089_;
  wire _12090_;
  wire _12091_;
  wire _12092_;
  wire _12093_;
  wire _12094_;
  wire _12095_;
  wire _12096_;
  wire _12097_;
  wire _12098_;
  wire _12099_;
  wire _12100_;
  wire _12101_;
  wire _12102_;
  wire _12103_;
  wire _12104_;
  wire _12105_;
  wire _12106_;
  wire _12107_;
  wire _12108_;
  wire _12109_;
  wire _12110_;
  wire _12111_;
  wire _12112_;
  wire _12113_;
  wire _12114_;
  wire _12115_;
  wire _12116_;
  wire _12117_;
  wire _12118_;
  wire _12119_;
  wire _12120_;
  wire _12121_;
  wire _12122_;
  wire _12123_;
  wire _12124_;
  wire _12125_;
  wire _12126_;
  wire _12127_;
  wire _12128_;
  wire _12129_;
  wire _12130_;
  wire _12131_;
  wire _12132_;
  wire _12133_;
  wire _12134_;
  wire _12135_;
  wire _12136_;
  wire _12137_;
  wire _12138_;
  wire _12139_;
  wire _12140_;
  wire _12141_;
  wire _12142_;
  wire _12143_;
  wire _12144_;
  wire _12145_;
  wire _12146_;
  wire _12147_;
  wire _12148_;
  wire _12149_;
  wire _12150_;
  wire _12151_;
  wire _12152_;
  wire _12153_;
  wire _12154_;
  wire _12155_;
  wire _12156_;
  wire _12157_;
  wire _12158_;
  wire _12159_;
  wire _12160_;
  wire _12161_;
  wire _12162_;
  wire _12163_;
  wire _12164_;
  wire _12165_;
  wire _12166_;
  wire _12167_;
  wire _12168_;
  wire _12169_;
  wire _12170_;
  wire _12171_;
  wire _12172_;
  wire _12173_;
  wire _12174_;
  wire _12175_;
  wire _12176_;
  wire _12177_;
  wire _12178_;
  wire _12179_;
  wire _12180_;
  wire _12181_;
  wire _12182_;
  wire _12183_;
  wire _12184_;
  wire _12185_;
  wire _12186_;
  wire _12187_;
  wire _12188_;
  wire _12189_;
  wire _12190_;
  wire _12191_;
  wire _12192_;
  wire _12193_;
  wire _12194_;
  wire _12195_;
  wire _12196_;
  wire _12197_;
  wire _12198_;
  wire _12199_;
  wire _12200_;
  wire _12201_;
  wire _12202_;
  wire _12203_;
  wire _12204_;
  wire _12205_;
  wire _12206_;
  wire _12207_;
  wire _12208_;
  wire _12209_;
  wire _12210_;
  wire _12211_;
  wire _12212_;
  wire _12213_;
  wire _12214_;
  wire _12215_;
  wire _12216_;
  wire _12217_;
  wire _12218_;
  wire _12219_;
  wire _12220_;
  wire _12221_;
  wire _12222_;
  wire _12223_;
  wire _12224_;
  wire _12225_;
  wire _12226_;
  wire _12227_;
  wire _12228_;
  wire _12229_;
  wire _12230_;
  wire _12231_;
  wire _12232_;
  wire _12233_;
  wire _12234_;
  wire _12235_;
  wire _12236_;
  wire _12237_;
  wire _12238_;
  wire _12239_;
  wire _12240_;
  wire _12241_;
  wire _12242_;
  wire _12243_;
  wire _12244_;
  wire _12245_;
  wire _12246_;
  wire _12247_;
  wire _12248_;
  wire _12249_;
  wire _12250_;
  wire _12251_;
  wire _12252_;
  wire _12253_;
  wire _12254_;
  wire _12255_;
  wire _12256_;
  wire _12257_;
  wire _12258_;
  wire _12259_;
  wire _12260_;
  wire _12261_;
  wire _12262_;
  wire _12263_;
  wire _12264_;
  wire _12265_;
  wire _12266_;
  wire _12267_;
  wire _12268_;
  wire _12269_;
  wire _12270_;
  wire _12271_;
  wire _12272_;
  wire _12273_;
  wire _12274_;
  wire _12275_;
  wire _12276_;
  wire _12277_;
  wire _12278_;
  wire _12279_;
  wire _12280_;
  wire _12281_;
  wire _12282_;
  wire _12283_;
  wire _12284_;
  wire _12285_;
  wire _12286_;
  wire _12287_;
  wire _12288_;
  wire _12289_;
  wire _12290_;
  wire _12291_;
  wire _12292_;
  wire _12293_;
  wire _12294_;
  wire _12295_;
  wire _12296_;
  wire _12297_;
  wire _12298_;
  wire _12299_;
  wire _12300_;
  wire _12301_;
  wire _12302_;
  wire _12303_;
  wire _12304_;
  wire _12305_;
  wire _12306_;
  wire _12307_;
  wire _12308_;
  wire _12309_;
  wire _12310_;
  wire _12311_;
  wire _12312_;
  wire _12313_;
  wire _12314_;
  wire _12315_;
  wire _12316_;
  wire _12317_;
  wire _12318_;
  wire _12319_;
  wire _12320_;
  wire _12321_;
  wire _12322_;
  wire _12323_;
  wire _12324_;
  wire _12325_;
  wire _12326_;
  wire _12327_;
  wire _12328_;
  wire _12329_;
  wire _12330_;
  wire _12331_;
  wire _12332_;
  wire _12333_;
  wire _12334_;
  wire _12335_;
  wire _12336_;
  wire _12337_;
  wire _12338_;
  wire _12339_;
  wire _12340_;
  wire _12341_;
  wire _12342_;
  wire _12343_;
  wire _12344_;
  wire _12345_;
  wire _12346_;
  wire _12347_;
  wire _12348_;
  wire _12349_;
  wire _12350_;
  wire _12351_;
  wire _12352_;
  wire _12353_;
  wire _12354_;
  wire _12355_;
  wire _12356_;
  wire _12357_;
  wire _12358_;
  wire _12359_;
  wire _12360_;
  wire _12361_;
  wire _12362_;
  wire _12363_;
  wire _12364_;
  wire _12365_;
  wire _12366_;
  wire _12367_;
  wire _12368_;
  wire _12369_;
  wire _12370_;
  wire _12371_;
  wire _12372_;
  wire _12373_;
  wire _12374_;
  wire _12375_;
  wire _12376_;
  wire _12377_;
  wire _12378_;
  wire _12379_;
  wire _12380_;
  wire _12381_;
  wire _12382_;
  wire _12383_;
  wire _12384_;
  wire _12385_;
  wire _12386_;
  wire _12387_;
  wire _12388_;
  wire _12389_;
  wire _12390_;
  wire _12391_;
  wire _12392_;
  wire _12393_;
  wire _12394_;
  wire _12395_;
  wire _12396_;
  wire _12397_;
  wire _12398_;
  wire _12399_;
  wire _12400_;
  wire _12401_;
  wire _12402_;
  wire _12403_;
  wire _12404_;
  wire _12405_;
  wire _12406_;
  wire _12407_;
  wire _12408_;
  wire _12409_;
  wire _12410_;
  wire _12411_;
  wire _12412_;
  wire _12413_;
  wire _12414_;
  wire _12415_;
  wire _12416_;
  wire _12417_;
  wire _12418_;
  wire _12419_;
  wire _12420_;
  wire _12421_;
  wire _12422_;
  wire _12423_;
  wire _12424_;
  wire _12425_;
  wire _12426_;
  wire _12427_;
  wire _12428_;
  wire _12429_;
  wire _12430_;
  wire _12431_;
  wire _12432_;
  wire _12433_;
  wire _12434_;
  wire _12435_;
  wire _12436_;
  wire _12437_;
  wire _12438_;
  wire _12439_;
  wire _12440_;
  wire _12441_;
  wire _12442_;
  wire _12443_;
  wire _12444_;
  wire _12445_;
  wire _12446_;
  wire _12447_;
  wire _12448_;
  wire _12449_;
  wire _12450_;
  wire _12451_;
  wire _12452_;
  wire _12453_;
  wire _12454_;
  wire _12455_;
  wire _12456_;
  wire _12457_;
  wire _12458_;
  wire _12459_;
  wire _12460_;
  wire _12461_;
  wire _12462_;
  wire _12463_;
  wire _12464_;
  wire _12465_;
  wire _12466_;
  wire _12467_;
  wire _12468_;
  wire _12469_;
  wire _12470_;
  wire _12471_;
  wire _12472_;
  wire _12473_;
  wire _12474_;
  wire _12475_;
  wire _12476_;
  wire _12477_;
  wire _12478_;
  wire _12479_;
  wire _12480_;
  wire _12481_;
  wire _12482_;
  wire _12483_;
  wire _12484_;
  wire _12485_;
  wire _12486_;
  wire _12487_;
  wire _12488_;
  wire _12489_;
  wire _12490_;
  wire _12491_;
  wire _12492_;
  wire _12493_;
  wire _12494_;
  wire _12495_;
  wire _12496_;
  wire _12497_;
  wire _12498_;
  wire _12499_;
  wire _12500_;
  wire _12501_;
  wire _12502_;
  wire _12503_;
  wire _12504_;
  wire _12505_;
  wire _12506_;
  wire _12507_;
  wire _12508_;
  wire _12509_;
  wire _12510_;
  wire _12511_;
  wire _12512_;
  wire _12513_;
  wire _12514_;
  wire _12515_;
  wire _12516_;
  wire _12517_;
  wire _12518_;
  wire _12519_;
  wire _12520_;
  wire _12521_;
  wire _12522_;
  wire _12523_;
  wire _12524_;
  wire _12525_;
  wire _12526_;
  wire _12527_;
  wire _12528_;
  wire _12529_;
  wire _12530_;
  wire _12531_;
  wire _12532_;
  wire _12533_;
  wire _12534_;
  wire _12535_;
  wire _12536_;
  wire _12537_;
  wire _12538_;
  wire _12539_;
  wire _12540_;
  wire _12541_;
  wire _12542_;
  wire _12543_;
  wire _12544_;
  wire _12545_;
  wire _12546_;
  wire _12547_;
  wire _12548_;
  wire _12549_;
  wire _12550_;
  wire _12551_;
  wire _12552_;
  wire _12553_;
  wire _12554_;
  wire _12555_;
  wire _12556_;
  wire _12557_;
  wire _12558_;
  wire _12559_;
  wire _12560_;
  wire _12561_;
  wire _12562_;
  wire _12563_;
  wire _12564_;
  wire _12565_;
  wire _12566_;
  wire _12567_;
  wire _12568_;
  wire _12569_;
  wire _12570_;
  wire _12571_;
  wire _12572_;
  wire _12573_;
  wire _12574_;
  wire _12575_;
  wire _12576_;
  wire _12577_;
  wire _12578_;
  wire _12579_;
  wire _12580_;
  wire _12581_;
  wire _12582_;
  wire _12583_;
  wire _12584_;
  wire _12585_;
  wire _12586_;
  wire _12587_;
  wire _12588_;
  wire _12589_;
  wire _12590_;
  wire _12591_;
  wire _12592_;
  wire _12593_;
  wire _12594_;
  wire _12595_;
  wire _12596_;
  wire _12597_;
  wire _12598_;
  wire _12599_;
  wire _12600_;
  wire _12601_;
  wire _12602_;
  wire _12603_;
  wire _12604_;
  wire _12605_;
  wire _12606_;
  wire _12607_;
  wire _12608_;
  wire _12609_;
  wire _12610_;
  wire _12611_;
  wire _12612_;
  wire _12613_;
  wire _12614_;
  wire _12615_;
  wire _12616_;
  wire _12617_;
  wire _12618_;
  wire _12619_;
  wire _12620_;
  wire _12621_;
  wire _12622_;
  wire _12623_;
  wire _12624_;
  wire _12625_;
  wire _12626_;
  wire _12627_;
  wire _12628_;
  wire _12629_;
  wire _12630_;
  wire _12631_;
  wire _12632_;
  wire _12633_;
  wire _12634_;
  wire _12635_;
  wire _12636_;
  wire _12637_;
  wire _12638_;
  wire _12639_;
  wire _12640_;
  wire _12641_;
  wire _12642_;
  wire _12643_;
  wire _12644_;
  wire _12645_;
  wire _12646_;
  wire _12647_;
  wire _12648_;
  wire _12649_;
  wire _12650_;
  wire _12651_;
  wire _12652_;
  wire _12653_;
  wire _12654_;
  wire _12655_;
  wire _12656_;
  wire _12657_;
  wire _12658_;
  wire _12659_;
  wire _12660_;
  wire _12661_;
  wire _12662_;
  wire _12663_;
  wire _12664_;
  wire _12665_;
  wire _12666_;
  wire _12667_;
  wire _12668_;
  wire _12669_;
  wire _12670_;
  wire _12671_;
  wire _12672_;
  wire _12673_;
  wire _12674_;
  wire _12675_;
  wire _12676_;
  wire _12677_;
  wire _12678_;
  wire _12679_;
  wire _12680_;
  wire _12681_;
  wire _12682_;
  wire _12683_;
  wire _12684_;
  wire _12685_;
  wire _12686_;
  wire _12687_;
  wire _12688_;
  wire _12689_;
  wire _12690_;
  wire _12691_;
  wire _12692_;
  wire _12693_;
  wire _12694_;
  wire _12695_;
  wire _12696_;
  wire _12697_;
  wire _12698_;
  wire _12699_;
  wire _12700_;
  wire _12701_;
  wire _12702_;
  wire _12703_;
  wire _12704_;
  wire _12705_;
  wire _12706_;
  wire _12707_;
  wire _12708_;
  wire _12709_;
  wire _12710_;
  wire _12711_;
  wire _12712_;
  wire _12713_;
  wire _12714_;
  wire _12715_;
  wire _12716_;
  wire _12717_;
  wire _12718_;
  wire _12719_;
  wire _12720_;
  wire _12721_;
  wire _12722_;
  wire _12723_;
  wire _12724_;
  wire _12725_;
  wire _12726_;
  wire _12727_;
  wire _12728_;
  wire _12729_;
  wire _12730_;
  wire _12731_;
  wire _12732_;
  wire _12733_;
  wire _12734_;
  wire _12735_;
  wire _12736_;
  wire _12737_;
  wire _12738_;
  wire _12739_;
  wire _12740_;
  wire _12741_;
  wire _12742_;
  wire _12743_;
  wire _12744_;
  wire _12745_;
  wire _12746_;
  wire _12747_;
  wire _12748_;
  wire _12749_;
  wire _12750_;
  wire _12751_;
  wire _12752_;
  wire _12753_;
  wire _12754_;
  wire _12755_;
  wire _12756_;
  wire _12757_;
  wire _12758_;
  wire _12759_;
  wire _12760_;
  wire _12761_;
  wire _12762_;
  wire _12763_;
  wire _12764_;
  wire _12765_;
  wire _12766_;
  wire _12767_;
  wire _12768_;
  wire _12769_;
  wire _12770_;
  wire _12771_;
  wire _12772_;
  wire _12773_;
  wire _12774_;
  wire _12775_;
  wire _12776_;
  wire _12777_;
  wire _12778_;
  wire _12779_;
  wire _12780_;
  wire _12781_;
  wire _12782_;
  wire _12783_;
  wire _12784_;
  wire _12785_;
  wire _12786_;
  wire _12787_;
  wire _12788_;
  wire _12789_;
  wire _12790_;
  wire _12791_;
  wire _12792_;
  wire _12793_;
  wire _12794_;
  wire _12795_;
  wire _12796_;
  wire _12797_;
  wire _12798_;
  wire _12799_;
  wire _12800_;
  wire _12801_;
  wire _12802_;
  wire _12803_;
  wire _12804_;
  wire _12805_;
  wire _12806_;
  wire _12807_;
  wire _12808_;
  wire _12809_;
  wire _12810_;
  wire _12811_;
  wire _12812_;
  wire _12813_;
  wire _12814_;
  wire _12815_;
  wire _12816_;
  wire _12817_;
  wire _12818_;
  wire _12819_;
  wire _12820_;
  wire _12821_;
  wire _12822_;
  wire _12823_;
  wire _12824_;
  wire _12825_;
  wire _12826_;
  wire _12827_;
  wire _12828_;
  wire _12829_;
  wire _12830_;
  wire _12831_;
  wire _12832_;
  wire _12833_;
  wire _12834_;
  wire _12835_;
  wire _12836_;
  wire _12837_;
  wire _12838_;
  wire _12839_;
  wire _12840_;
  wire _12841_;
  wire _12842_;
  wire _12843_;
  wire _12844_;
  wire _12845_;
  wire _12846_;
  wire _12847_;
  wire _12848_;
  wire _12849_;
  wire _12850_;
  wire _12851_;
  wire _12852_;
  wire _12853_;
  wire _12854_;
  wire _12855_;
  wire _12856_;
  wire _12857_;
  wire _12858_;
  wire _12859_;
  wire _12860_;
  wire _12861_;
  wire _12862_;
  wire _12863_;
  wire _12864_;
  wire _12865_;
  wire _12866_;
  wire _12867_;
  wire _12868_;
  wire _12869_;
  wire _12870_;
  wire _12871_;
  wire _12872_;
  wire _12873_;
  wire _12874_;
  wire _12875_;
  wire _12876_;
  wire _12877_;
  wire _12878_;
  wire _12879_;
  wire _12880_;
  wire _12881_;
  wire _12882_;
  wire _12883_;
  wire _12884_;
  wire _12885_;
  wire _12886_;
  wire _12887_;
  wire _12888_;
  wire _12889_;
  wire _12890_;
  wire _12891_;
  wire _12892_;
  wire _12893_;
  wire _12894_;
  wire _12895_;
  wire _12896_;
  wire _12897_;
  wire _12898_;
  wire _12899_;
  wire _12900_;
  wire _12901_;
  wire _12902_;
  wire _12903_;
  wire _12904_;
  wire _12905_;
  wire _12906_;
  wire _12907_;
  wire _12908_;
  wire _12909_;
  wire _12910_;
  wire _12911_;
  wire _12912_;
  wire _12913_;
  wire _12914_;
  wire _12915_;
  wire _12916_;
  wire _12917_;
  wire _12918_;
  wire _12919_;
  wire _12920_;
  wire _12921_;
  wire _12922_;
  wire _12923_;
  wire _12924_;
  wire _12925_;
  wire _12926_;
  wire _12927_;
  wire _12928_;
  wire _12929_;
  wire _12930_;
  wire _12931_;
  wire _12932_;
  wire _12933_;
  wire _12934_;
  wire _12935_;
  wire _12936_;
  wire _12937_;
  wire _12938_;
  wire _12939_;
  wire _12940_;
  wire _12941_;
  wire _12942_;
  wire _12943_;
  wire _12944_;
  wire _12945_;
  wire _12946_;
  wire _12947_;
  wire _12948_;
  wire _12949_;
  wire _12950_;
  wire _12951_;
  wire _12952_;
  wire _12953_;
  wire _12954_;
  wire _12955_;
  wire _12956_;
  wire _12957_;
  wire _12958_;
  wire _12959_;
  wire _12960_;
  wire _12961_;
  wire _12962_;
  wire _12963_;
  wire _12964_;
  wire _12965_;
  wire _12966_;
  wire _12967_;
  wire _12968_;
  wire _12969_;
  wire _12970_;
  wire _12971_;
  wire _12972_;
  wire _12973_;
  wire _12974_;
  wire _12975_;
  wire _12976_;
  wire _12977_;
  wire _12978_;
  wire _12979_;
  wire _12980_;
  wire _12981_;
  wire _12982_;
  wire _12983_;
  wire _12984_;
  wire _12985_;
  wire _12986_;
  wire _12987_;
  wire _12988_;
  wire _12989_;
  wire _12990_;
  wire _12991_;
  wire _12992_;
  wire _12993_;
  wire _12994_;
  wire _12995_;
  wire _12996_;
  wire _12997_;
  wire _12998_;
  wire _12999_;
  wire _13000_;
  wire _13001_;
  wire _13002_;
  wire _13003_;
  wire _13004_;
  wire _13005_;
  wire _13006_;
  wire _13007_;
  wire _13008_;
  wire _13009_;
  wire _13010_;
  wire _13011_;
  wire _13012_;
  wire _13013_;
  wire _13014_;
  wire _13015_;
  wire _13016_;
  wire _13017_;
  wire _13018_;
  wire _13019_;
  wire _13020_;
  wire _13021_;
  wire _13022_;
  wire _13023_;
  wire _13024_;
  wire _13025_;
  wire _13026_;
  wire _13027_;
  wire _13028_;
  wire _13029_;
  wire _13030_;
  wire _13031_;
  wire _13032_;
  wire _13033_;
  wire _13034_;
  wire _13035_;
  wire _13036_;
  wire _13037_;
  wire _13038_;
  wire _13039_;
  wire _13040_;
  wire _13041_;
  wire _13042_;
  wire _13043_;
  wire _13044_;
  wire _13045_;
  wire _13046_;
  wire _13047_;
  wire _13048_;
  wire _13049_;
  wire _13050_;
  wire _13051_;
  wire _13052_;
  wire _13053_;
  wire _13054_;
  wire _13055_;
  wire _13056_;
  wire _13057_;
  wire _13058_;
  wire _13059_;
  wire _13060_;
  wire _13061_;
  wire _13062_;
  wire _13063_;
  wire _13064_;
  wire _13065_;
  wire _13066_;
  wire _13067_;
  wire _13068_;
  wire _13069_;
  wire _13070_;
  wire _13071_;
  wire _13072_;
  wire _13073_;
  wire _13074_;
  wire _13075_;
  wire _13076_;
  wire _13077_;
  wire _13078_;
  wire _13079_;
  wire _13080_;
  wire _13081_;
  wire _13082_;
  wire _13083_;
  wire _13084_;
  wire _13085_;
  wire _13086_;
  wire _13087_;
  wire _13088_;
  wire _13089_;
  wire _13090_;
  wire _13091_;
  wire _13092_;
  wire _13093_;
  wire _13094_;
  wire _13095_;
  wire _13096_;
  wire _13097_;
  wire _13098_;
  wire _13099_;
  wire _13100_;
  wire _13101_;
  wire _13102_;
  wire _13103_;
  wire _13104_;
  wire _13105_;
  wire _13106_;
  wire _13107_;
  wire _13108_;
  wire _13109_;
  wire _13110_;
  wire _13111_;
  wire _13112_;
  wire _13113_;
  wire _13114_;
  wire _13115_;
  wire _13116_;
  wire _13117_;
  wire _13118_;
  wire _13119_;
  wire _13120_;
  wire _13121_;
  wire _13122_;
  wire _13123_;
  wire _13124_;
  wire _13125_;
  wire _13126_;
  wire _13127_;
  wire _13128_;
  wire _13129_;
  wire _13130_;
  wire _13131_;
  wire _13132_;
  wire _13133_;
  wire _13134_;
  wire _13135_;
  wire _13136_;
  wire _13137_;
  wire _13138_;
  wire _13139_;
  wire _13140_;
  wire _13141_;
  wire _13142_;
  wire _13143_;
  wire _13144_;
  wire _13145_;
  wire _13146_;
  wire _13147_;
  wire _13148_;
  wire _13149_;
  wire _13150_;
  wire _13151_;
  wire _13152_;
  wire _13153_;
  wire _13154_;
  wire _13155_;
  wire _13156_;
  wire _13157_;
  wire _13158_;
  wire _13159_;
  wire _13160_;
  wire _13161_;
  wire _13162_;
  wire _13163_;
  wire _13164_;
  wire _13165_;
  wire _13166_;
  wire _13167_;
  wire _13168_;
  wire _13169_;
  wire _13170_;
  wire _13171_;
  wire _13172_;
  wire _13173_;
  wire _13174_;
  wire _13175_;
  wire _13176_;
  wire _13177_;
  wire _13178_;
  wire _13179_;
  wire _13180_;
  wire _13181_;
  wire _13182_;
  wire _13183_;
  wire _13184_;
  wire _13185_;
  wire _13186_;
  wire _13187_;
  wire _13188_;
  wire _13189_;
  wire _13190_;
  wire _13191_;
  wire _13192_;
  wire _13193_;
  wire _13194_;
  wire _13195_;
  wire _13196_;
  wire _13197_;
  wire _13198_;
  wire _13199_;
  wire _13200_;
  wire _13201_;
  wire _13202_;
  wire _13203_;
  wire _13204_;
  wire _13205_;
  wire _13206_;
  wire _13207_;
  wire _13208_;
  wire _13209_;
  wire _13210_;
  wire _13211_;
  wire _13212_;
  wire _13213_;
  wire _13214_;
  wire _13215_;
  wire _13216_;
  wire _13217_;
  wire _13218_;
  wire _13219_;
  wire _13220_;
  wire _13221_;
  wire _13222_;
  wire _13223_;
  wire _13224_;
  wire _13225_;
  wire _13226_;
  wire _13227_;
  wire _13228_;
  wire _13229_;
  wire _13230_;
  wire _13231_;
  wire _13232_;
  wire _13233_;
  wire _13234_;
  wire _13235_;
  wire _13236_;
  wire _13237_;
  wire _13238_;
  wire _13239_;
  wire _13240_;
  wire _13241_;
  wire _13242_;
  wire _13243_;
  wire _13244_;
  wire _13245_;
  wire _13246_;
  wire _13247_;
  wire _13248_;
  wire _13249_;
  wire _13250_;
  wire _13251_;
  wire _13252_;
  wire _13253_;
  wire _13254_;
  wire _13255_;
  wire _13256_;
  wire _13257_;
  wire _13258_;
  wire _13259_;
  wire _13260_;
  wire _13261_;
  wire _13262_;
  wire _13263_;
  wire _13264_;
  wire _13265_;
  wire _13266_;
  wire _13267_;
  wire _13268_;
  wire _13269_;
  wire _13270_;
  wire _13271_;
  wire _13272_;
  wire _13273_;
  wire _13274_;
  wire _13275_;
  wire _13276_;
  wire _13277_;
  wire _13278_;
  wire _13279_;
  wire _13280_;
  wire _13281_;
  wire _13282_;
  wire _13283_;
  wire _13284_;
  wire _13285_;
  wire _13286_;
  wire _13287_;
  wire _13288_;
  wire _13289_;
  wire _13290_;
  wire _13291_;
  wire _13292_;
  wire _13293_;
  wire _13294_;
  wire _13295_;
  wire _13296_;
  wire _13297_;
  wire _13298_;
  wire _13299_;
  wire _13300_;
  wire _13301_;
  wire _13302_;
  wire _13303_;
  wire _13304_;
  wire _13305_;
  wire _13306_;
  wire _13307_;
  wire _13308_;
  wire _13309_;
  wire _13310_;
  wire _13311_;
  wire _13312_;
  wire _13313_;
  wire _13314_;
  wire _13315_;
  wire _13316_;
  wire _13317_;
  wire _13318_;
  wire _13319_;
  wire _13320_;
  wire _13321_;
  wire _13322_;
  wire _13323_;
  wire _13324_;
  wire _13325_;
  wire _13326_;
  wire _13327_;
  wire _13328_;
  wire _13329_;
  wire _13330_;
  wire _13331_;
  wire _13332_;
  wire _13333_;
  wire _13334_;
  wire _13335_;
  wire _13336_;
  wire _13337_;
  wire _13338_;
  wire _13339_;
  wire _13340_;
  wire _13341_;
  wire _13342_;
  wire _13343_;
  wire _13344_;
  wire _13345_;
  wire _13346_;
  wire _13347_;
  wire _13348_;
  wire _13349_;
  wire _13350_;
  wire _13351_;
  wire _13352_;
  wire _13353_;
  wire _13354_;
  wire _13355_;
  wire _13356_;
  wire _13357_;
  wire _13358_;
  wire _13359_;
  wire _13360_;
  wire _13361_;
  wire _13362_;
  wire _13363_;
  wire _13364_;
  wire _13365_;
  wire _13366_;
  wire _13367_;
  wire _13368_;
  wire _13369_;
  wire _13370_;
  wire _13371_;
  wire _13372_;
  wire _13373_;
  wire _13374_;
  wire _13375_;
  wire _13376_;
  wire _13377_;
  wire _13378_;
  wire _13379_;
  wire _13380_;
  wire _13381_;
  wire _13382_;
  wire _13383_;
  wire _13384_;
  wire _13385_;
  wire _13386_;
  wire _13387_;
  wire _13388_;
  wire _13389_;
  wire _13390_;
  wire _13391_;
  wire _13392_;
  wire _13393_;
  wire _13394_;
  wire _13395_;
  wire _13396_;
  wire _13397_;
  wire _13398_;
  wire _13399_;
  wire _13400_;
  wire _13401_;
  wire _13402_;
  wire _13403_;
  wire _13404_;
  wire _13405_;
  wire _13406_;
  wire _13407_;
  wire _13408_;
  wire _13409_;
  wire _13410_;
  wire _13411_;
  wire _13412_;
  wire _13413_;
  wire _13414_;
  wire _13415_;
  wire _13416_;
  wire _13417_;
  wire _13418_;
  wire _13419_;
  wire _13420_;
  wire _13421_;
  wire _13422_;
  wire _13423_;
  wire _13424_;
  wire _13425_;
  wire _13426_;
  wire _13427_;
  wire _13428_;
  wire _13429_;
  wire _13430_;
  wire _13431_;
  wire _13432_;
  wire _13433_;
  wire _13434_;
  wire _13435_;
  wire _13436_;
  wire _13437_;
  wire _13438_;
  wire _13439_;
  wire _13440_;
  wire _13441_;
  wire _13442_;
  wire _13443_;
  wire _13444_;
  wire _13445_;
  wire _13446_;
  wire _13447_;
  wire _13448_;
  wire _13449_;
  wire _13450_;
  wire _13451_;
  wire _13452_;
  wire _13453_;
  wire _13454_;
  wire _13455_;
  wire _13456_;
  wire _13457_;
  wire _13458_;
  wire _13459_;
  wire _13460_;
  wire _13461_;
  wire _13462_;
  wire _13463_;
  wire _13464_;
  wire _13465_;
  wire _13466_;
  wire _13467_;
  wire _13468_;
  wire _13469_;
  wire _13470_;
  wire _13471_;
  wire _13472_;
  wire _13473_;
  wire _13474_;
  wire _13475_;
  wire _13476_;
  wire _13477_;
  wire _13478_;
  wire _13479_;
  wire _13480_;
  wire _13481_;
  wire _13482_;
  wire _13483_;
  wire _13484_;
  wire _13485_;
  wire _13486_;
  wire _13487_;
  wire _13488_;
  wire _13489_;
  wire _13490_;
  wire _13491_;
  wire _13492_;
  wire _13493_;
  wire _13494_;
  wire _13495_;
  wire _13496_;
  wire _13497_;
  wire _13498_;
  wire _13499_;
  wire _13500_;
  wire _13501_;
  wire _13502_;
  wire _13503_;
  wire _13504_;
  wire _13505_;
  wire _13506_;
  wire _13507_;
  wire _13508_;
  wire _13509_;
  wire _13510_;
  wire _13511_;
  wire _13512_;
  wire _13513_;
  wire _13514_;
  wire _13515_;
  wire _13516_;
  wire _13517_;
  wire _13518_;
  wire _13519_;
  wire _13520_;
  wire _13521_;
  wire _13522_;
  wire _13523_;
  wire _13524_;
  wire _13525_;
  wire _13526_;
  wire _13527_;
  wire _13528_;
  wire _13529_;
  wire _13530_;
  wire _13531_;
  wire _13532_;
  wire _13533_;
  wire _13534_;
  wire _13535_;
  wire _13536_;
  wire _13537_;
  wire _13538_;
  wire _13539_;
  wire _13540_;
  wire _13541_;
  wire _13542_;
  wire _13543_;
  wire _13544_;
  wire _13545_;
  wire _13546_;
  wire _13547_;
  wire _13548_;
  wire _13549_;
  wire _13550_;
  wire _13551_;
  wire _13552_;
  wire _13553_;
  wire _13554_;
  wire _13555_;
  wire _13556_;
  wire _13557_;
  wire _13558_;
  wire _13559_;
  wire _13560_;
  wire _13561_;
  wire _13562_;
  wire _13563_;
  wire _13564_;
  wire _13565_;
  wire _13566_;
  wire _13567_;
  wire _13568_;
  wire _13569_;
  wire _13570_;
  wire _13571_;
  wire _13572_;
  wire _13573_;
  wire _13574_;
  wire _13575_;
  wire _13576_;
  wire _13577_;
  wire _13578_;
  wire _13579_;
  wire _13580_;
  wire _13581_;
  wire _13582_;
  wire _13583_;
  wire _13584_;
  wire _13585_;
  wire _13586_;
  wire _13587_;
  wire _13588_;
  wire _13589_;
  wire _13590_;
  wire _13591_;
  wire _13592_;
  wire _13593_;
  wire _13594_;
  wire _13595_;
  wire _13596_;
  wire _13597_;
  wire _13598_;
  wire _13599_;
  wire _13600_;
  wire _13601_;
  wire _13602_;
  wire _13603_;
  wire _13604_;
  wire _13605_;
  wire _13606_;
  wire _13607_;
  wire _13608_;
  wire _13609_;
  wire _13610_;
  wire _13611_;
  wire _13612_;
  wire _13613_;
  wire _13614_;
  wire _13615_;
  wire _13616_;
  wire _13617_;
  wire _13618_;
  wire _13619_;
  wire _13620_;
  wire _13621_;
  wire _13622_;
  wire _13623_;
  wire _13624_;
  wire _13625_;
  wire _13626_;
  wire _13627_;
  wire _13628_;
  wire _13629_;
  wire _13630_;
  wire _13631_;
  wire _13632_;
  wire _13633_;
  wire _13634_;
  wire _13635_;
  wire _13636_;
  wire _13637_;
  wire _13638_;
  wire _13639_;
  wire _13640_;
  wire _13641_;
  wire _13642_;
  wire _13643_;
  wire _13644_;
  wire _13645_;
  wire _13646_;
  wire _13647_;
  wire _13648_;
  wire _13649_;
  wire _13650_;
  wire _13651_;
  wire _13652_;
  wire _13653_;
  wire _13654_;
  wire _13655_;
  wire _13656_;
  wire _13657_;
  wire _13658_;
  wire _13659_;
  wire _13660_;
  wire _13661_;
  wire _13662_;
  wire _13663_;
  wire _13664_;
  wire _13665_;
  wire _13666_;
  wire _13667_;
  wire _13668_;
  wire _13669_;
  wire _13670_;
  wire _13671_;
  wire _13672_;
  wire _13673_;
  wire _13674_;
  wire _13675_;
  wire _13676_;
  wire _13677_;
  wire _13678_;
  wire _13679_;
  wire _13680_;
  wire _13681_;
  wire _13682_;
  wire _13683_;
  wire _13684_;
  wire _13685_;
  wire _13686_;
  wire _13687_;
  wire _13688_;
  wire _13689_;
  wire _13690_;
  wire _13691_;
  wire _13692_;
  wire _13693_;
  wire _13694_;
  wire _13695_;
  wire _13696_;
  wire _13697_;
  wire _13698_;
  wire _13699_;
  wire _13700_;
  wire _13701_;
  wire _13702_;
  wire _13703_;
  wire _13704_;
  wire _13705_;
  wire _13706_;
  wire _13707_;
  wire _13708_;
  wire _13709_;
  wire _13710_;
  wire _13711_;
  wire _13712_;
  wire _13713_;
  wire _13714_;
  wire _13715_;
  wire _13716_;
  wire _13717_;
  wire _13718_;
  wire _13719_;
  wire _13720_;
  wire _13721_;
  wire _13722_;
  wire _13723_;
  wire _13724_;
  wire _13725_;
  wire _13726_;
  wire _13727_;
  wire _13728_;
  wire _13729_;
  wire _13730_;
  wire _13731_;
  wire _13732_;
  wire _13733_;
  wire _13734_;
  wire _13735_;
  wire _13736_;
  wire _13737_;
  wire _13738_;
  wire _13739_;
  wire _13740_;
  wire _13741_;
  wire _13742_;
  wire _13743_;
  wire _13744_;
  wire _13745_;
  wire _13746_;
  wire _13747_;
  wire _13748_;
  wire _13749_;
  wire _13750_;
  wire _13751_;
  wire _13752_;
  wire _13753_;
  wire _13754_;
  wire _13755_;
  wire _13756_;
  wire _13757_;
  wire _13758_;
  wire _13759_;
  wire _13760_;
  wire _13761_;
  wire _13762_;
  wire _13763_;
  wire _13764_;
  wire _13765_;
  wire _13766_;
  wire _13767_;
  wire _13768_;
  wire _13769_;
  wire _13770_;
  wire _13771_;
  wire _13772_;
  wire _13773_;
  wire _13774_;
  wire _13775_;
  wire _13776_;
  wire _13777_;
  wire _13778_;
  wire _13779_;
  wire _13780_;
  wire _13781_;
  wire _13782_;
  wire _13783_;
  wire _13784_;
  wire _13785_;
  wire _13786_;
  wire _13787_;
  wire _13788_;
  wire _13789_;
  wire _13790_;
  wire _13791_;
  wire _13792_;
  wire _13793_;
  wire _13794_;
  wire _13795_;
  wire _13796_;
  wire _13797_;
  wire _13798_;
  wire _13799_;
  wire _13800_;
  wire _13801_;
  wire _13802_;
  wire _13803_;
  wire _13804_;
  wire _13805_;
  wire _13806_;
  wire _13807_;
  wire _13808_;
  wire _13809_;
  wire _13810_;
  wire _13811_;
  wire _13812_;
  wire _13813_;
  wire _13814_;
  wire _13815_;
  wire _13816_;
  wire _13817_;
  wire _13818_;
  wire _13819_;
  wire _13820_;
  wire _13821_;
  wire _13822_;
  wire _13823_;
  wire _13824_;
  wire _13825_;
  wire _13826_;
  wire _13827_;
  wire _13828_;
  wire _13829_;
  wire _13830_;
  wire _13831_;
  wire _13832_;
  wire _13833_;
  wire _13834_;
  wire _13835_;
  wire _13836_;
  wire _13837_;
  wire _13838_;
  wire _13839_;
  wire _13840_;
  wire _13841_;
  wire _13842_;
  wire _13843_;
  wire _13844_;
  wire _13845_;
  wire _13846_;
  wire _13847_;
  wire _13848_;
  wire _13849_;
  wire _13850_;
  wire _13851_;
  wire _13852_;
  wire _13853_;
  wire _13854_;
  wire _13855_;
  wire _13856_;
  wire _13857_;
  wire _13858_;
  wire _13859_;
  wire _13860_;
  wire _13861_;
  wire _13862_;
  wire _13863_;
  wire _13864_;
  wire _13865_;
  wire _13866_;
  wire _13867_;
  wire _13868_;
  wire _13869_;
  wire _13870_;
  wire _13871_;
  wire _13872_;
  wire _13873_;
  wire _13874_;
  wire _13875_;
  wire _13876_;
  wire _13877_;
  wire _13878_;
  wire _13879_;
  wire _13880_;
  wire _13881_;
  wire _13882_;
  wire _13883_;
  wire _13884_;
  wire _13885_;
  wire _13886_;
  wire _13887_;
  wire _13888_;
  wire _13889_;
  wire _13890_;
  wire _13891_;
  wire _13892_;
  wire _13893_;
  wire _13894_;
  wire _13895_;
  wire _13896_;
  wire _13897_;
  wire _13898_;
  wire _13899_;
  wire _13900_;
  wire _13901_;
  wire _13902_;
  wire _13903_;
  wire _13904_;
  wire _13905_;
  wire _13906_;
  wire _13907_;
  wire _13908_;
  wire _13909_;
  wire _13910_;
  wire _13911_;
  wire _13912_;
  wire _13913_;
  wire _13914_;
  wire _13915_;
  wire _13916_;
  wire _13917_;
  wire _13918_;
  wire _13919_;
  wire _13920_;
  wire _13921_;
  wire _13922_;
  wire _13923_;
  wire _13924_;
  wire _13925_;
  wire _13926_;
  wire _13927_;
  wire _13928_;
  wire _13929_;
  wire _13930_;
  wire _13931_;
  wire _13932_;
  wire _13933_;
  wire _13934_;
  wire _13935_;
  wire _13936_;
  wire _13937_;
  wire _13938_;
  wire _13939_;
  wire _13940_;
  wire _13941_;
  wire _13942_;
  wire _13943_;
  wire _13944_;
  wire _13945_;
  wire _13946_;
  wire _13947_;
  wire _13948_;
  wire _13949_;
  wire _13950_;
  wire _13951_;
  wire _13952_;
  wire _13953_;
  wire _13954_;
  wire _13955_;
  wire _13956_;
  wire _13957_;
  wire _13958_;
  wire _13959_;
  wire _13960_;
  wire _13961_;
  wire _13962_;
  wire _13963_;
  wire _13964_;
  wire _13965_;
  wire _13966_;
  wire _13967_;
  wire _13968_;
  wire _13969_;
  wire _13970_;
  wire _13971_;
  wire _13972_;
  wire _13973_;
  wire _13974_;
  wire _13975_;
  wire _13976_;
  wire _13977_;
  wire _13978_;
  wire _13979_;
  wire _13980_;
  wire _13981_;
  wire _13982_;
  wire _13983_;
  wire _13984_;
  wire _13985_;
  wire _13986_;
  wire _13987_;
  wire _13988_;
  wire _13989_;
  wire _13990_;
  wire _13991_;
  wire _13992_;
  wire _13993_;
  wire _13994_;
  wire _13995_;
  wire _13996_;
  wire _13997_;
  wire _13998_;
  wire _13999_;
  wire _14000_;
  wire _14001_;
  wire _14002_;
  wire _14003_;
  wire _14004_;
  wire _14005_;
  wire _14006_;
  wire _14007_;
  wire _14008_;
  wire _14009_;
  wire _14010_;
  wire _14011_;
  wire _14012_;
  wire _14013_;
  wire _14014_;
  wire _14015_;
  wire _14016_;
  wire _14017_;
  wire _14018_;
  wire _14019_;
  wire _14020_;
  wire _14021_;
  wire _14022_;
  wire _14023_;
  wire _14024_;
  wire _14025_;
  wire _14026_;
  wire _14027_;
  wire _14028_;
  wire _14029_;
  wire _14030_;
  wire _14031_;
  wire _14032_;
  wire _14033_;
  wire _14034_;
  wire _14035_;
  wire _14036_;
  wire _14037_;
  wire _14038_;
  wire _14039_;
  wire _14040_;
  wire _14041_;
  wire _14042_;
  wire _14043_;
  wire _14044_;
  wire _14045_;
  wire _14046_;
  wire _14047_;
  wire _14048_;
  wire _14049_;
  wire _14050_;
  wire _14051_;
  wire _14052_;
  wire _14053_;
  wire _14054_;
  wire _14055_;
  wire _14056_;
  wire _14057_;
  wire _14058_;
  wire _14059_;
  wire _14060_;
  wire _14061_;
  wire _14062_;
  wire _14063_;
  wire _14064_;
  wire _14065_;
  wire _14066_;
  wire _14067_;
  wire _14068_;
  wire _14069_;
  wire _14070_;
  wire _14071_;
  wire _14072_;
  wire _14073_;
  wire _14074_;
  wire _14075_;
  wire _14076_;
  wire _14077_;
  wire _14078_;
  wire _14079_;
  wire _14080_;
  wire _14081_;
  wire _14082_;
  wire _14083_;
  wire _14084_;
  wire _14085_;
  wire _14086_;
  wire _14087_;
  wire _14088_;
  wire _14089_;
  wire _14090_;
  wire _14091_;
  wire _14092_;
  wire _14093_;
  wire _14094_;
  wire _14095_;
  wire _14096_;
  wire _14097_;
  wire _14098_;
  wire _14099_;
  wire _14100_;
  wire _14101_;
  wire _14102_;
  wire _14103_;
  wire _14104_;
  wire _14105_;
  wire _14106_;
  wire _14107_;
  wire _14108_;
  wire _14109_;
  wire _14110_;
  wire _14111_;
  wire _14112_;
  wire _14113_;
  wire _14114_;
  wire _14115_;
  wire _14116_;
  wire _14117_;
  wire _14118_;
  wire _14119_;
  wire _14120_;
  wire _14121_;
  wire _14122_;
  wire _14123_;
  wire _14124_;
  wire _14125_;
  wire _14126_;
  wire _14127_;
  wire _14128_;
  wire _14129_;
  wire _14130_;
  wire _14131_;
  wire _14132_;
  wire _14133_;
  wire _14134_;
  wire _14135_;
  wire _14136_;
  wire _14137_;
  wire _14138_;
  wire _14139_;
  wire _14140_;
  wire _14141_;
  wire _14142_;
  wire _14143_;
  wire _14144_;
  wire _14145_;
  wire _14146_;
  wire _14147_;
  wire _14148_;
  wire _14149_;
  wire _14150_;
  wire _14151_;
  wire _14152_;
  wire _14153_;
  wire _14154_;
  wire _14155_;
  wire _14156_;
  wire _14157_;
  wire _14158_;
  wire _14159_;
  wire _14160_;
  wire _14161_;
  wire _14162_;
  wire _14163_;
  wire _14164_;
  wire _14165_;
  wire _14166_;
  wire _14167_;
  wire _14168_;
  wire _14169_;
  wire _14170_;
  wire _14171_;
  wire _14172_;
  wire _14173_;
  wire _14174_;
  wire _14175_;
  wire _14176_;
  wire _14177_;
  wire _14178_;
  wire _14179_;
  wire _14180_;
  wire _14181_;
  wire _14182_;
  wire _14183_;
  wire _14184_;
  wire _14185_;
  wire _14186_;
  wire _14187_;
  wire _14188_;
  wire _14189_;
  wire _14190_;
  wire _14191_;
  wire _14192_;
  wire _14193_;
  wire _14194_;
  wire _14195_;
  wire _14196_;
  wire _14197_;
  wire _14198_;
  wire _14199_;
  wire _14200_;
  wire _14201_;
  wire _14202_;
  wire _14203_;
  wire _14204_;
  wire _14205_;
  wire _14206_;
  wire _14207_;
  wire _14208_;
  wire _14209_;
  wire _14210_;
  wire _14211_;
  wire _14212_;
  wire _14213_;
  wire _14214_;
  wire _14215_;
  wire _14216_;
  wire _14217_;
  wire _14218_;
  wire _14219_;
  wire _14220_;
  wire _14221_;
  wire _14222_;
  wire _14223_;
  wire _14224_;
  wire _14225_;
  wire _14226_;
  wire _14227_;
  wire _14228_;
  wire _14229_;
  wire _14230_;
  wire _14231_;
  wire _14232_;
  wire _14233_;
  wire _14234_;
  wire _14235_;
  wire _14236_;
  wire _14237_;
  wire _14238_;
  wire _14239_;
  wire _14240_;
  wire _14241_;
  wire _14242_;
  wire _14243_;
  wire _14244_;
  wire _14245_;
  wire _14246_;
  wire _14247_;
  wire _14248_;
  wire _14249_;
  wire _14250_;
  wire _14251_;
  wire _14252_;
  wire _14253_;
  wire _14254_;
  wire _14255_;
  wire _14256_;
  wire _14257_;
  wire _14258_;
  wire _14259_;
  wire _14260_;
  wire _14261_;
  wire _14262_;
  wire _14263_;
  wire _14264_;
  wire _14265_;
  wire _14266_;
  wire _14267_;
  wire _14268_;
  wire _14269_;
  wire _14270_;
  wire _14271_;
  wire _14272_;
  wire _14273_;
  wire _14274_;
  wire _14275_;
  wire _14276_;
  wire _14277_;
  wire _14278_;
  wire _14279_;
  wire _14280_;
  wire _14281_;
  wire _14282_;
  wire _14283_;
  wire _14284_;
  wire _14285_;
  wire _14286_;
  wire _14287_;
  wire _14288_;
  wire _14289_;
  wire _14290_;
  wire _14291_;
  wire _14292_;
  wire _14293_;
  wire _14294_;
  wire _14295_;
  wire _14296_;
  wire _14297_;
  wire _14298_;
  wire _14299_;
  wire _14300_;
  wire _14301_;
  wire _14302_;
  wire _14303_;
  wire _14304_;
  wire _14305_;
  wire _14306_;
  wire _14307_;
  wire _14308_;
  wire _14309_;
  wire _14310_;
  wire _14311_;
  wire _14312_;
  wire _14313_;
  wire _14314_;
  wire _14315_;
  wire _14316_;
  wire _14317_;
  wire _14318_;
  wire _14319_;
  wire _14320_;
  wire _14321_;
  wire _14322_;
  wire _14323_;
  wire _14324_;
  wire _14325_;
  wire _14326_;
  wire _14327_;
  wire _14328_;
  wire _14329_;
  wire _14330_;
  wire _14331_;
  wire _14332_;
  wire _14333_;
  wire _14334_;
  wire _14335_;
  wire _14336_;
  wire _14337_;
  wire _14338_;
  wire _14339_;
  wire _14340_;
  wire _14341_;
  wire _14342_;
  wire _14343_;
  wire _14344_;
  wire _14345_;
  wire _14346_;
  wire _14347_;
  wire _14348_;
  wire _14349_;
  wire _14350_;
  wire _14351_;
  wire _14352_;
  wire _14353_;
  wire _14354_;
  wire _14355_;
  wire _14356_;
  wire _14357_;
  wire _14358_;
  wire _14359_;
  wire _14360_;
  wire _14361_;
  wire _14362_;
  wire _14363_;
  wire _14364_;
  wire _14365_;
  wire _14366_;
  wire _14367_;
  wire _14368_;
  wire _14369_;
  wire _14370_;
  wire _14371_;
  wire _14372_;
  wire _14373_;
  wire _14374_;
  wire _14375_;
  wire _14376_;
  wire _14377_;
  wire _14378_;
  wire _14379_;
  wire _14380_;
  wire _14381_;
  wire _14382_;
  wire _14383_;
  wire _14384_;
  wire _14385_;
  wire _14386_;
  wire _14387_;
  wire _14388_;
  wire _14389_;
  wire _14390_;
  wire _14391_;
  wire _14392_;
  wire _14393_;
  wire _14394_;
  wire _14395_;
  wire _14396_;
  wire _14397_;
  wire _14398_;
  wire _14399_;
  wire _14400_;
  wire _14401_;
  wire _14402_;
  wire _14403_;
  wire _14404_;
  wire _14405_;
  wire _14406_;
  wire _14407_;
  wire _14408_;
  wire _14409_;
  wire _14410_;
  wire _14411_;
  wire _14412_;
  wire _14413_;
  wire _14414_;
  wire _14415_;
  wire _14416_;
  wire _14417_;
  wire _14418_;
  wire _14419_;
  wire _14420_;
  wire _14421_;
  wire _14422_;
  wire _14423_;
  wire _14424_;
  wire _14425_;
  wire _14426_;
  wire _14427_;
  wire _14428_;
  wire _14429_;
  wire _14430_;
  wire _14431_;
  wire _14432_;
  wire _14433_;
  wire _14434_;
  wire _14435_;
  wire _14436_;
  wire _14437_;
  wire _14438_;
  wire _14439_;
  wire _14440_;
  wire _14441_;
  wire _14442_;
  wire _14443_;
  wire _14444_;
  wire _14445_;
  wire _14446_;
  wire _14447_;
  wire _14448_;
  wire _14449_;
  wire _14450_;
  wire _14451_;
  wire _14452_;
  wire _14453_;
  wire _14454_;
  wire _14455_;
  wire _14456_;
  wire _14457_;
  wire _14458_;
  wire _14459_;
  wire _14460_;
  wire _14461_;
  wire _14462_;
  wire _14463_;
  wire _14464_;
  wire _14465_;
  wire _14466_;
  wire _14467_;
  wire _14468_;
  wire _14469_;
  wire _14470_;
  wire _14471_;
  wire _14472_;
  wire _14473_;
  wire _14474_;
  wire _14475_;
  wire _14476_;
  wire _14477_;
  wire _14478_;
  wire _14479_;
  wire _14480_;
  wire _14481_;
  wire _14482_;
  wire _14483_;
  wire _14484_;
  wire _14485_;
  wire _14486_;
  wire _14487_;
  wire _14488_;
  wire _14489_;
  wire _14490_;
  wire _14491_;
  wire _14492_;
  wire _14493_;
  wire _14494_;
  wire _14495_;
  wire _14496_;
  wire _14497_;
  wire _14498_;
  wire _14499_;
  wire _14500_;
  wire _14501_;
  wire _14502_;
  wire _14503_;
  wire _14504_;
  wire _14505_;
  wire _14506_;
  wire _14507_;
  wire _14508_;
  wire _14509_;
  wire _14510_;
  wire _14511_;
  wire _14512_;
  wire _14513_;
  wire _14514_;
  wire _14515_;
  wire _14516_;
  wire _14517_;
  wire _14518_;
  wire _14519_;
  wire _14520_;
  wire _14521_;
  wire _14522_;
  wire _14523_;
  wire _14524_;
  wire _14525_;
  wire _14526_;
  wire _14527_;
  wire _14528_;
  wire _14529_;
  wire _14530_;
  wire _14531_;
  wire _14532_;
  wire _14533_;
  wire _14534_;
  wire _14535_;
  wire _14536_;
  wire _14537_;
  wire _14538_;
  wire _14539_;
  wire _14540_;
  wire _14541_;
  wire _14542_;
  wire _14543_;
  wire _14544_;
  wire _14545_;
  wire _14546_;
  wire _14547_;
  wire _14548_;
  wire _14549_;
  wire _14550_;
  wire _14551_;
  wire _14552_;
  wire _14553_;
  wire _14554_;
  wire _14555_;
  wire _14556_;
  wire _14557_;
  wire _14558_;
  wire _14559_;
  wire _14560_;
  wire _14561_;
  wire _14562_;
  wire _14563_;
  wire _14564_;
  wire _14565_;
  wire _14566_;
  wire _14567_;
  wire _14568_;
  wire _14569_;
  wire _14570_;
  wire _14571_;
  wire _14572_;
  wire _14573_;
  wire _14574_;
  wire _14575_;
  wire _14576_;
  wire _14577_;
  wire _14578_;
  wire _14579_;
  wire _14580_;
  wire _14581_;
  wire _14582_;
  wire _14583_;
  wire _14584_;
  wire _14585_;
  wire _14586_;
  wire _14587_;
  wire _14588_;
  wire _14589_;
  wire _14590_;
  wire _14591_;
  wire _14592_;
  wire _14593_;
  wire _14594_;
  wire _14595_;
  wire _14596_;
  wire _14597_;
  wire _14598_;
  wire _14599_;
  wire _14600_;
  wire _14601_;
  wire _14602_;
  wire _14603_;
  wire _14604_;
  wire _14605_;
  wire _14606_;
  wire _14607_;
  wire _14608_;
  wire _14609_;
  wire _14610_;
  wire _14611_;
  wire _14612_;
  wire _14613_;
  wire _14614_;
  wire _14615_;
  wire _14616_;
  wire _14617_;
  wire _14618_;
  wire _14619_;
  wire _14620_;
  wire _14621_;
  wire _14622_;
  wire _14623_;
  wire _14624_;
  wire _14625_;
  wire _14626_;
  wire _14627_;
  wire _14628_;
  wire _14629_;
  wire _14630_;
  wire _14631_;
  wire _14632_;
  wire _14633_;
  wire _14634_;
  wire _14635_;
  wire _14636_;
  wire _14637_;
  wire _14638_;
  wire _14639_;
  wire _14640_;
  wire _14641_;
  wire _14642_;
  wire _14643_;
  wire _14644_;
  wire _14645_;
  wire _14646_;
  wire _14647_;
  wire _14648_;
  wire _14649_;
  wire _14650_;
  wire _14651_;
  wire _14652_;
  wire _14653_;
  wire _14654_;
  wire _14655_;
  wire _14656_;
  wire _14657_;
  wire _14658_;
  wire _14659_;
  wire _14660_;
  wire _14661_;
  wire _14662_;
  wire _14663_;
  wire _14664_;
  wire _14665_;
  wire _14666_;
  wire _14667_;
  wire _14668_;
  wire _14669_;
  wire _14670_;
  wire _14671_;
  wire _14672_;
  wire _14673_;
  wire _14674_;
  wire _14675_;
  wire _14676_;
  wire _14677_;
  wire _14678_;
  wire _14679_;
  wire _14680_;
  wire _14681_;
  wire _14682_;
  wire _14683_;
  wire _14684_;
  wire _14685_;
  wire _14686_;
  wire _14687_;
  wire _14688_;
  wire _14689_;
  wire _14690_;
  wire _14691_;
  wire _14692_;
  wire _14693_;
  wire _14694_;
  wire _14695_;
  wire _14696_;
  wire _14697_;
  wire _14698_;
  wire _14699_;
  wire _14700_;
  wire _14701_;
  wire _14702_;
  wire _14703_;
  wire _14704_;
  wire _14705_;
  wire _14706_;
  wire _14707_;
  wire _14708_;
  wire _14709_;
  wire _14710_;
  wire _14711_;
  wire _14712_;
  wire _14713_;
  wire _14714_;
  wire _14715_;
  wire _14716_;
  wire _14717_;
  wire _14718_;
  wire _14719_;
  wire _14720_;
  wire _14721_;
  wire _14722_;
  wire _14723_;
  wire _14724_;
  wire _14725_;
  wire _14726_;
  wire _14727_;
  wire _14728_;
  wire _14729_;
  wire _14730_;
  wire _14731_;
  wire _14732_;
  wire _14733_;
  wire _14734_;
  wire _14735_;
  wire _14736_;
  wire _14737_;
  wire _14738_;
  wire _14739_;
  wire _14740_;
  wire _14741_;
  wire _14742_;
  wire _14743_;
  wire _14744_;
  wire _14745_;
  wire _14746_;
  wire _14747_;
  wire _14748_;
  wire _14749_;
  wire _14750_;
  wire _14751_;
  wire _14752_;
  wire _14753_;
  wire _14754_;
  wire _14755_;
  wire _14756_;
  wire _14757_;
  wire _14758_;
  wire _14759_;
  wire _14760_;
  wire _14761_;
  wire _14762_;
  wire _14763_;
  wire _14764_;
  wire _14765_;
  wire _14766_;
  wire _14767_;
  wire _14768_;
  wire _14769_;
  wire _14770_;
  wire _14771_;
  wire _14772_;
  wire _14773_;
  wire _14774_;
  wire _14775_;
  wire _14776_;
  wire _14777_;
  wire _14778_;
  wire _14779_;
  wire _14780_;
  wire _14781_;
  wire _14782_;
  wire _14783_;
  wire _14784_;
  wire _14785_;
  wire _14786_;
  wire _14787_;
  wire _14788_;
  wire _14789_;
  wire _14790_;
  wire _14791_;
  wire _14792_;
  wire _14793_;
  wire _14794_;
  wire _14795_;
  wire _14796_;
  wire _14797_;
  wire _14798_;
  wire _14799_;
  wire _14800_;
  wire _14801_;
  wire _14802_;
  wire _14803_;
  wire _14804_;
  wire _14805_;
  wire _14806_;
  wire _14807_;
  wire _14808_;
  wire _14809_;
  wire _14810_;
  wire _14811_;
  wire _14812_;
  wire _14813_;
  wire _14814_;
  wire _14815_;
  wire _14816_;
  wire _14817_;
  wire _14818_;
  wire _14819_;
  wire _14820_;
  wire _14821_;
  wire _14822_;
  wire _14823_;
  wire _14824_;
  wire _14825_;
  wire _14826_;
  wire _14827_;
  wire _14828_;
  wire _14829_;
  wire _14830_;
  wire _14831_;
  wire _14832_;
  wire _14833_;
  wire _14834_;
  wire _14835_;
  wire _14836_;
  wire _14837_;
  wire _14838_;
  wire _14839_;
  wire _14840_;
  wire _14841_;
  wire _14842_;
  wire _14843_;
  wire _14844_;
  wire _14845_;
  wire _14846_;
  wire _14847_;
  wire _14848_;
  wire _14849_;
  wire _14850_;
  wire _14851_;
  wire _14852_;
  wire _14853_;
  wire _14854_;
  wire _14855_;
  wire _14856_;
  wire _14857_;
  wire _14858_;
  wire _14859_;
  wire _14860_;
  wire _14861_;
  wire _14862_;
  wire _14863_;
  wire _14864_;
  wire _14865_;
  wire _14866_;
  wire _14867_;
  wire _14868_;
  wire _14869_;
  wire _14870_;
  wire _14871_;
  wire _14872_;
  wire _14873_;
  wire _14874_;
  wire _14875_;
  wire _14876_;
  wire _14877_;
  wire _14878_;
  wire _14879_;
  wire _14880_;
  wire _14881_;
  wire _14882_;
  wire _14883_;
  wire _14884_;
  wire _14885_;
  wire _14886_;
  wire _14887_;
  wire _14888_;
  wire _14889_;
  wire _14890_;
  wire _14891_;
  wire _14892_;
  wire _14893_;
  wire _14894_;
  wire _14895_;
  wire _14896_;
  wire _14897_;
  wire _14898_;
  wire _14899_;
  wire _14900_;
  wire _14901_;
  wire _14902_;
  wire _14903_;
  wire _14904_;
  wire _14905_;
  wire _14906_;
  wire _14907_;
  wire _14908_;
  wire _14909_;
  wire _14910_;
  wire _14911_;
  wire _14912_;
  wire _14913_;
  wire _14914_;
  wire _14915_;
  wire _14916_;
  wire _14917_;
  wire _14918_;
  wire _14919_;
  wire _14920_;
  wire _14921_;
  wire _14922_;
  wire _14923_;
  wire _14924_;
  wire _14925_;
  wire _14926_;
  wire _14927_;
  wire _14928_;
  wire _14929_;
  wire _14930_;
  wire _14931_;
  wire _14932_;
  wire _14933_;
  wire _14934_;
  wire _14935_;
  wire _14936_;
  wire _14937_;
  wire _14938_;
  wire _14939_;
  wire _14940_;
  wire _14941_;
  wire _14942_;
  wire _14943_;
  wire _14944_;
  wire _14945_;
  wire _14946_;
  wire _14947_;
  wire _14948_;
  wire _14949_;
  wire _14950_;
  wire _14951_;
  wire _14952_;
  wire _14953_;
  wire _14954_;
  wire _14955_;
  wire _14956_;
  wire _14957_;
  wire _14958_;
  wire _14959_;
  wire _14960_;
  wire _14961_;
  wire _14962_;
  wire _14963_;
  wire _14964_;
  wire _14965_;
  wire _14966_;
  wire _14967_;
  wire _14968_;
  wire _14969_;
  wire _14970_;
  wire _14971_;
  wire _14972_;
  wire _14973_;
  wire _14974_;
  wire _14975_;
  wire _14976_;
  wire _14977_;
  wire _14978_;
  wire _14979_;
  wire _14980_;
  wire _14981_;
  wire _14982_;
  wire _14983_;
  wire _14984_;
  wire _14985_;
  wire _14986_;
  wire _14987_;
  wire _14988_;
  wire _14989_;
  wire _14990_;
  wire _14991_;
  wire _14992_;
  wire _14993_;
  wire _14994_;
  wire _14995_;
  wire _14996_;
  wire _14997_;
  wire _14998_;
  wire _14999_;
  wire _15000_;
  wire _15001_;
  wire _15002_;
  wire _15003_;
  wire _15004_;
  wire _15005_;
  wire _15006_;
  wire _15007_;
  wire _15008_;
  wire _15009_;
  wire _15010_;
  wire _15011_;
  wire _15012_;
  wire _15013_;
  wire _15014_;
  wire _15015_;
  wire _15016_;
  wire _15017_;
  wire _15018_;
  wire _15019_;
  wire _15020_;
  wire _15021_;
  wire _15022_;
  wire _15023_;
  wire _15024_;
  wire _15025_;
  wire _15026_;
  wire _15027_;
  wire _15028_;
  wire _15029_;
  wire _15030_;
  wire _15031_;
  wire _15032_;
  wire _15033_;
  wire _15034_;
  wire _15035_;
  wire _15036_;
  wire _15037_;
  wire _15038_;
  wire _15039_;
  wire _15040_;
  wire _15041_;
  wire _15042_;
  wire _15043_;
  wire _15044_;
  wire _15045_;
  wire _15046_;
  wire _15047_;
  wire _15048_;
  wire _15049_;
  wire _15050_;
  wire _15051_;
  wire _15052_;
  wire _15053_;
  wire _15054_;
  wire _15055_;
  wire _15056_;
  wire _15057_;
  wire _15058_;
  wire _15059_;
  wire _15060_;
  wire _15061_;
  wire _15062_;
  wire _15063_;
  wire _15064_;
  wire _15065_;
  wire _15066_;
  wire _15067_;
  wire _15068_;
  wire _15069_;
  wire _15070_;
  wire _15071_;
  wire _15072_;
  wire _15073_;
  wire _15074_;
  wire _15075_;
  wire _15076_;
  wire _15077_;
  wire _15078_;
  wire _15079_;
  wire _15080_;
  wire _15081_;
  wire _15082_;
  wire _15083_;
  wire _15084_;
  wire _15085_;
  wire _15086_;
  wire _15087_;
  wire _15088_;
  wire _15089_;
  wire _15090_;
  wire _15091_;
  wire _15092_;
  wire _15093_;
  wire _15094_;
  wire _15095_;
  wire _15096_;
  wire _15097_;
  wire _15098_;
  wire _15099_;
  wire _15100_;
  wire _15101_;
  wire _15102_;
  wire _15103_;
  wire _15104_;
  wire _15105_;
  wire _15106_;
  wire _15107_;
  wire _15108_;
  wire _15109_;
  wire _15110_;
  wire _15111_;
  wire _15112_;
  wire _15113_;
  wire _15114_;
  wire _15115_;
  wire _15116_;
  wire _15117_;
  wire _15118_;
  wire _15119_;
  wire _15120_;
  wire _15121_;
  wire _15122_;
  wire _15123_;
  wire _15124_;
  wire _15125_;
  wire _15126_;
  wire _15127_;
  wire _15128_;
  wire _15129_;
  wire _15130_;
  wire _15131_;
  wire _15132_;
  wire _15133_;
  wire _15134_;
  wire _15135_;
  wire _15136_;
  wire _15137_;
  wire _15138_;
  wire _15139_;
  wire _15140_;
  wire _15141_;
  wire _15142_;
  wire _15143_;
  wire _15144_;
  wire _15145_;
  wire _15146_;
  wire _15147_;
  wire _15148_;
  wire _15149_;
  wire _15150_;
  wire _15151_;
  wire _15152_;
  wire _15153_;
  wire _15154_;
  wire _15155_;
  wire _15156_;
  wire _15157_;
  wire _15158_;
  wire _15159_;
  wire _15160_;
  wire _15161_;
  wire _15162_;
  wire _15163_;
  wire _15164_;
  wire _15165_;
  wire _15166_;
  wire _15167_;
  wire _15168_;
  wire _15169_;
  wire _15170_;
  wire _15171_;
  wire _15172_;
  wire _15173_;
  wire _15174_;
  wire _15175_;
  wire _15176_;
  wire _15177_;
  wire _15178_;
  wire _15179_;
  wire _15180_;
  wire _15181_;
  wire _15182_;
  wire _15183_;
  wire _15184_;
  wire _15185_;
  wire _15186_;
  wire _15187_;
  wire _15188_;
  wire _15189_;
  wire _15190_;
  wire _15191_;
  wire _15192_;
  wire _15193_;
  wire _15194_;
  wire _15195_;
  wire _15196_;
  wire _15197_;
  wire _15198_;
  wire _15199_;
  wire _15200_;
  wire _15201_;
  wire _15202_;
  wire _15203_;
  wire _15204_;
  wire _15205_;
  wire _15206_;
  wire _15207_;
  wire _15208_;
  wire _15209_;
  wire _15210_;
  wire _15211_;
  wire _15212_;
  wire _15213_;
  wire _15214_;
  wire _15215_;
  wire _15216_;
  wire _15217_;
  wire _15218_;
  wire _15219_;
  wire _15220_;
  wire _15221_;
  wire _15222_;
  wire _15223_;
  wire _15224_;
  wire _15225_;
  wire _15226_;
  wire _15227_;
  wire _15228_;
  wire _15229_;
  wire _15230_;
  wire _15231_;
  wire _15232_;
  wire _15233_;
  wire _15234_;
  wire _15235_;
  wire _15236_;
  wire _15237_;
  wire _15238_;
  wire _15239_;
  wire _15240_;
  wire _15241_;
  wire _15242_;
  wire _15243_;
  wire _15244_;
  wire _15245_;
  wire _15246_;
  wire _15247_;
  wire _15248_;
  wire _15249_;
  wire _15250_;
  wire _15251_;
  wire _15252_;
  wire _15253_;
  wire _15254_;
  wire _15255_;
  wire _15256_;
  wire _15257_;
  wire _15258_;
  wire _15259_;
  wire _15260_;
  wire _15261_;
  wire _15262_;
  wire _15263_;
  wire _15264_;
  wire _15265_;
  wire _15266_;
  wire _15267_;
  wire _15268_;
  wire _15269_;
  wire _15270_;
  wire _15271_;
  wire _15272_;
  wire _15273_;
  wire _15274_;
  wire _15275_;
  wire _15276_;
  wire _15277_;
  wire _15278_;
  wire _15279_;
  wire _15280_;
  wire _15281_;
  wire _15282_;
  wire _15283_;
  wire _15284_;
  wire _15285_;
  wire _15286_;
  wire _15287_;
  wire _15288_;
  wire _15289_;
  wire _15290_;
  wire _15291_;
  wire _15292_;
  wire _15293_;
  wire _15294_;
  wire _15295_;
  wire _15296_;
  wire _15297_;
  wire _15298_;
  wire _15299_;
  wire _15300_;
  wire _15301_;
  wire _15302_;
  wire _15303_;
  wire _15304_;
  wire _15305_;
  wire _15306_;
  wire _15307_;
  wire _15308_;
  wire _15309_;
  wire _15310_;
  wire _15311_;
  wire _15312_;
  wire _15313_;
  wire _15314_;
  wire _15315_;
  wire _15316_;
  wire _15317_;
  wire _15318_;
  wire _15319_;
  wire _15320_;
  wire _15321_;
  wire _15322_;
  wire _15323_;
  wire _15324_;
  wire _15325_;
  wire _15326_;
  wire _15327_;
  wire _15328_;
  wire _15329_;
  wire _15330_;
  wire _15331_;
  wire _15332_;
  wire _15333_;
  wire _15334_;
  wire _15335_;
  wire _15336_;
  wire _15337_;
  wire _15338_;
  wire _15339_;
  wire _15340_;
  wire _15341_;
  wire _15342_;
  wire _15343_;
  wire _15344_;
  wire _15345_;
  wire _15346_;
  wire _15347_;
  wire _15348_;
  wire _15349_;
  wire _15350_;
  wire _15351_;
  wire _15352_;
  wire _15353_;
  wire _15354_;
  wire _15355_;
  wire _15356_;
  wire _15357_;
  wire _15358_;
  wire _15359_;
  wire _15360_;
  wire _15361_;
  wire _15362_;
  wire _15363_;
  wire _15364_;
  wire _15365_;
  wire _15366_;
  wire _15367_;
  wire _15368_;
  wire _15369_;
  wire _15370_;
  wire _15371_;
  wire _15372_;
  wire _15373_;
  wire _15374_;
  wire _15375_;
  wire _15376_;
  wire _15377_;
  wire _15378_;
  wire _15379_;
  wire _15380_;
  wire _15381_;
  wire _15382_;
  wire _15383_;
  wire _15384_;
  wire _15385_;
  wire _15386_;
  wire _15387_;
  wire _15388_;
  wire _15389_;
  wire _15390_;
  wire _15391_;
  wire _15392_;
  wire _15393_;
  wire _15394_;
  wire _15395_;
  wire _15396_;
  wire _15397_;
  wire _15398_;
  wire _15399_;
  wire _15400_;
  wire _15401_;
  wire _15402_;
  wire _15403_;
  wire _15404_;
  wire _15405_;
  wire _15406_;
  wire _15407_;
  wire _15408_;
  wire _15409_;
  wire _15410_;
  wire _15411_;
  wire _15412_;
  wire _15413_;
  wire _15414_;
  wire _15415_;
  wire _15416_;
  wire _15417_;
  wire _15418_;
  wire _15419_;
  wire _15420_;
  wire _15421_;
  wire _15422_;
  wire _15423_;
  wire _15424_;
  wire _15425_;
  wire _15426_;
  wire _15427_;
  wire _15428_;
  wire _15429_;
  wire _15430_;
  wire _15431_;
  wire _15432_;
  wire _15433_;
  wire _15434_;
  wire _15435_;
  wire _15436_;
  wire _15437_;
  wire _15438_;
  wire _15439_;
  wire _15440_;
  wire _15441_;
  wire _15442_;
  wire _15443_;
  wire _15444_;
  wire _15445_;
  wire _15446_;
  wire _15447_;
  wire _15448_;
  wire _15449_;
  wire _15450_;
  wire _15451_;
  wire _15452_;
  wire _15453_;
  wire _15454_;
  wire _15455_;
  wire _15456_;
  wire _15457_;
  wire _15458_;
  wire _15459_;
  wire _15460_;
  wire _15461_;
  wire _15462_;
  wire _15463_;
  wire _15464_;
  wire _15465_;
  wire _15466_;
  wire _15467_;
  wire _15468_;
  wire _15469_;
  wire _15470_;
  wire _15471_;
  wire _15472_;
  wire _15473_;
  wire _15474_;
  wire _15475_;
  wire _15476_;
  wire _15477_;
  wire _15478_;
  wire _15479_;
  wire _15480_;
  wire _15481_;
  wire _15482_;
  wire _15483_;
  wire _15484_;
  wire _15485_;
  wire _15486_;
  wire _15487_;
  wire _15488_;
  wire _15489_;
  wire _15490_;
  wire _15491_;
  wire _15492_;
  wire _15493_;
  wire _15494_;
  wire _15495_;
  wire _15496_;
  wire _15497_;
  wire _15498_;
  wire _15499_;
  wire _15500_;
  wire _15501_;
  wire _15502_;
  wire _15503_;
  wire _15504_;
  wire _15505_;
  wire _15506_;
  wire _15507_;
  wire _15508_;
  wire _15509_;
  wire _15510_;
  wire _15511_;
  wire _15512_;
  wire _15513_;
  wire _15514_;
  wire _15515_;
  wire _15516_;
  wire _15517_;
  wire _15518_;
  wire _15519_;
  wire _15520_;
  wire _15521_;
  wire _15522_;
  wire _15523_;
  wire _15524_;
  wire _15525_;
  wire _15526_;
  wire _15527_;
  wire _15528_;
  wire _15529_;
  wire _15530_;
  wire _15531_;
  wire _15532_;
  wire _15533_;
  wire _15534_;
  wire _15535_;
  wire _15536_;
  wire _15537_;
  wire _15538_;
  wire _15539_;
  wire _15540_;
  wire _15541_;
  wire _15542_;
  wire _15543_;
  wire _15544_;
  wire _15545_;
  wire _15546_;
  wire _15547_;
  wire _15548_;
  wire _15549_;
  wire _15550_;
  wire _15551_;
  wire _15552_;
  wire _15553_;
  wire _15554_;
  wire _15555_;
  wire _15556_;
  wire _15557_;
  wire _15558_;
  wire _15559_;
  wire _15560_;
  wire _15561_;
  wire _15562_;
  wire _15563_;
  wire _15564_;
  wire _15565_;
  wire _15566_;
  wire _15567_;
  wire _15568_;
  wire _15569_;
  wire _15570_;
  wire _15571_;
  wire _15572_;
  wire _15573_;
  wire _15574_;
  wire _15575_;
  wire _15576_;
  wire _15577_;
  wire _15578_;
  wire _15579_;
  wire _15580_;
  wire _15581_;
  wire _15582_;
  wire _15583_;
  wire _15584_;
  wire _15585_;
  wire _15586_;
  wire _15587_;
  wire _15588_;
  wire _15589_;
  wire _15590_;
  wire _15591_;
  wire _15592_;
  wire _15593_;
  wire _15594_;
  wire _15595_;
  wire _15596_;
  wire _15597_;
  wire _15598_;
  wire _15599_;
  wire _15600_;
  wire _15601_;
  wire _15602_;
  wire _15603_;
  wire _15604_;
  wire _15605_;
  wire _15606_;
  wire _15607_;
  wire _15608_;
  wire _15609_;
  wire _15610_;
  wire _15611_;
  wire _15612_;
  wire _15613_;
  wire _15614_;
  wire _15615_;
  wire _15616_;
  wire _15617_;
  wire _15618_;
  wire _15619_;
  wire _15620_;
  wire _15621_;
  wire _15622_;
  wire _15623_;
  wire _15624_;
  wire _15625_;
  wire _15626_;
  wire _15627_;
  wire _15628_;
  wire _15629_;
  wire _15630_;
  wire _15631_;
  wire _15632_;
  wire _15633_;
  wire _15634_;
  wire _15635_;
  wire _15636_;
  wire _15637_;
  wire _15638_;
  wire _15639_;
  wire _15640_;
  wire _15641_;
  wire _15642_;
  wire _15643_;
  wire _15644_;
  wire _15645_;
  wire _15646_;
  wire _15647_;
  wire _15648_;
  wire _15649_;
  wire _15650_;
  wire _15651_;
  wire _15652_;
  wire _15653_;
  wire _15654_;
  wire _15655_;
  wire _15656_;
  wire _15657_;
  wire _15658_;
  wire _15659_;
  wire _15660_;
  wire _15661_;
  wire _15662_;
  wire _15663_;
  wire _15664_;
  wire _15665_;
  wire _15666_;
  wire _15667_;
  wire _15668_;
  wire _15669_;
  wire _15670_;
  wire _15671_;
  wire _15672_;
  wire _15673_;
  wire _15674_;
  wire _15675_;
  wire _15676_;
  wire _15677_;
  wire _15678_;
  wire _15679_;
  wire _15680_;
  wire _15681_;
  wire _15682_;
  wire _15683_;
  wire _15684_;
  wire _15685_;
  wire _15686_;
  wire _15687_;
  wire _15688_;
  wire _15689_;
  wire _15690_;
  wire _15691_;
  wire _15692_;
  wire _15693_;
  wire _15694_;
  wire _15695_;
  wire _15696_;
  wire _15697_;
  wire _15698_;
  wire _15699_;
  wire _15700_;
  wire _15701_;
  wire _15702_;
  wire _15703_;
  wire _15704_;
  wire _15705_;
  wire _15706_;
  wire _15707_;
  wire _15708_;
  wire _15709_;
  wire _15710_;
  wire _15711_;
  wire _15712_;
  wire _15713_;
  wire _15714_;
  wire _15715_;
  wire _15716_;
  wire _15717_;
  wire _15718_;
  wire _15719_;
  wire _15720_;
  wire _15721_;
  wire _15722_;
  wire _15723_;
  wire _15724_;
  wire _15725_;
  wire _15726_;
  wire _15727_;
  wire _15728_;
  wire _15729_;
  wire _15730_;
  wire _15731_;
  wire _15732_;
  wire _15733_;
  wire _15734_;
  wire _15735_;
  wire _15736_;
  wire _15737_;
  wire _15738_;
  wire _15739_;
  wire _15740_;
  wire _15741_;
  wire _15742_;
  wire _15743_;
  wire _15744_;
  wire _15745_;
  wire _15746_;
  wire _15747_;
  wire _15748_;
  wire _15749_;
  wire _15750_;
  wire _15751_;
  wire _15752_;
  wire _15753_;
  wire _15754_;
  wire _15755_;
  wire _15756_;
  wire _15757_;
  wire _15758_;
  wire _15759_;
  wire _15760_;
  wire _15761_;
  wire _15762_;
  wire _15763_;
  wire _15764_;
  wire _15765_;
  wire _15766_;
  wire _15767_;
  wire _15768_;
  wire _15769_;
  wire _15770_;
  wire _15771_;
  wire _15772_;
  wire _15773_;
  wire _15774_;
  wire _15775_;
  wire _15776_;
  wire _15777_;
  wire _15778_;
  wire _15779_;
  wire _15780_;
  wire _15781_;
  wire _15782_;
  wire _15783_;
  wire _15784_;
  wire _15785_;
  wire _15786_;
  wire _15787_;
  wire _15788_;
  wire _15789_;
  wire _15790_;
  wire _15791_;
  wire _15792_;
  wire _15793_;
  wire _15794_;
  wire _15795_;
  wire _15796_;
  wire _15797_;
  wire _15798_;
  wire _15799_;
  wire _15800_;
  wire _15801_;
  wire _15802_;
  wire _15803_;
  wire _15804_;
  wire _15805_;
  wire _15806_;
  wire _15807_;
  wire _15808_;
  wire _15809_;
  wire _15810_;
  wire _15811_;
  wire _15812_;
  wire _15813_;
  wire _15814_;
  wire _15815_;
  wire _15816_;
  wire _15817_;
  wire _15818_;
  wire _15819_;
  wire _15820_;
  wire _15821_;
  wire _15822_;
  wire _15823_;
  wire _15824_;
  wire _15825_;
  wire _15826_;
  wire _15827_;
  wire _15828_;
  wire _15829_;
  wire _15830_;
  wire _15831_;
  wire _15832_;
  wire _15833_;
  wire _15834_;
  wire _15835_;
  wire _15836_;
  wire _15837_;
  wire _15838_;
  wire _15839_;
  wire _15840_;
  wire _15841_;
  wire _15842_;
  wire _15843_;
  wire _15844_;
  wire _15845_;
  wire _15846_;
  wire _15847_;
  wire _15848_;
  wire _15849_;
  wire _15850_;
  wire _15851_;
  wire _15852_;
  wire _15853_;
  wire _15854_;
  wire _15855_;
  wire _15856_;
  wire _15857_;
  wire _15858_;
  wire _15859_;
  wire _15860_;
  wire _15861_;
  wire _15862_;
  wire _15863_;
  wire _15864_;
  wire _15865_;
  wire _15866_;
  wire _15867_;
  wire _15868_;
  wire _15869_;
  wire _15870_;
  wire _15871_;
  wire _15872_;
  wire _15873_;
  wire _15874_;
  wire _15875_;
  wire _15876_;
  wire _15877_;
  wire _15878_;
  wire _15879_;
  wire _15880_;
  wire _15881_;
  wire _15882_;
  wire _15883_;
  wire _15884_;
  wire _15885_;
  wire _15886_;
  wire _15887_;
  wire _15888_;
  wire _15889_;
  wire _15890_;
  wire _15891_;
  wire _15892_;
  wire _15893_;
  wire _15894_;
  wire _15895_;
  wire _15896_;
  wire _15897_;
  wire _15898_;
  wire _15899_;
  wire _15900_;
  wire _15901_;
  wire _15902_;
  wire _15903_;
  wire _15904_;
  wire _15905_;
  wire _15906_;
  wire _15907_;
  wire _15908_;
  wire _15909_;
  wire _15910_;
  wire _15911_;
  wire _15912_;
  wire _15913_;
  wire _15914_;
  wire _15915_;
  wire _15916_;
  wire _15917_;
  wire _15918_;
  wire _15919_;
  wire _15920_;
  wire _15921_;
  wire _15922_;
  wire _15923_;
  wire _15924_;
  wire _15925_;
  wire _15926_;
  wire _15927_;
  wire _15928_;
  wire _15929_;
  wire _15930_;
  wire _15931_;
  wire _15932_;
  wire _15933_;
  wire _15934_;
  wire _15935_;
  wire _15936_;
  wire _15937_;
  wire _15938_;
  wire _15939_;
  wire _15940_;
  wire _15941_;
  wire _15942_;
  wire _15943_;
  wire _15944_;
  wire _15945_;
  wire _15946_;
  wire _15947_;
  wire _15948_;
  wire _15949_;
  wire _15950_;
  wire _15951_;
  wire _15952_;
  wire _15953_;
  wire _15954_;
  wire _15955_;
  wire _15956_;
  wire _15957_;
  wire _15958_;
  wire _15959_;
  wire _15960_;
  wire _15961_;
  wire _15962_;
  wire _15963_;
  wire _15964_;
  wire _15965_;
  wire _15966_;
  wire _15967_;
  wire _15968_;
  wire _15969_;
  wire _15970_;
  wire _15971_;
  wire _15972_;
  wire _15973_;
  wire _15974_;
  wire _15975_;
  wire _15976_;
  wire _15977_;
  wire _15978_;
  wire _15979_;
  wire _15980_;
  wire _15981_;
  wire _15982_;
  wire _15983_;
  wire _15984_;
  wire _15985_;
  wire _15986_;
  wire _15987_;
  wire _15988_;
  wire _15989_;
  wire _15990_;
  wire _15991_;
  wire _15992_;
  wire _15993_;
  wire _15994_;
  wire _15995_;
  wire _15996_;
  wire _15997_;
  wire _15998_;
  wire _15999_;
  wire _16000_;
  wire _16001_;
  wire _16002_;
  wire _16003_;
  wire _16004_;
  wire _16005_;
  wire _16006_;
  wire _16007_;
  wire _16008_;
  wire _16009_;
  wire _16010_;
  wire _16011_;
  wire _16012_;
  wire _16013_;
  wire _16014_;
  wire _16015_;
  wire _16016_;
  wire _16017_;
  wire _16018_;
  wire _16019_;
  wire _16020_;
  wire _16021_;
  wire _16022_;
  wire _16023_;
  wire _16024_;
  wire _16025_;
  wire _16026_;
  wire _16027_;
  wire _16028_;
  wire _16029_;
  wire _16030_;
  wire _16031_;
  wire _16032_;
  wire _16033_;
  wire _16034_;
  wire _16035_;
  wire _16036_;
  wire _16037_;
  wire _16038_;
  wire _16039_;
  wire _16040_;
  wire _16041_;
  wire _16042_;
  wire _16043_;
  wire _16044_;
  wire _16045_;
  wire _16046_;
  wire _16047_;
  wire _16048_;
  wire _16049_;
  wire _16050_;
  wire _16051_;
  wire _16052_;
  wire _16053_;
  wire _16054_;
  wire _16055_;
  wire _16056_;
  wire _16057_;
  wire _16058_;
  wire _16059_;
  wire _16060_;
  wire _16061_;
  wire _16062_;
  wire _16063_;
  wire _16064_;
  wire _16065_;
  wire _16066_;
  wire _16067_;
  wire _16068_;
  wire _16069_;
  wire _16070_;
  wire _16071_;
  wire _16072_;
  wire _16073_;
  wire _16074_;
  wire _16075_;
  wire _16076_;
  wire _16077_;
  wire _16078_;
  wire _16079_;
  wire _16080_;
  wire _16081_;
  wire _16082_;
  wire _16083_;
  wire _16084_;
  wire _16085_;
  wire _16086_;
  wire _16087_;
  wire _16088_;
  wire _16089_;
  wire _16090_;
  wire _16091_;
  wire _16092_;
  wire _16093_;
  wire _16094_;
  wire _16095_;
  wire _16096_;
  wire _16097_;
  wire _16098_;
  wire _16099_;
  wire _16100_;
  wire _16101_;
  wire _16102_;
  wire _16103_;
  wire _16104_;
  wire _16105_;
  wire _16106_;
  wire _16107_;
  wire _16108_;
  wire _16109_;
  wire _16110_;
  wire _16111_;
  wire _16112_;
  wire _16113_;
  wire _16114_;
  wire _16115_;
  wire _16116_;
  wire _16117_;
  wire _16118_;
  wire _16119_;
  wire _16120_;
  wire _16121_;
  wire _16122_;
  wire _16123_;
  wire _16124_;
  wire _16125_;
  wire _16126_;
  wire _16127_;
  wire _16128_;
  wire _16129_;
  wire _16130_;
  wire _16131_;
  wire _16132_;
  wire _16133_;
  wire _16134_;
  wire _16135_;
  wire _16136_;
  wire _16137_;
  wire _16138_;
  wire _16139_;
  wire _16140_;
  wire _16141_;
  wire _16142_;
  wire _16143_;
  wire _16144_;
  wire _16145_;
  wire _16146_;
  wire _16147_;
  wire _16148_;
  wire _16149_;
  wire _16150_;
  wire _16151_;
  wire _16152_;
  wire _16153_;
  wire _16154_;
  wire _16155_;
  wire _16156_;
  wire _16157_;
  wire _16158_;
  wire _16159_;
  wire _16160_;
  wire _16161_;
  wire _16162_;
  wire _16163_;
  wire _16164_;
  wire _16165_;
  wire _16166_;
  wire _16167_;
  wire _16168_;
  wire _16169_;
  wire _16170_;
  wire _16171_;
  wire _16172_;
  wire _16173_;
  wire _16174_;
  wire _16175_;
  wire _16176_;
  wire _16177_;
  wire _16178_;
  wire _16179_;
  wire _16180_;
  wire _16181_;
  wire _16182_;
  wire _16183_;
  wire _16184_;
  wire _16185_;
  wire _16186_;
  wire _16187_;
  wire _16188_;
  wire _16189_;
  wire _16190_;
  wire _16191_;
  wire _16192_;
  wire _16193_;
  wire _16194_;
  wire _16195_;
  wire _16196_;
  wire _16197_;
  wire _16198_;
  wire _16199_;
  wire _16200_;
  wire _16201_;
  wire _16202_;
  wire _16203_;
  wire _16204_;
  wire _16205_;
  wire _16206_;
  wire _16207_;
  wire _16208_;
  wire _16209_;
  wire _16210_;
  wire _16211_;
  wire _16212_;
  wire _16213_;
  wire _16214_;
  wire _16215_;
  wire _16216_;
  wire _16217_;
  wire _16218_;
  wire _16219_;
  wire _16220_;
  wire _16221_;
  wire _16222_;
  wire _16223_;
  wire _16224_;
  wire _16225_;
  wire _16226_;
  wire _16227_;
  wire _16228_;
  wire _16229_;
  wire _16230_;
  wire _16231_;
  wire _16232_;
  wire _16233_;
  wire _16234_;
  wire _16235_;
  wire _16236_;
  wire _16237_;
  wire _16238_;
  wire _16239_;
  wire _16240_;
  wire _16241_;
  wire _16242_;
  wire _16243_;
  wire _16244_;
  wire _16245_;
  wire _16246_;
  wire _16247_;
  wire _16248_;
  wire _16249_;
  wire _16250_;
  wire _16251_;
  wire _16252_;
  wire _16253_;
  wire _16254_;
  wire _16255_;
  wire _16256_;
  wire _16257_;
  wire _16258_;
  wire _16259_;
  wire _16260_;
  wire _16261_;
  wire _16262_;
  wire _16263_;
  wire _16264_;
  wire _16265_;
  wire _16266_;
  wire _16267_;
  wire _16268_;
  wire _16269_;
  wire _16270_;
  wire _16271_;
  wire _16272_;
  wire _16273_;
  wire _16274_;
  wire _16275_;
  wire _16276_;
  wire _16277_;
  wire _16278_;
  wire _16279_;
  wire _16280_;
  wire _16281_;
  wire _16282_;
  wire _16283_;
  wire _16284_;
  wire _16285_;
  wire _16286_;
  wire _16287_;
  wire _16288_;
  wire _16289_;
  wire _16290_;
  wire _16291_;
  wire _16292_;
  wire _16293_;
  wire _16294_;
  wire _16295_;
  wire _16296_;
  wire _16297_;
  wire _16298_;
  wire _16299_;
  wire _16300_;
  wire _16301_;
  wire _16302_;
  wire _16303_;
  wire _16304_;
  wire _16305_;
  wire _16306_;
  wire _16307_;
  wire _16308_;
  wire _16309_;
  wire _16310_;
  wire _16311_;
  wire _16312_;
  wire _16313_;
  wire _16314_;
  wire _16315_;
  wire _16316_;
  wire _16317_;
  wire _16318_;
  wire _16319_;
  wire _16320_;
  wire _16321_;
  wire _16322_;
  wire _16323_;
  wire _16324_;
  wire _16325_;
  wire _16326_;
  wire _16327_;
  wire _16328_;
  wire _16329_;
  wire _16330_;
  wire _16331_;
  wire _16332_;
  wire _16333_;
  wire _16334_;
  wire _16335_;
  wire _16336_;
  wire _16337_;
  wire _16338_;
  wire _16339_;
  wire _16340_;
  wire _16341_;
  wire _16342_;
  wire _16343_;
  wire _16344_;
  wire _16345_;
  wire _16346_;
  wire _16347_;
  wire _16348_;
  wire _16349_;
  wire _16350_;
  wire _16351_;
  wire _16352_;
  wire _16353_;
  wire _16354_;
  wire _16355_;
  wire _16356_;
  wire _16357_;
  wire _16358_;
  wire _16359_;
  wire _16360_;
  wire _16361_;
  wire _16362_;
  wire _16363_;
  wire _16364_;
  wire _16365_;
  wire _16366_;
  wire _16367_;
  wire _16368_;
  wire _16369_;
  wire _16370_;
  wire _16371_;
  wire _16372_;
  wire _16373_;
  wire _16374_;
  wire _16375_;
  wire _16376_;
  wire _16377_;
  wire _16378_;
  wire _16379_;
  wire _16380_;
  wire _16381_;
  wire _16382_;
  wire _16383_;
  wire _16384_;
  wire _16385_;
  wire _16386_;
  wire _16387_;
  wire _16388_;
  wire _16389_;
  wire _16390_;
  wire _16391_;
  wire _16392_;
  wire _16393_;
  wire _16394_;
  wire _16395_;
  wire _16396_;
  wire _16397_;
  wire _16398_;
  wire _16399_;
  wire _16400_;
  wire _16401_;
  wire _16402_;
  wire _16403_;
  wire _16404_;
  wire _16405_;
  wire _16406_;
  wire _16407_;
  wire _16408_;
  wire _16409_;
  wire _16410_;
  wire _16411_;
  wire _16412_;
  wire _16413_;
  wire _16414_;
  wire _16415_;
  wire _16416_;
  wire _16417_;
  wire _16418_;
  wire _16419_;
  wire _16420_;
  wire _16421_;
  wire _16422_;
  wire _16423_;
  wire _16424_;
  wire _16425_;
  wire _16426_;
  wire _16427_;
  wire _16428_;
  wire _16429_;
  wire _16430_;
  wire _16431_;
  wire _16432_;
  wire _16433_;
  wire _16434_;
  wire _16435_;
  wire _16436_;
  wire _16437_;
  wire _16438_;
  wire _16439_;
  wire _16440_;
  wire _16441_;
  wire _16442_;
  wire _16443_;
  wire _16444_;
  wire _16445_;
  wire _16446_;
  wire _16447_;
  wire _16448_;
  wire _16449_;
  wire _16450_;
  wire _16451_;
  wire _16452_;
  wire _16453_;
  wire _16454_;
  wire _16455_;
  wire _16456_;
  wire _16457_;
  wire _16458_;
  wire _16459_;
  wire _16460_;
  wire _16461_;
  wire _16462_;
  wire _16463_;
  wire _16464_;
  wire _16465_;
  wire _16466_;
  wire _16467_;
  wire _16468_;
  wire _16469_;
  wire _16470_;
  wire _16471_;
  wire _16472_;
  wire _16473_;
  wire _16474_;
  wire _16475_;
  wire _16476_;
  wire _16477_;
  wire _16478_;
  wire _16479_;
  wire _16480_;
  wire _16481_;
  wire _16482_;
  wire _16483_;
  wire _16484_;
  wire _16485_;
  wire _16486_;
  wire _16487_;
  wire _16488_;
  wire _16489_;
  wire _16490_;
  wire _16491_;
  wire _16492_;
  wire _16493_;
  wire _16494_;
  wire _16495_;
  wire _16496_;
  wire _16497_;
  wire _16498_;
  wire _16499_;
  wire _16500_;
  wire _16501_;
  wire _16502_;
  wire _16503_;
  wire _16504_;
  wire _16505_;
  wire _16506_;
  wire _16507_;
  wire _16508_;
  wire _16509_;
  wire _16510_;
  wire _16511_;
  wire _16512_;
  wire _16513_;
  wire _16514_;
  wire _16515_;
  wire _16516_;
  wire _16517_;
  wire _16518_;
  wire _16519_;
  wire _16520_;
  wire _16521_;
  wire _16522_;
  wire _16523_;
  wire _16524_;
  wire _16525_;
  wire _16526_;
  wire _16527_;
  wire _16528_;
  wire _16529_;
  wire _16530_;
  wire _16531_;
  wire _16532_;
  wire _16533_;
  wire _16534_;
  wire _16535_;
  wire _16536_;
  wire _16537_;
  wire _16538_;
  wire _16539_;
  wire _16540_;
  wire _16541_;
  wire _16542_;
  wire _16543_;
  wire _16544_;
  wire _16545_;
  wire _16546_;
  wire _16547_;
  wire _16548_;
  wire _16549_;
  wire _16550_;
  wire _16551_;
  wire _16552_;
  wire _16553_;
  wire _16554_;
  wire _16555_;
  wire _16556_;
  wire _16557_;
  wire _16558_;
  wire _16559_;
  wire _16560_;
  wire _16561_;
  wire _16562_;
  wire _16563_;
  wire _16564_;
  wire _16565_;
  wire _16566_;
  wire _16567_;
  wire _16568_;
  wire _16569_;
  wire _16570_;
  wire _16571_;
  wire _16572_;
  wire _16573_;
  wire _16574_;
  wire _16575_;
  wire _16576_;
  wire _16577_;
  wire _16578_;
  wire _16579_;
  wire _16580_;
  wire _16581_;
  wire _16582_;
  wire _16583_;
  wire _16584_;
  wire _16585_;
  wire _16586_;
  wire _16587_;
  wire _16588_;
  wire _16589_;
  wire _16590_;
  wire _16591_;
  wire _16592_;
  wire _16593_;
  wire _16594_;
  wire _16595_;
  wire _16596_;
  wire _16597_;
  wire _16598_;
  wire _16599_;
  wire _16600_;
  wire _16601_;
  wire _16602_;
  wire _16603_;
  wire _16604_;
  wire _16605_;
  wire _16606_;
  wire _16607_;
  wire _16608_;
  wire _16609_;
  wire _16610_;
  wire _16611_;
  wire _16612_;
  wire _16613_;
  wire _16614_;
  wire _16615_;
  wire _16616_;
  wire _16617_;
  wire _16618_;
  wire _16619_;
  wire _16620_;
  wire _16621_;
  wire _16622_;
  wire _16623_;
  wire _16624_;
  wire _16625_;
  wire _16626_;
  wire _16627_;
  wire _16628_;
  wire _16629_;
  wire _16630_;
  wire _16631_;
  wire _16632_;
  wire _16633_;
  wire _16634_;
  wire _16635_;
  wire _16636_;
  wire _16637_;
  wire _16638_;
  wire _16639_;
  wire _16640_;
  wire _16641_;
  wire _16642_;
  wire _16643_;
  wire _16644_;
  wire _16645_;
  wire _16646_;
  wire _16647_;
  wire _16648_;
  wire _16649_;
  wire _16650_;
  wire _16651_;
  wire _16652_;
  wire _16653_;
  wire _16654_;
  wire _16655_;
  wire _16656_;
  wire _16657_;
  wire _16658_;
  wire _16659_;
  wire _16660_;
  wire _16661_;
  wire _16662_;
  wire _16663_;
  wire _16664_;
  wire _16665_;
  wire _16666_;
  wire _16667_;
  wire _16668_;
  wire _16669_;
  wire _16670_;
  wire _16671_;
  wire _16672_;
  wire _16673_;
  wire _16674_;
  wire _16675_;
  wire _16676_;
  wire _16677_;
  wire _16678_;
  wire _16679_;
  wire _16680_;
  wire _16681_;
  wire _16682_;
  wire _16683_;
  wire _16684_;
  wire _16685_;
  wire _16686_;
  wire _16687_;
  wire _16688_;
  wire _16689_;
  wire _16690_;
  wire _16691_;
  wire _16692_;
  wire _16693_;
  wire _16694_;
  wire _16695_;
  wire _16696_;
  wire _16697_;
  wire _16698_;
  wire _16699_;
  wire _16700_;
  wire _16701_;
  wire _16702_;
  wire _16703_;
  wire _16704_;
  wire _16705_;
  wire _16706_;
  wire _16707_;
  wire _16708_;
  wire _16709_;
  wire _16710_;
  wire _16711_;
  wire _16712_;
  wire _16713_;
  wire _16714_;
  wire _16715_;
  wire _16716_;
  wire _16717_;
  wire _16718_;
  wire _16719_;
  wire _16720_;
  wire _16721_;
  wire _16722_;
  wire _16723_;
  wire _16724_;
  wire _16725_;
  wire _16726_;
  wire _16727_;
  wire _16728_;
  wire _16729_;
  wire _16730_;
  wire _16731_;
  wire _16732_;
  wire _16733_;
  wire _16734_;
  wire _16735_;
  wire _16736_;
  wire _16737_;
  wire _16738_;
  wire _16739_;
  wire _16740_;
  wire _16741_;
  wire _16742_;
  wire _16743_;
  wire _16744_;
  wire _16745_;
  wire _16746_;
  wire _16747_;
  wire _16748_;
  wire _16749_;
  wire _16750_;
  wire _16751_;
  wire _16752_;
  wire _16753_;
  wire _16754_;
  wire _16755_;
  wire _16756_;
  wire _16757_;
  wire _16758_;
  wire _16759_;
  wire _16760_;
  wire _16761_;
  wire _16762_;
  wire _16763_;
  wire _16764_;
  wire _16765_;
  wire _16766_;
  wire _16767_;
  wire _16768_;
  wire _16769_;
  wire _16770_;
  wire _16771_;
  wire _16772_;
  wire _16773_;
  wire _16774_;
  wire _16775_;
  wire _16776_;
  wire _16777_;
  wire _16778_;
  wire _16779_;
  wire _16780_;
  wire _16781_;
  wire _16782_;
  wire _16783_;
  wire _16784_;
  wire _16785_;
  wire _16786_;
  wire _16787_;
  wire _16788_;
  wire _16789_;
  wire _16790_;
  wire _16791_;
  wire _16792_;
  wire _16793_;
  wire _16794_;
  wire _16795_;
  wire _16796_;
  wire _16797_;
  wire _16798_;
  wire _16799_;
  wire _16800_;
  wire _16801_;
  wire _16802_;
  wire _16803_;
  wire _16804_;
  wire _16805_;
  wire _16806_;
  wire _16807_;
  wire _16808_;
  wire _16809_;
  wire _16810_;
  wire _16811_;
  wire _16812_;
  wire _16813_;
  wire _16814_;
  wire _16815_;
  wire _16816_;
  wire _16817_;
  wire _16818_;
  wire _16819_;
  wire _16820_;
  wire _16821_;
  wire _16822_;
  wire _16823_;
  wire _16824_;
  wire _16825_;
  wire _16826_;
  wire _16827_;
  wire _16828_;
  wire _16829_;
  wire _16830_;
  wire _16831_;
  wire _16832_;
  wire _16833_;
  wire _16834_;
  wire _16835_;
  wire _16836_;
  wire _16837_;
  wire _16838_;
  wire _16839_;
  wire _16840_;
  wire _16841_;
  wire _16842_;
  wire _16843_;
  wire _16844_;
  wire _16845_;
  wire _16846_;
  wire _16847_;
  wire _16848_;
  wire _16849_;
  wire _16850_;
  wire _16851_;
  wire _16852_;
  wire _16853_;
  wire _16854_;
  wire _16855_;
  wire _16856_;
  wire _16857_;
  wire _16858_;
  wire _16859_;
  wire _16860_;
  wire _16861_;
  wire _16862_;
  wire _16863_;
  wire _16864_;
  wire _16865_;
  wire _16866_;
  wire _16867_;
  wire _16868_;
  wire _16869_;
  wire _16870_;
  wire _16871_;
  wire _16872_;
  wire _16873_;
  wire _16874_;
  wire _16875_;
  wire _16876_;
  wire _16877_;
  wire _16878_;
  wire _16879_;
  wire _16880_;
  wire _16881_;
  wire _16882_;
  wire _16883_;
  wire _16884_;
  wire _16885_;
  wire _16886_;
  wire _16887_;
  wire _16888_;
  wire _16889_;
  wire _16890_;
  wire _16891_;
  wire _16892_;
  wire _16893_;
  wire _16894_;
  wire _16895_;
  wire _16896_;
  wire _16897_;
  wire _16898_;
  wire _16899_;
  wire _16900_;
  wire _16901_;
  wire _16902_;
  wire _16903_;
  wire _16904_;
  wire _16905_;
  wire _16906_;
  wire _16907_;
  wire _16908_;
  wire _16909_;
  wire _16910_;
  wire _16911_;
  wire _16912_;
  wire _16913_;
  wire _16914_;
  wire _16915_;
  wire _16916_;
  wire _16917_;
  wire _16918_;
  wire _16919_;
  wire _16920_;
  wire _16921_;
  wire _16922_;
  wire _16923_;
  wire _16924_;
  wire _16925_;
  wire _16926_;
  wire _16927_;
  wire _16928_;
  wire _16929_;
  wire _16930_;
  wire _16931_;
  wire _16932_;
  wire _16933_;
  wire _16934_;
  wire _16935_;
  wire _16936_;
  wire _16937_;
  wire _16938_;
  wire _16939_;
  wire _16940_;
  wire _16941_;
  wire _16942_;
  wire _16943_;
  wire _16944_;
  wire _16945_;
  wire _16946_;
  wire _16947_;
  wire _16948_;
  wire _16949_;
  wire _16950_;
  wire _16951_;
  wire _16952_;
  wire _16953_;
  wire _16954_;
  wire _16955_;
  wire _16956_;
  wire _16957_;
  wire _16958_;
  wire _16959_;
  wire _16960_;
  wire _16961_;
  wire _16962_;
  wire _16963_;
  wire _16964_;
  wire _16965_;
  wire _16966_;
  wire _16967_;
  wire _16968_;
  wire _16969_;
  wire _16970_;
  wire _16971_;
  wire _16972_;
  wire _16973_;
  wire _16974_;
  wire _16975_;
  wire _16976_;
  wire _16977_;
  wire _16978_;
  wire _16979_;
  wire _16980_;
  wire _16981_;
  wire _16982_;
  wire _16983_;
  wire _16984_;
  wire _16985_;
  wire _16986_;
  wire _16987_;
  wire _16988_;
  wire _16989_;
  wire _16990_;
  wire _16991_;
  wire _16992_;
  wire _16993_;
  wire _16994_;
  wire _16995_;
  wire _16996_;
  wire _16997_;
  wire _16998_;
  wire _16999_;
  wire _17000_;
  wire _17001_;
  wire _17002_;
  wire _17003_;
  wire _17004_;
  wire _17005_;
  wire _17006_;
  wire _17007_;
  wire _17008_;
  wire _17009_;
  wire _17010_;
  wire _17011_;
  wire _17012_;
  wire _17013_;
  wire _17014_;
  wire _17015_;
  wire _17016_;
  wire _17017_;
  wire _17018_;
  wire _17019_;
  wire _17020_;
  wire _17021_;
  wire _17022_;
  wire _17023_;
  wire _17024_;
  wire _17025_;
  wire _17026_;
  wire _17027_;
  wire _17028_;
  wire _17029_;
  wire _17030_;
  wire _17031_;
  wire _17032_;
  wire _17033_;
  wire _17034_;
  wire _17035_;
  wire _17036_;
  wire _17037_;
  wire _17038_;
  wire _17039_;
  wire _17040_;
  wire _17041_;
  wire _17042_;
  wire _17043_;
  wire _17044_;
  wire _17045_;
  wire _17046_;
  wire _17047_;
  wire _17048_;
  wire _17049_;
  wire _17050_;
  wire _17051_;
  wire _17052_;
  wire _17053_;
  wire _17054_;
  wire _17055_;
  wire _17056_;
  wire _17057_;
  wire _17058_;
  wire _17059_;
  wire _17060_;
  wire _17061_;
  wire _17062_;
  wire _17063_;
  wire _17064_;
  wire _17065_;
  wire _17066_;
  wire _17067_;
  wire _17068_;
  wire _17069_;
  wire _17070_;
  wire _17071_;
  wire _17072_;
  wire _17073_;
  wire _17074_;
  wire _17075_;
  wire _17076_;
  wire _17077_;
  wire _17078_;
  wire _17079_;
  wire _17080_;
  wire _17081_;
  wire _17082_;
  wire _17083_;
  wire _17084_;
  wire _17085_;
  wire _17086_;
  wire _17087_;
  wire _17088_;
  wire _17089_;
  wire _17090_;
  wire _17091_;
  wire _17092_;
  wire _17093_;
  wire _17094_;
  wire _17095_;
  wire _17096_;
  wire _17097_;
  wire _17098_;
  wire _17099_;
  wire _17100_;
  wire _17101_;
  wire _17102_;
  wire _17103_;
  wire _17104_;
  wire _17105_;
  wire _17106_;
  wire _17107_;
  wire _17108_;
  wire _17109_;
  wire _17110_;
  wire _17111_;
  wire _17112_;
  wire _17113_;
  wire _17114_;
  wire _17115_;
  wire _17116_;
  wire _17117_;
  wire _17118_;
  wire _17119_;
  wire _17120_;
  wire _17121_;
  wire _17122_;
  wire _17123_;
  wire _17124_;
  wire _17125_;
  wire _17126_;
  wire _17127_;
  wire _17128_;
  wire _17129_;
  wire _17130_;
  wire _17131_;
  wire _17132_;
  wire _17133_;
  wire _17134_;
  wire _17135_;
  wire _17136_;
  wire _17137_;
  wire _17138_;
  wire _17139_;
  wire _17140_;
  wire _17141_;
  wire _17142_;
  wire _17143_;
  wire _17144_;
  wire _17145_;
  wire _17146_;
  wire _17147_;
  wire _17148_;
  wire _17149_;
  wire _17150_;
  wire _17151_;
  wire _17152_;
  wire _17153_;
  wire _17154_;
  wire _17155_;
  wire _17156_;
  wire _17157_;
  wire _17158_;
  wire _17159_;
  wire _17160_;
  wire _17161_;
  wire _17162_;
  wire _17163_;
  wire _17164_;
  wire _17165_;
  wire _17166_;
  wire _17167_;
  wire _17168_;
  wire _17169_;
  wire _17170_;
  wire _17171_;
  wire _17172_;
  wire _17173_;
  wire _17174_;
  wire _17175_;
  wire _17176_;
  wire _17177_;
  wire _17178_;
  wire _17179_;
  wire _17180_;
  wire _17181_;
  wire _17182_;
  wire _17183_;
  wire _17184_;
  wire _17185_;
  wire _17186_;
  wire _17187_;
  wire _17188_;
  wire _17189_;
  wire _17190_;
  wire _17191_;
  wire _17192_;
  wire _17193_;
  wire _17194_;
  wire _17195_;
  wire _17196_;
  wire _17197_;
  wire _17198_;
  wire _17199_;
  wire _17200_;
  wire _17201_;
  wire _17202_;
  wire _17203_;
  wire _17204_;
  wire _17205_;
  wire _17206_;
  wire _17207_;
  wire _17208_;
  wire _17209_;
  wire _17210_;
  wire _17211_;
  wire _17212_;
  wire _17213_;
  wire _17214_;
  wire _17215_;
  wire _17216_;
  wire _17217_;
  wire _17218_;
  wire _17219_;
  wire _17220_;
  wire _17221_;
  wire _17222_;
  wire _17223_;
  wire _17224_;
  wire _17225_;
  wire _17226_;
  wire _17227_;
  wire _17228_;
  wire _17229_;
  wire _17230_;
  wire _17231_;
  wire _17232_;
  wire _17233_;
  wire _17234_;
  wire _17235_;
  wire _17236_;
  wire _17237_;
  wire _17238_;
  wire _17239_;
  wire _17240_;
  wire _17241_;
  wire _17242_;
  wire _17243_;
  wire _17244_;
  wire _17245_;
  wire _17246_;
  wire _17247_;
  wire _17248_;
  wire _17249_;
  wire _17250_;
  wire _17251_;
  wire _17252_;
  wire _17253_;
  wire _17254_;
  wire _17255_;
  wire _17256_;
  wire _17257_;
  wire _17258_;
  wire _17259_;
  wire _17260_;
  wire _17261_;
  wire _17262_;
  wire _17263_;
  wire _17264_;
  wire _17265_;
  wire _17266_;
  wire _17267_;
  wire _17268_;
  wire _17269_;
  wire _17270_;
  wire _17271_;
  wire _17272_;
  wire _17273_;
  wire _17274_;
  wire _17275_;
  wire _17276_;
  wire _17277_;
  wire _17278_;
  wire _17279_;
  wire _17280_;
  wire _17281_;
  wire _17282_;
  wire _17283_;
  wire _17284_;
  wire _17285_;
  wire _17286_;
  wire _17287_;
  wire _17288_;
  wire _17289_;
  wire _17290_;
  wire _17291_;
  wire _17292_;
  wire _17293_;
  wire _17294_;
  wire _17295_;
  wire _17296_;
  wire _17297_;
  wire _17298_;
  wire _17299_;
  wire _17300_;
  wire _17301_;
  wire _17302_;
  wire _17303_;
  wire _17304_;
  wire _17305_;
  wire _17306_;
  wire _17307_;
  wire _17308_;
  wire _17309_;
  wire _17310_;
  wire _17311_;
  wire _17312_;
  wire _17313_;
  wire _17314_;
  wire _17315_;
  wire _17316_;
  wire _17317_;
  wire _17318_;
  wire _17319_;
  wire _17320_;
  wire _17321_;
  wire _17322_;
  wire _17323_;
  wire _17324_;
  wire _17325_;
  wire _17326_;
  wire _17327_;
  wire _17328_;
  wire _17329_;
  wire _17330_;
  wire _17331_;
  wire _17332_;
  wire _17333_;
  wire _17334_;
  wire _17335_;
  wire _17336_;
  wire _17337_;
  wire _17338_;
  wire _17339_;
  wire _17340_;
  wire _17341_;
  wire _17342_;
  wire _17343_;
  wire _17344_;
  wire _17345_;
  wire _17346_;
  wire _17347_;
  wire _17348_;
  wire _17349_;
  wire _17350_;
  wire _17351_;
  wire _17352_;
  wire _17353_;
  wire _17354_;
  wire _17355_;
  wire _17356_;
  wire _17357_;
  wire _17358_;
  wire _17359_;
  wire _17360_;
  wire _17361_;
  wire _17362_;
  wire _17363_;
  wire _17364_;
  wire _17365_;
  wire _17366_;
  wire _17367_;
  wire _17368_;
  wire _17369_;
  wire _17370_;
  wire _17371_;
  wire _17372_;
  wire _17373_;
  wire _17374_;
  wire _17375_;
  wire _17376_;
  wire _17377_;
  wire _17378_;
  wire _17379_;
  wire _17380_;
  wire _17381_;
  wire _17382_;
  wire _17383_;
  wire _17384_;
  wire _17385_;
  wire _17386_;
  wire _17387_;
  wire _17388_;
  wire _17389_;
  wire _17390_;
  wire _17391_;
  wire _17392_;
  wire _17393_;
  wire _17394_;
  wire _17395_;
  wire _17396_;
  wire _17397_;
  wire _17398_;
  wire _17399_;
  wire _17400_;
  wire _17401_;
  wire _17402_;
  wire _17403_;
  wire _17404_;
  wire _17405_;
  wire _17406_;
  wire _17407_;
  wire _17408_;
  wire _17409_;
  wire _17410_;
  wire _17411_;
  wire _17412_;
  wire _17413_;
  wire _17414_;
  wire _17415_;
  wire _17416_;
  wire _17417_;
  wire _17418_;
  wire _17419_;
  wire _17420_;
  wire _17421_;
  wire _17422_;
  wire _17423_;
  wire _17424_;
  wire _17425_;
  wire _17426_;
  wire _17427_;
  wire _17428_;
  wire _17429_;
  wire _17430_;
  wire _17431_;
  wire _17432_;
  wire _17433_;
  wire _17434_;
  wire _17435_;
  wire _17436_;
  wire _17437_;
  wire _17438_;
  wire _17439_;
  wire _17440_;
  wire _17441_;
  wire _17442_;
  wire _17443_;
  wire _17444_;
  wire _17445_;
  wire _17446_;
  wire _17447_;
  wire _17448_;
  wire _17449_;
  wire _17450_;
  wire _17451_;
  wire _17452_;
  wire _17453_;
  wire _17454_;
  wire _17455_;
  wire _17456_;
  wire _17457_;
  wire _17458_;
  wire _17459_;
  wire _17460_;
  wire _17461_;
  wire _17462_;
  wire _17463_;
  wire _17464_;
  wire _17465_;
  wire _17466_;
  wire _17467_;
  wire _17468_;
  wire _17469_;
  wire _17470_;
  wire _17471_;
  wire _17472_;
  wire _17473_;
  wire _17474_;
  wire _17475_;
  wire _17476_;
  wire _17477_;
  wire _17478_;
  wire _17479_;
  wire _17480_;
  wire _17481_;
  wire _17482_;
  wire _17483_;
  wire _17484_;
  wire _17485_;
  wire _17486_;
  wire _17487_;
  wire _17488_;
  wire _17489_;
  wire _17490_;
  wire _17491_;
  wire _17492_;
  wire _17493_;
  wire _17494_;
  wire _17495_;
  wire _17496_;
  wire _17497_;
  wire _17498_;
  wire _17499_;
  wire _17500_;
  wire _17501_;
  wire _17502_;
  wire _17503_;
  wire _17504_;
  wire _17505_;
  wire _17506_;
  wire _17507_;
  wire _17508_;
  wire _17509_;
  wire _17510_;
  wire _17511_;
  wire _17512_;
  wire _17513_;
  wire _17514_;
  wire _17515_;
  wire _17516_;
  wire _17517_;
  wire _17518_;
  wire _17519_;
  wire _17520_;
  wire _17521_;
  wire _17522_;
  wire _17523_;
  wire _17524_;
  wire _17525_;
  wire _17526_;
  wire _17527_;
  wire _17528_;
  wire _17529_;
  wire _17530_;
  wire _17531_;
  wire _17532_;
  wire _17533_;
  wire _17534_;
  wire _17535_;
  wire _17536_;
  wire _17537_;
  wire _17538_;
  wire _17539_;
  wire _17540_;
  wire _17541_;
  wire _17542_;
  wire _17543_;
  wire _17544_;
  wire _17545_;
  wire _17546_;
  wire _17547_;
  wire _17548_;
  wire _17549_;
  wire _17550_;
  wire _17551_;
  wire _17552_;
  wire _17553_;
  wire _17554_;
  wire _17555_;
  wire _17556_;
  wire _17557_;
  wire _17558_;
  wire _17559_;
  wire _17560_;
  wire _17561_;
  wire _17562_;
  wire _17563_;
  wire _17564_;
  wire _17565_;
  wire _17566_;
  wire _17567_;
  wire _17568_;
  wire _17569_;
  wire _17570_;
  wire _17571_;
  wire _17572_;
  wire _17573_;
  wire _17574_;
  wire _17575_;
  wire _17576_;
  wire _17577_;
  wire _17578_;
  wire _17579_;
  wire _17580_;
  wire _17581_;
  wire _17582_;
  wire _17583_;
  wire _17584_;
  wire _17585_;
  wire _17586_;
  wire _17587_;
  wire _17588_;
  wire _17589_;
  wire _17590_;
  wire _17591_;
  wire _17592_;
  wire _17593_;
  wire _17594_;
  wire _17595_;
  wire _17596_;
  wire _17597_;
  wire _17598_;
  wire _17599_;
  wire _17600_;
  wire _17601_;
  wire _17602_;
  wire _17603_;
  wire _17604_;
  wire _17605_;
  wire _17606_;
  wire _17607_;
  wire _17608_;
  wire _17609_;
  wire _17610_;
  wire _17611_;
  wire _17612_;
  wire _17613_;
  wire _17614_;
  wire _17615_;
  wire _17616_;
  wire _17617_;
  wire _17618_;
  wire _17619_;
  wire _17620_;
  wire _17621_;
  wire _17622_;
  wire _17623_;
  wire _17624_;
  wire _17625_;
  wire _17626_;
  wire _17627_;
  wire _17628_;
  wire _17629_;
  wire _17630_;
  wire _17631_;
  wire _17632_;
  wire _17633_;
  wire _17634_;
  wire _17635_;
  wire _17636_;
  wire _17637_;
  wire _17638_;
  wire _17639_;
  wire _17640_;
  wire _17641_;
  wire _17642_;
  wire _17643_;
  wire _17644_;
  wire _17645_;
  wire _17646_;
  wire _17647_;
  wire _17648_;
  wire _17649_;
  wire _17650_;
  wire _17651_;
  wire _17652_;
  wire _17653_;
  wire _17654_;
  wire _17655_;
  wire _17656_;
  wire _17657_;
  wire _17658_;
  wire _17659_;
  wire _17660_;
  wire _17661_;
  wire _17662_;
  wire _17663_;
  wire _17664_;
  wire _17665_;
  wire _17666_;
  wire _17667_;
  wire _17668_;
  wire _17669_;
  wire _17670_;
  wire _17671_;
  wire _17672_;
  wire _17673_;
  wire _17674_;
  wire _17675_;
  wire _17676_;
  wire _17677_;
  wire _17678_;
  wire _17679_;
  wire _17680_;
  wire _17681_;
  wire _17682_;
  wire _17683_;
  wire _17684_;
  wire _17685_;
  wire _17686_;
  wire _17687_;
  wire _17688_;
  wire _17689_;
  wire _17690_;
  wire _17691_;
  wire _17692_;
  wire _17693_;
  wire _17694_;
  wire _17695_;
  wire _17696_;
  wire _17697_;
  wire _17698_;
  wire _17699_;
  wire _17700_;
  wire _17701_;
  wire _17702_;
  wire _17703_;
  wire _17704_;
  wire _17705_;
  wire _17706_;
  wire _17707_;
  wire _17708_;
  wire _17709_;
  wire _17710_;
  wire _17711_;
  wire _17712_;
  wire _17713_;
  wire _17714_;
  wire _17715_;
  wire _17716_;
  wire _17717_;
  wire _17718_;
  wire _17719_;
  wire _17720_;
  wire _17721_;
  wire _17722_;
  wire _17723_;
  wire _17724_;
  wire _17725_;
  wire _17726_;
  wire _17727_;
  wire _17728_;
  wire _17729_;
  wire _17730_;
  wire _17731_;
  wire _17732_;
  wire _17733_;
  wire _17734_;
  wire _17735_;
  wire _17736_;
  wire _17737_;
  wire _17738_;
  wire _17739_;
  wire _17740_;
  wire _17741_;
  wire _17742_;
  wire _17743_;
  wire _17744_;
  wire _17745_;
  wire _17746_;
  wire _17747_;
  wire _17748_;
  wire _17749_;
  wire _17750_;
  wire _17751_;
  wire _17752_;
  wire _17753_;
  wire _17754_;
  wire _17755_;
  wire _17756_;
  wire _17757_;
  wire _17758_;
  wire _17759_;
  wire _17760_;
  wire _17761_;
  wire _17762_;
  wire _17763_;
  wire _17764_;
  wire _17765_;
  wire _17766_;
  wire _17767_;
  wire _17768_;
  wire _17769_;
  wire _17770_;
  wire _17771_;
  wire _17772_;
  wire _17773_;
  wire _17774_;
  wire _17775_;
  wire _17776_;
  wire _17777_;
  wire _17778_;
  wire _17779_;
  wire _17780_;
  wire _17781_;
  wire _17782_;
  wire _17783_;
  wire _17784_;
  wire _17785_;
  wire _17786_;
  wire _17787_;
  wire _17788_;
  wire _17789_;
  wire _17790_;
  wire _17791_;
  wire _17792_;
  wire _17793_;
  wire _17794_;
  wire _17795_;
  wire _17796_;
  wire _17797_;
  wire _17798_;
  wire _17799_;
  wire _17800_;
  wire _17801_;
  wire _17802_;
  wire _17803_;
  wire _17804_;
  wire _17805_;
  wire _17806_;
  wire _17807_;
  wire _17808_;
  wire _17809_;
  wire _17810_;
  wire _17811_;
  wire _17812_;
  wire _17813_;
  wire _17814_;
  wire _17815_;
  wire _17816_;
  wire _17817_;
  wire _17818_;
  wire _17819_;
  wire _17820_;
  wire _17821_;
  wire _17822_;
  wire _17823_;
  wire _17824_;
  wire _17825_;
  wire _17826_;
  wire _17827_;
  wire _17828_;
  wire _17829_;
  wire _17830_;
  wire _17831_;
  wire _17832_;
  wire _17833_;
  wire _17834_;
  wire _17835_;
  wire _17836_;
  wire _17837_;
  wire _17838_;
  wire _17839_;
  wire _17840_;
  wire _17841_;
  wire _17842_;
  wire _17843_;
  wire _17844_;
  wire _17845_;
  wire _17846_;
  wire _17847_;
  wire _17848_;
  wire _17849_;
  wire _17850_;
  wire _17851_;
  wire _17852_;
  wire _17853_;
  wire _17854_;
  wire _17855_;
  wire _17856_;
  wire _17857_;
  wire _17858_;
  wire _17859_;
  wire _17860_;
  wire _17861_;
  wire _17862_;
  wire _17863_;
  wire _17864_;
  wire _17865_;
  wire _17866_;
  wire _17867_;
  wire _17868_;
  wire _17869_;
  wire _17870_;
  wire _17871_;
  wire _17872_;
  wire _17873_;
  wire _17874_;
  wire _17875_;
  wire _17876_;
  wire _17877_;
  wire _17878_;
  wire _17879_;
  wire _17880_;
  wire _17881_;
  wire _17882_;
  wire _17883_;
  wire _17884_;
  wire _17885_;
  wire _17886_;
  wire _17887_;
  wire _17888_;
  wire _17889_;
  wire _17890_;
  wire _17891_;
  wire _17892_;
  wire _17893_;
  wire _17894_;
  wire _17895_;
  wire _17896_;
  wire _17897_;
  wire _17898_;
  wire _17899_;
  wire _17900_;
  wire _17901_;
  wire _17902_;
  wire _17903_;
  wire _17904_;
  wire _17905_;
  wire _17906_;
  wire _17907_;
  wire _17908_;
  wire _17909_;
  wire _17910_;
  wire _17911_;
  wire _17912_;
  wire _17913_;
  wire _17914_;
  wire _17915_;
  wire _17916_;
  wire _17917_;
  wire _17918_;
  wire _17919_;
  wire _17920_;
  wire _17921_;
  wire _17922_;
  wire _17923_;
  wire _17924_;
  wire _17925_;
  wire _17926_;
  wire _17927_;
  wire _17928_;
  wire _17929_;
  wire _17930_;
  wire _17931_;
  wire _17932_;
  wire _17933_;
  wire _17934_;
  wire _17935_;
  wire _17936_;
  wire _17937_;
  wire _17938_;
  wire _17939_;
  wire _17940_;
  wire _17941_;
  wire _17942_;
  wire _17943_;
  wire _17944_;
  wire _17945_;
  wire _17946_;
  wire _17947_;
  wire _17948_;
  wire _17949_;
  wire _17950_;
  wire _17951_;
  wire _17952_;
  wire _17953_;
  wire _17954_;
  wire _17955_;
  wire _17956_;
  wire _17957_;
  wire _17958_;
  wire _17959_;
  wire _17960_;
  wire _17961_;
  wire _17962_;
  wire _17963_;
  wire _17964_;
  wire _17965_;
  wire _17966_;
  wire _17967_;
  wire _17968_;
  wire _17969_;
  wire _17970_;
  wire _17971_;
  wire _17972_;
  wire _17973_;
  wire _17974_;
  wire _17975_;
  wire _17976_;
  wire _17977_;
  wire _17978_;
  wire _17979_;
  wire _17980_;
  wire _17981_;
  wire _17982_;
  wire _17983_;
  wire _17984_;
  wire _17985_;
  wire _17986_;
  wire _17987_;
  wire _17988_;
  wire _17989_;
  wire _17990_;
  wire _17991_;
  wire _17992_;
  wire _17993_;
  wire _17994_;
  wire _17995_;
  wire _17996_;
  wire _17997_;
  wire _17998_;
  wire _17999_;
  wire _18000_;
  wire _18001_;
  wire _18002_;
  wire _18003_;
  wire _18004_;
  wire _18005_;
  wire _18006_;
  wire _18007_;
  wire _18008_;
  wire _18009_;
  wire _18010_;
  wire _18011_;
  wire _18012_;
  wire _18013_;
  wire _18014_;
  wire _18015_;
  wire _18016_;
  wire _18017_;
  wire _18018_;
  wire _18019_;
  wire _18020_;
  wire _18021_;
  wire _18022_;
  wire _18023_;
  wire _18024_;
  wire _18025_;
  wire _18026_;
  wire _18027_;
  wire _18028_;
  wire _18029_;
  wire _18030_;
  wire _18031_;
  wire _18032_;
  wire _18033_;
  wire _18034_;
  wire _18035_;
  wire _18036_;
  wire _18037_;
  wire _18038_;
  wire _18039_;
  wire _18040_;
  wire _18041_;
  wire _18042_;
  wire _18043_;
  wire _18044_;
  wire _18045_;
  wire _18046_;
  wire _18047_;
  wire _18048_;
  wire _18049_;
  wire _18050_;
  wire _18051_;
  wire _18052_;
  wire _18053_;
  wire _18054_;
  wire _18055_;
  wire _18056_;
  wire _18057_;
  wire _18058_;
  wire _18059_;
  wire _18060_;
  wire _18061_;
  wire _18062_;
  wire _18063_;
  wire _18064_;
  wire _18065_;
  wire _18066_;
  wire _18067_;
  wire _18068_;
  wire _18069_;
  wire _18070_;
  wire _18071_;
  wire _18072_;
  wire _18073_;
  wire _18074_;
  wire _18075_;
  wire _18076_;
  wire _18077_;
  wire _18078_;
  wire _18079_;
  wire _18080_;
  wire _18081_;
  wire _18082_;
  wire _18083_;
  wire _18084_;
  wire _18085_;
  wire _18086_;
  wire _18087_;
  wire _18088_;
  wire _18089_;
  wire _18090_;
  wire _18091_;
  wire _18092_;
  wire _18093_;
  wire _18094_;
  wire _18095_;
  wire _18096_;
  wire _18097_;
  wire _18098_;
  wire _18099_;
  wire _18100_;
  wire _18101_;
  wire _18102_;
  wire _18103_;
  wire _18104_;
  wire _18105_;
  wire _18106_;
  wire _18107_;
  wire _18108_;
  wire _18109_;
  wire _18110_;
  wire _18111_;
  wire _18112_;
  wire _18113_;
  wire _18114_;
  wire _18115_;
  wire _18116_;
  wire _18117_;
  wire _18118_;
  wire _18119_;
  wire _18120_;
  wire _18121_;
  wire _18122_;
  wire _18123_;
  wire _18124_;
  wire _18125_;
  wire _18126_;
  wire _18127_;
  wire _18128_;
  wire _18129_;
  wire _18130_;
  wire _18131_;
  wire _18132_;
  wire _18133_;
  wire _18134_;
  wire _18135_;
  wire _18136_;
  wire _18137_;
  wire _18138_;
  wire _18139_;
  wire _18140_;
  wire _18141_;
  wire _18142_;
  wire _18143_;
  wire _18144_;
  wire _18145_;
  wire _18146_;
  wire _18147_;
  wire _18148_;
  wire _18149_;
  wire _18150_;
  wire _18151_;
  wire _18152_;
  wire _18153_;
  wire _18154_;
  wire _18155_;
  wire _18156_;
  wire _18157_;
  wire _18158_;
  wire _18159_;
  wire _18160_;
  wire _18161_;
  wire _18162_;
  wire _18163_;
  wire _18164_;
  wire _18165_;
  wire _18166_;
  wire _18167_;
  wire _18168_;
  wire _18169_;
  wire _18170_;
  wire _18171_;
  wire _18172_;
  wire _18173_;
  wire _18174_;
  wire _18175_;
  wire _18176_;
  wire _18177_;
  wire _18178_;
  wire _18179_;
  wire _18180_;
  wire _18181_;
  wire _18182_;
  wire _18183_;
  wire _18184_;
  wire _18185_;
  wire _18186_;
  wire _18187_;
  wire _18188_;
  wire _18189_;
  wire _18190_;
  wire _18191_;
  wire _18192_;
  wire _18193_;
  wire _18194_;
  wire _18195_;
  wire _18196_;
  wire _18197_;
  wire _18198_;
  wire _18199_;
  wire _18200_;
  wire _18201_;
  wire _18202_;
  wire _18203_;
  wire _18204_;
  wire _18205_;
  wire _18206_;
  wire _18207_;
  wire _18208_;
  wire _18209_;
  wire _18210_;
  wire _18211_;
  wire _18212_;
  wire _18213_;
  wire _18214_;
  wire _18215_;
  wire _18216_;
  wire _18217_;
  wire _18218_;
  wire _18219_;
  wire _18220_;
  wire _18221_;
  wire _18222_;
  wire _18223_;
  wire _18224_;
  wire _18225_;
  wire _18226_;
  wire _18227_;
  wire _18228_;
  wire _18229_;
  wire _18230_;
  wire _18231_;
  wire _18232_;
  wire _18233_;
  wire _18234_;
  wire _18235_;
  wire _18236_;
  wire _18237_;
  wire _18238_;
  wire _18239_;
  wire _18240_;
  wire _18241_;
  wire _18242_;
  wire _18243_;
  wire _18244_;
  wire _18245_;
  wire _18246_;
  wire _18247_;
  wire _18248_;
  wire _18249_;
  wire _18250_;
  wire _18251_;
  wire _18252_;
  wire _18253_;
  wire _18254_;
  wire _18255_;
  wire _18256_;
  wire _18257_;
  wire _18258_;
  wire _18259_;
  wire _18260_;
  wire _18261_;
  wire _18262_;
  wire _18263_;
  wire _18264_;
  wire _18265_;
  wire _18266_;
  wire _18267_;
  wire _18268_;
  wire _18269_;
  wire _18270_;
  wire _18271_;
  wire _18272_;
  wire _18273_;
  wire _18274_;
  wire _18275_;
  wire _18276_;
  wire _18277_;
  wire _18278_;
  wire _18279_;
  wire _18280_;
  wire _18281_;
  wire _18282_;
  wire _18283_;
  wire _18284_;
  wire _18285_;
  wire _18286_;
  wire _18287_;
  wire _18288_;
  wire _18289_;
  wire _18290_;
  wire _18291_;
  wire _18292_;
  wire _18293_;
  wire _18294_;
  wire _18295_;
  wire _18296_;
  wire _18297_;
  wire _18298_;
  wire _18299_;
  wire _18300_;
  wire _18301_;
  wire _18302_;
  wire _18303_;
  wire _18304_;
  wire _18305_;
  wire _18306_;
  wire _18307_;
  wire _18308_;
  wire _18309_;
  wire _18310_;
  wire _18311_;
  wire _18312_;
  wire _18313_;
  wire _18314_;
  wire _18315_;
  wire _18316_;
  wire _18317_;
  wire _18318_;
  wire _18319_;
  wire _18320_;
  wire _18321_;
  wire _18322_;
  wire _18323_;
  wire _18324_;
  wire _18325_;
  wire _18326_;
  wire _18327_;
  wire _18328_;
  wire _18329_;
  wire _18330_;
  wire _18331_;
  wire _18332_;
  wire _18333_;
  wire _18334_;
  wire _18335_;
  wire _18336_;
  wire _18337_;
  wire _18338_;
  wire _18339_;
  wire _18340_;
  wire _18341_;
  wire _18342_;
  wire _18343_;
  wire _18344_;
  wire _18345_;
  wire _18346_;
  wire _18347_;
  wire _18348_;
  wire _18349_;
  wire _18350_;
  wire _18351_;
  wire _18352_;
  wire _18353_;
  wire _18354_;
  wire _18355_;
  wire _18356_;
  wire _18357_;
  wire _18358_;
  wire _18359_;
  wire _18360_;
  wire _18361_;
  wire _18362_;
  wire _18363_;
  wire _18364_;
  wire _18365_;
  wire _18366_;
  wire _18367_;
  wire _18368_;
  wire _18369_;
  wire _18370_;
  wire _18371_;
  wire _18372_;
  wire _18373_;
  wire _18374_;
  wire _18375_;
  wire _18376_;
  wire _18377_;
  wire _18378_;
  wire _18379_;
  wire _18380_;
  wire _18381_;
  wire _18382_;
  wire _18383_;
  wire _18384_;
  wire _18385_;
  wire _18386_;
  wire _18387_;
  wire _18388_;
  wire _18389_;
  wire _18390_;
  wire _18391_;
  wire _18392_;
  wire _18393_;
  wire _18394_;
  wire _18395_;
  wire _18396_;
  wire _18397_;
  wire _18398_;
  wire _18399_;
  wire _18400_;
  wire _18401_;
  wire _18402_;
  wire _18403_;
  wire _18404_;
  wire _18405_;
  wire _18406_;
  wire _18407_;
  wire _18408_;
  wire _18409_;
  wire _18410_;
  wire _18411_;
  wire _18412_;
  wire _18413_;
  wire _18414_;
  wire _18415_;
  wire _18416_;
  wire _18417_;
  wire _18418_;
  wire _18419_;
  wire _18420_;
  wire _18421_;
  wire _18422_;
  wire _18423_;
  wire _18424_;
  wire _18425_;
  wire _18426_;
  wire _18427_;
  wire _18428_;
  wire _18429_;
  wire _18430_;
  wire _18431_;
  wire _18432_;
  wire _18433_;
  wire _18434_;
  wire _18435_;
  wire _18436_;
  wire _18437_;
  wire _18438_;
  wire _18439_;
  wire _18440_;
  wire _18441_;
  wire _18442_;
  wire _18443_;
  wire _18444_;
  wire _18445_;
  wire _18446_;
  wire _18447_;
  wire _18448_;
  wire _18449_;
  wire _18450_;
  wire _18451_;
  wire _18452_;
  wire _18453_;
  wire _18454_;
  wire _18455_;
  wire _18456_;
  wire _18457_;
  wire _18458_;
  wire _18459_;
  wire _18460_;
  wire _18461_;
  wire _18462_;
  wire _18463_;
  wire _18464_;
  wire _18465_;
  wire _18466_;
  wire _18467_;
  wire _18468_;
  wire _18469_;
  wire _18470_;
  wire _18471_;
  wire _18472_;
  wire _18473_;
  wire _18474_;
  wire _18475_;
  wire _18476_;
  wire _18477_;
  wire _18478_;
  wire _18479_;
  wire _18480_;
  wire _18481_;
  wire _18482_;
  wire _18483_;
  wire _18484_;
  wire _18485_;
  wire _18486_;
  wire _18487_;
  wire _18488_;
  wire _18489_;
  wire _18490_;
  wire _18491_;
  wire _18492_;
  wire _18493_;
  wire _18494_;
  wire _18495_;
  wire _18496_;
  wire _18497_;
  wire _18498_;
  wire _18499_;
  wire _18500_;
  wire _18501_;
  wire _18502_;
  wire _18503_;
  wire _18504_;
  wire _18505_;
  wire _18506_;
  wire _18507_;
  wire _18508_;
  wire _18509_;
  wire _18510_;
  wire _18511_;
  wire _18512_;
  wire _18513_;
  wire _18514_;
  wire _18515_;
  wire _18516_;
  wire _18517_;
  wire _18518_;
  wire _18519_;
  wire _18520_;
  wire _18521_;
  wire _18522_;
  wire _18523_;
  wire _18524_;
  wire _18525_;
  wire _18526_;
  wire _18527_;
  wire _18528_;
  wire _18529_;
  wire _18530_;
  wire _18531_;
  wire _18532_;
  wire _18533_;
  wire _18534_;
  wire _18535_;
  wire _18536_;
  wire _18537_;
  wire _18538_;
  wire _18539_;
  wire _18540_;
  wire _18541_;
  wire _18542_;
  wire _18543_;
  wire _18544_;
  wire _18545_;
  wire _18546_;
  wire _18547_;
  wire _18548_;
  wire _18549_;
  wire _18550_;
  wire _18551_;
  wire _18552_;
  wire _18553_;
  wire _18554_;
  wire _18555_;
  wire _18556_;
  wire _18557_;
  wire _18558_;
  wire _18559_;
  wire _18560_;
  wire _18561_;
  wire _18562_;
  wire _18563_;
  wire _18564_;
  wire _18565_;
  wire _18566_;
  wire _18567_;
  wire _18568_;
  wire _18569_;
  wire _18570_;
  wire _18571_;
  wire _18572_;
  wire _18573_;
  wire _18574_;
  wire _18575_;
  wire _18576_;
  wire _18577_;
  wire _18578_;
  wire _18579_;
  wire _18580_;
  wire _18581_;
  wire _18582_;
  wire _18583_;
  wire _18584_;
  wire _18585_;
  wire _18586_;
  wire _18587_;
  wire _18588_;
  wire _18589_;
  wire _18590_;
  wire _18591_;
  wire _18592_;
  wire _18593_;
  wire _18594_;
  wire _18595_;
  wire _18596_;
  wire _18597_;
  wire _18598_;
  wire _18599_;
  wire _18600_;
  wire _18601_;
  wire _18602_;
  wire _18603_;
  wire _18604_;
  wire _18605_;
  wire _18606_;
  wire _18607_;
  wire _18608_;
  wire _18609_;
  wire _18610_;
  wire _18611_;
  wire _18612_;
  wire _18613_;
  wire _18614_;
  wire _18615_;
  wire _18616_;
  wire _18617_;
  wire _18618_;
  wire _18619_;
  wire _18620_;
  wire _18621_;
  wire _18622_;
  wire _18623_;
  wire _18624_;
  wire _18625_;
  wire _18626_;
  wire _18627_;
  wire _18628_;
  wire _18629_;
  wire _18630_;
  wire _18631_;
  wire _18632_;
  wire _18633_;
  wire _18634_;
  wire _18635_;
  wire _18636_;
  wire _18637_;
  wire _18638_;
  wire _18639_;
  wire _18640_;
  wire _18641_;
  wire _18642_;
  wire _18643_;
  wire _18644_;
  wire _18645_;
  wire _18646_;
  wire _18647_;
  wire _18648_;
  wire _18649_;
  wire _18650_;
  wire _18651_;
  wire _18652_;
  wire _18653_;
  wire _18654_;
  wire _18655_;
  wire _18656_;
  wire _18657_;
  wire _18658_;
  wire _18659_;
  wire _18660_;
  wire _18661_;
  wire _18662_;
  wire _18663_;
  wire _18664_;
  wire _18665_;
  wire _18666_;
  wire _18667_;
  wire _18668_;
  wire _18669_;
  wire _18670_;
  wire _18671_;
  wire _18672_;
  wire _18673_;
  wire _18674_;
  wire _18675_;
  wire _18676_;
  wire _18677_;
  wire _18678_;
  wire _18679_;
  wire _18680_;
  wire _18681_;
  wire _18682_;
  wire _18683_;
  wire _18684_;
  wire _18685_;
  wire _18686_;
  wire _18687_;
  wire _18688_;
  wire _18689_;
  wire _18690_;
  wire _18691_;
  wire _18692_;
  wire _18693_;
  wire _18694_;
  wire _18695_;
  wire _18696_;
  wire _18697_;
  wire _18698_;
  wire _18699_;
  wire _18700_;
  wire _18701_;
  wire _18702_;
  wire _18703_;
  wire _18704_;
  wire _18705_;
  wire _18706_;
  wire _18707_;
  wire _18708_;
  wire _18709_;
  wire _18710_;
  wire _18711_;
  wire _18712_;
  wire _18713_;
  wire _18714_;
  wire _18715_;
  wire _18716_;
  wire _18717_;
  wire _18718_;
  wire _18719_;
  wire _18720_;
  wire _18721_;
  wire _18722_;
  wire _18723_;
  wire _18724_;
  wire _18725_;
  wire _18726_;
  wire _18727_;
  wire _18728_;
  wire _18729_;
  wire _18730_;
  wire _18731_;
  wire _18732_;
  wire _18733_;
  wire _18734_;
  wire _18735_;
  wire _18736_;
  wire _18737_;
  wire _18738_;
  wire _18739_;
  wire _18740_;
  wire _18741_;
  wire _18742_;
  wire _18743_;
  wire _18744_;
  wire _18745_;
  wire _18746_;
  wire _18747_;
  wire _18748_;
  wire _18749_;
  wire _18750_;
  wire _18751_;
  wire _18752_;
  wire _18753_;
  wire _18754_;
  wire _18755_;
  wire _18756_;
  wire _18757_;
  wire _18758_;
  wire _18759_;
  wire _18760_;
  wire _18761_;
  wire _18762_;
  wire _18763_;
  wire _18764_;
  wire _18765_;
  wire _18766_;
  wire _18767_;
  wire _18768_;
  wire _18769_;
  wire _18770_;
  wire _18771_;
  wire _18772_;
  wire _18773_;
  wire _18774_;
  wire _18775_;
  wire _18776_;
  wire _18777_;
  wire _18778_;
  wire _18779_;
  wire _18780_;
  wire _18781_;
  wire _18782_;
  wire _18783_;
  wire _18784_;
  wire _18785_;
  wire _18786_;
  wire _18787_;
  wire _18788_;
  wire _18789_;
  wire _18790_;
  wire _18791_;
  wire _18792_;
  wire _18793_;
  wire _18794_;
  wire _18795_;
  wire _18796_;
  wire _18797_;
  wire _18798_;
  wire _18799_;
  wire _18800_;
  wire _18801_;
  wire _18802_;
  wire _18803_;
  wire _18804_;
  wire _18805_;
  wire _18806_;
  wire _18807_;
  wire _18808_;
  wire _18809_;
  wire _18810_;
  wire _18811_;
  wire _18812_;
  wire _18813_;
  wire _18814_;
  wire _18815_;
  wire _18816_;
  wire _18817_;
  wire _18818_;
  wire _18819_;
  wire _18820_;
  wire _18821_;
  wire _18822_;
  wire _18823_;
  wire _18824_;
  wire _18825_;
  wire _18826_;
  wire _18827_;
  wire _18828_;
  wire _18829_;
  wire _18830_;
  wire _18831_;
  wire _18832_;
  wire _18833_;
  wire _18834_;
  wire _18835_;
  wire _18836_;
  wire _18837_;
  wire _18838_;
  wire _18839_;
  wire _18840_;
  wire _18841_;
  wire _18842_;
  wire _18843_;
  wire _18844_;
  wire _18845_;
  wire _18846_;
  wire _18847_;
  wire _18848_;
  wire _18849_;
  wire _18850_;
  wire _18851_;
  wire _18852_;
  wire _18853_;
  wire _18854_;
  wire _18855_;
  wire _18856_;
  wire _18857_;
  wire _18858_;
  wire _18859_;
  wire _18860_;
  wire _18861_;
  wire _18862_;
  wire _18863_;
  wire _18864_;
  wire _18865_;
  wire _18866_;
  wire _18867_;
  wire _18868_;
  wire _18869_;
  wire _18870_;
  wire _18871_;
  wire _18872_;
  wire _18873_;
  wire _18874_;
  wire _18875_;
  wire _18876_;
  wire _18877_;
  wire _18878_;
  wire _18879_;
  wire _18880_;
  wire _18881_;
  wire _18882_;
  wire _18883_;
  wire _18884_;
  wire _18885_;
  wire _18886_;
  wire _18887_;
  wire _18888_;
  wire _18889_;
  wire _18890_;
  wire _18891_;
  wire _18892_;
  wire _18893_;
  wire _18894_;
  wire _18895_;
  wire _18896_;
  wire _18897_;
  wire _18898_;
  wire _18899_;
  wire _18900_;
  wire _18901_;
  wire _18902_;
  wire _18903_;
  wire _18904_;
  wire _18905_;
  wire _18906_;
  wire _18907_;
  wire _18908_;
  wire _18909_;
  wire _18910_;
  wire _18911_;
  wire _18912_;
  wire _18913_;
  wire _18914_;
  wire _18915_;
  wire _18916_;
  wire _18917_;
  wire _18918_;
  wire _18919_;
  wire _18920_;
  wire _18921_;
  wire _18922_;
  wire _18923_;
  wire _18924_;
  wire _18925_;
  wire _18926_;
  wire _18927_;
  wire _18928_;
  wire _18929_;
  wire _18930_;
  wire _18931_;
  wire _18932_;
  wire _18933_;
  wire _18934_;
  wire _18935_;
  wire _18936_;
  wire _18937_;
  wire _18938_;
  wire _18939_;
  wire _18940_;
  wire _18941_;
  wire _18942_;
  wire _18943_;
  wire _18944_;
  wire _18945_;
  wire _18946_;
  wire _18947_;
  wire _18948_;
  wire _18949_;
  wire _18950_;
  wire _18951_;
  wire _18952_;
  wire _18953_;
  wire _18954_;
  wire _18955_;
  wire _18956_;
  wire _18957_;
  wire _18958_;
  wire _18959_;
  wire _18960_;
  wire _18961_;
  wire _18962_;
  wire _18963_;
  wire _18964_;
  wire _18965_;
  wire _18966_;
  wire _18967_;
  wire _18968_;
  wire _18969_;
  wire _18970_;
  wire _18971_;
  wire _18972_;
  wire _18973_;
  wire _18974_;
  wire _18975_;
  wire _18976_;
  wire _18977_;
  wire _18978_;
  wire _18979_;
  wire _18980_;
  wire _18981_;
  wire _18982_;
  wire _18983_;
  wire _18984_;
  wire _18985_;
  wire _18986_;
  wire _18987_;
  wire _18988_;
  wire _18989_;
  wire _18990_;
  wire _18991_;
  wire _18992_;
  wire _18993_;
  wire _18994_;
  wire _18995_;
  wire _18996_;
  wire _18997_;
  wire _18998_;
  wire _18999_;
  wire _19000_;
  wire _19001_;
  wire _19002_;
  wire _19003_;
  wire _19004_;
  wire _19005_;
  wire _19006_;
  wire _19007_;
  wire _19008_;
  wire _19009_;
  wire _19010_;
  wire _19011_;
  wire _19012_;
  wire _19013_;
  wire _19014_;
  wire _19015_;
  wire _19016_;
  wire _19017_;
  wire _19018_;
  wire _19019_;
  wire _19020_;
  wire _19021_;
  wire _19022_;
  wire _19023_;
  wire _19024_;
  wire _19025_;
  wire _19026_;
  wire _19027_;
  wire _19028_;
  wire _19029_;
  wire _19030_;
  wire _19031_;
  wire _19032_;
  wire _19033_;
  wire _19034_;
  wire _19035_;
  wire _19036_;
  wire _19037_;
  wire _19038_;
  wire _19039_;
  wire _19040_;
  wire _19041_;
  wire _19042_;
  wire _19043_;
  wire _19044_;
  wire _19045_;
  wire _19046_;
  wire _19047_;
  wire _19048_;
  wire _19049_;
  wire _19050_;
  wire _19051_;
  wire _19052_;
  wire _19053_;
  wire _19054_;
  wire _19055_;
  wire _19056_;
  wire _19057_;
  wire _19058_;
  wire _19059_;
  wire _19060_;
  wire _19061_;
  wire _19062_;
  wire _19063_;
  wire _19064_;
  wire _19065_;
  wire _19066_;
  wire _19067_;
  wire _19068_;
  wire _19069_;
  wire _19070_;
  wire _19071_;
  wire _19072_;
  wire _19073_;
  wire _19074_;
  wire _19075_;
  wire _19076_;
  wire _19077_;
  wire _19078_;
  wire _19079_;
  wire _19080_;
  wire _19081_;
  wire _19082_;
  wire _19083_;
  wire _19084_;
  wire _19085_;
  wire _19086_;
  wire _19087_;
  wire _19088_;
  wire _19089_;
  wire _19090_;
  wire _19091_;
  wire _19092_;
  wire _19093_;
  wire _19094_;
  wire _19095_;
  wire _19096_;
  wire _19097_;
  wire _19098_;
  wire _19099_;
  wire _19100_;
  wire _19101_;
  wire _19102_;
  wire _19103_;
  wire _19104_;
  wire _19105_;
  wire _19106_;
  wire _19107_;
  wire _19108_;
  wire _19109_;
  wire _19110_;
  wire _19111_;
  wire _19112_;
  wire _19113_;
  wire _19114_;
  wire _19115_;
  wire _19116_;
  wire _19117_;
  wire _19118_;
  wire _19119_;
  wire _19120_;
  wire _19121_;
  wire _19122_;
  wire _19123_;
  wire _19124_;
  wire _19125_;
  wire _19126_;
  wire _19127_;
  wire _19128_;
  wire _19129_;
  wire _19130_;
  wire _19131_;
  wire _19132_;
  wire _19133_;
  wire _19134_;
  wire _19135_;
  wire _19136_;
  wire _19137_;
  wire _19138_;
  wire _19139_;
  wire _19140_;
  wire _19141_;
  wire _19142_;
  wire _19143_;
  wire _19144_;
  wire _19145_;
  wire _19146_;
  wire _19147_;
  wire _19148_;
  wire _19149_;
  wire _19150_;
  wire _19151_;
  wire _19152_;
  wire _19153_;
  wire _19154_;
  wire _19155_;
  wire _19156_;
  wire _19157_;
  wire _19158_;
  wire _19159_;
  wire _19160_;
  wire _19161_;
  wire _19162_;
  wire _19163_;
  wire _19164_;
  wire _19165_;
  wire _19166_;
  wire _19167_;
  wire _19168_;
  wire _19169_;
  wire _19170_;
  wire _19171_;
  wire _19172_;
  wire _19173_;
  wire _19174_;
  wire _19175_;
  wire _19176_;
  wire _19177_;
  wire _19178_;
  wire _19179_;
  wire _19180_;
  wire _19181_;
  wire _19182_;
  wire _19183_;
  wire _19184_;
  wire _19185_;
  wire _19186_;
  wire _19187_;
  wire _19188_;
  wire _19189_;
  wire _19190_;
  wire _19191_;
  wire _19192_;
  wire _19193_;
  wire _19194_;
  wire _19195_;
  wire _19196_;
  wire _19197_;
  wire _19198_;
  wire _19199_;
  wire _19200_;
  wire _19201_;
  wire _19202_;
  wire _19203_;
  wire _19204_;
  wire _19205_;
  wire _19206_;
  wire _19207_;
  wire _19208_;
  wire _19209_;
  wire _19210_;
  wire _19211_;
  wire _19212_;
  wire _19213_;
  wire _19214_;
  wire _19215_;
  wire _19216_;
  wire _19217_;
  wire _19218_;
  wire _19219_;
  wire _19220_;
  wire _19221_;
  wire _19222_;
  wire _19223_;
  wire _19224_;
  wire _19225_;
  wire _19226_;
  wire _19227_;
  wire _19228_;
  wire _19229_;
  wire _19230_;
  wire _19231_;
  wire _19232_;
  wire _19233_;
  wire _19234_;
  wire _19235_;
  wire _19236_;
  wire _19237_;
  wire _19238_;
  wire _19239_;
  wire _19240_;
  wire _19241_;
  wire _19242_;
  wire _19243_;
  wire _19244_;
  wire _19245_;
  wire _19246_;
  wire _19247_;
  wire _19248_;
  wire _19249_;
  wire _19250_;
  wire _19251_;
  wire _19252_;
  wire _19253_;
  wire _19254_;
  wire _19255_;
  wire _19256_;
  wire _19257_;
  wire _19258_;
  wire _19259_;
  wire _19260_;
  wire _19261_;
  wire _19262_;
  wire _19263_;
  wire _19264_;
  wire _19265_;
  wire _19266_;
  wire _19267_;
  wire _19268_;
  wire _19269_;
  wire _19270_;
  wire _19271_;
  wire _19272_;
  wire _19273_;
  wire _19274_;
  wire _19275_;
  wire _19276_;
  wire _19277_;
  wire _19278_;
  wire _19279_;
  wire _19280_;
  wire _19281_;
  wire _19282_;
  wire _19283_;
  wire _19284_;
  wire _19285_;
  wire _19286_;
  wire _19287_;
  wire _19288_;
  wire _19289_;
  wire _19290_;
  wire _19291_;
  wire _19292_;
  wire _19293_;
  wire _19294_;
  wire _19295_;
  wire _19296_;
  wire _19297_;
  wire _19298_;
  wire _19299_;
  wire _19300_;
  wire _19301_;
  wire _19302_;
  wire _19303_;
  wire _19304_;
  wire _19305_;
  wire _19306_;
  wire _19307_;
  wire _19308_;
  wire _19309_;
  wire _19310_;
  wire _19311_;
  wire _19312_;
  wire _19313_;
  wire _19314_;
  wire _19315_;
  wire _19316_;
  wire _19317_;
  wire _19318_;
  wire _19319_;
  wire _19320_;
  wire _19321_;
  wire _19322_;
  wire _19323_;
  wire _19324_;
  wire _19325_;
  wire _19326_;
  wire _19327_;
  wire _19328_;
  wire _19329_;
  wire _19330_;
  wire _19331_;
  wire _19332_;
  wire _19333_;
  wire _19334_;
  wire _19335_;
  wire _19336_;
  wire _19337_;
  wire _19338_;
  wire _19339_;
  wire _19340_;
  wire _19341_;
  wire _19342_;
  wire _19343_;
  wire _19344_;
  wire _19345_;
  wire _19346_;
  wire _19347_;
  wire _19348_;
  wire _19349_;
  wire _19350_;
  wire _19351_;
  wire _19352_;
  wire _19353_;
  wire _19354_;
  wire _19355_;
  wire _19356_;
  wire _19357_;
  wire _19358_;
  wire _19359_;
  wire _19360_;
  wire _19361_;
  wire _19362_;
  wire _19363_;
  wire _19364_;
  wire _19365_;
  wire _19366_;
  wire _19367_;
  wire _19368_;
  wire _19369_;
  wire _19370_;
  wire _19371_;
  wire _19372_;
  wire _19373_;
  wire _19374_;
  wire _19375_;
  wire _19376_;
  wire _19377_;
  wire _19378_;
  wire _19379_;
  wire _19380_;
  wire _19381_;
  wire _19382_;
  wire _19383_;
  wire _19384_;
  wire _19385_;
  wire _19386_;
  wire _19387_;
  wire _19388_;
  wire _19389_;
  wire _19390_;
  wire _19391_;
  wire _19392_;
  wire _19393_;
  wire _19394_;
  wire _19395_;
  wire _19396_;
  wire _19397_;
  wire _19398_;
  wire _19399_;
  wire _19400_;
  wire _19401_;
  wire _19402_;
  wire _19403_;
  wire _19404_;
  wire _19405_;
  wire _19406_;
  wire _19407_;
  wire _19408_;
  wire _19409_;
  wire _19410_;
  wire _19411_;
  wire _19412_;
  wire _19413_;
  wire _19414_;
  wire _19415_;
  wire _19416_;
  wire _19417_;
  wire _19418_;
  wire _19419_;
  wire _19420_;
  wire _19421_;
  wire _19422_;
  wire _19423_;
  wire _19424_;
  wire _19425_;
  wire _19426_;
  wire _19427_;
  wire _19428_;
  wire _19429_;
  wire _19430_;
  wire _19431_;
  wire _19432_;
  wire _19433_;
  wire _19434_;
  wire _19435_;
  wire _19436_;
  wire _19437_;
  wire _19438_;
  wire _19439_;
  wire _19440_;
  wire _19441_;
  wire _19442_;
  wire _19443_;
  wire _19444_;
  wire _19445_;
  wire _19446_;
  wire _19447_;
  wire _19448_;
  wire _19449_;
  wire _19450_;
  wire _19451_;
  wire _19452_;
  wire _19453_;
  wire _19454_;
  wire _19455_;
  wire _19456_;
  wire _19457_;
  wire _19458_;
  wire _19459_;
  wire _19460_;
  wire _19461_;
  wire _19462_;
  wire _19463_;
  wire _19464_;
  wire _19465_;
  wire _19466_;
  wire _19467_;
  wire _19468_;
  wire _19469_;
  wire _19470_;
  wire _19471_;
  wire _19472_;
  wire _19473_;
  wire _19474_;
  wire _19475_;
  wire _19476_;
  wire _19477_;
  wire _19478_;
  wire _19479_;
  wire _19480_;
  wire _19481_;
  wire _19482_;
  wire _19483_;
  wire _19484_;
  wire _19485_;
  wire _19486_;
  wire _19487_;
  wire _19488_;
  wire _19489_;
  wire _19490_;
  wire _19491_;
  wire _19492_;
  wire _19493_;
  wire _19494_;
  wire _19495_;
  wire _19496_;
  wire _19497_;
  wire _19498_;
  wire _19499_;
  wire _19500_;
  wire _19501_;
  wire _19502_;
  wire _19503_;
  wire _19504_;
  wire _19505_;
  wire _19506_;
  wire _19507_;
  wire _19508_;
  wire _19509_;
  wire _19510_;
  wire _19511_;
  wire _19512_;
  wire _19513_;
  wire _19514_;
  wire _19515_;
  wire _19516_;
  wire _19517_;
  wire _19518_;
  wire _19519_;
  wire _19520_;
  wire _19521_;
  wire _19522_;
  wire _19523_;
  wire _19524_;
  wire _19525_;
  wire _19526_;
  wire _19527_;
  wire _19528_;
  wire _19529_;
  wire _19530_;
  wire _19531_;
  wire _19532_;
  wire _19533_;
  wire _19534_;
  wire _19535_;
  wire _19536_;
  wire _19537_;
  wire _19538_;
  wire _19539_;
  wire _19540_;
  wire _19541_;
  wire _19542_;
  wire _19543_;
  wire _19544_;
  wire _19545_;
  wire _19546_;
  wire _19547_;
  wire _19548_;
  wire _19549_;
  wire _19550_;
  wire _19551_;
  wire _19552_;
  wire _19553_;
  wire _19554_;
  wire _19555_;
  wire _19556_;
  wire _19557_;
  wire _19558_;
  wire _19559_;
  wire _19560_;
  wire _19561_;
  wire _19562_;
  wire _19563_;
  wire _19564_;
  wire _19565_;
  wire _19566_;
  wire _19567_;
  wire _19568_;
  wire _19569_;
  wire _19570_;
  wire _19571_;
  wire _19572_;
  wire _19573_;
  wire _19574_;
  wire _19575_;
  wire _19576_;
  wire _19577_;
  wire _19578_;
  wire _19579_;
  wire _19580_;
  wire _19581_;
  wire _19582_;
  wire _19583_;
  wire _19584_;
  wire _19585_;
  wire _19586_;
  wire _19587_;
  wire _19588_;
  wire _19589_;
  wire _19590_;
  wire _19591_;
  wire _19592_;
  wire _19593_;
  wire _19594_;
  wire _19595_;
  wire _19596_;
  wire _19597_;
  wire _19598_;
  wire _19599_;
  wire _19600_;
  wire _19601_;
  wire _19602_;
  wire _19603_;
  wire _19604_;
  wire _19605_;
  wire _19606_;
  wire _19607_;
  wire _19608_;
  wire _19609_;
  wire _19610_;
  wire _19611_;
  wire _19612_;
  wire _19613_;
  wire _19614_;
  wire _19615_;
  wire _19616_;
  wire _19617_;
  wire _19618_;
  wire _19619_;
  wire _19620_;
  wire _19621_;
  wire _19622_;
  wire _19623_;
  wire _19624_;
  wire _19625_;
  wire _19626_;
  wire _19627_;
  wire _19628_;
  wire _19629_;
  wire _19630_;
  wire _19631_;
  wire _19632_;
  wire _19633_;
  wire _19634_;
  wire _19635_;
  wire _19636_;
  wire _19637_;
  wire _19638_;
  wire _19639_;
  wire _19640_;
  wire _19641_;
  wire _19642_;
  wire _19643_;
  wire _19644_;
  wire _19645_;
  wire _19646_;
  wire _19647_;
  wire _19648_;
  wire _19649_;
  wire _19650_;
  wire _19651_;
  wire _19652_;
  wire _19653_;
  wire _19654_;
  wire _19655_;
  wire _19656_;
  wire _19657_;
  wire _19658_;
  wire _19659_;
  wire _19660_;
  wire _19661_;
  wire _19662_;
  wire _19663_;
  wire _19664_;
  wire _19665_;
  wire _19666_;
  wire _19667_;
  wire _19668_;
  wire _19669_;
  wire _19670_;
  wire _19671_;
  wire _19672_;
  wire _19673_;
  wire _19674_;
  wire _19675_;
  wire _19676_;
  wire _19677_;
  wire _19678_;
  wire _19679_;
  wire _19680_;
  wire _19681_;
  wire _19682_;
  wire _19683_;
  wire _19684_;
  wire _19685_;
  wire _19686_;
  wire _19687_;
  wire _19688_;
  wire _19689_;
  wire _19690_;
  wire _19691_;
  wire _19692_;
  wire _19693_;
  wire _19694_;
  wire _19695_;
  wire _19696_;
  wire _19697_;
  wire _19698_;
  wire _19699_;
  wire _19700_;
  wire _19701_;
  wire _19702_;
  wire _19703_;
  wire _19704_;
  wire _19705_;
  wire _19706_;
  wire _19707_;
  wire _19708_;
  wire _19709_;
  wire _19710_;
  wire _19711_;
  wire _19712_;
  wire _19713_;
  wire _19714_;
  wire _19715_;
  wire _19716_;
  wire _19717_;
  wire _19718_;
  wire _19719_;
  wire _19720_;
  wire _19721_;
  wire _19722_;
  wire _19723_;
  wire _19724_;
  wire _19725_;
  wire _19726_;
  wire _19727_;
  wire _19728_;
  wire _19729_;
  wire _19730_;
  wire _19731_;
  wire _19732_;
  wire _19733_;
  wire _19734_;
  wire _19735_;
  wire _19736_;
  wire _19737_;
  wire _19738_;
  wire _19739_;
  wire _19740_;
  wire _19741_;
  wire _19742_;
  wire _19743_;
  wire _19744_;
  wire _19745_;
  wire _19746_;
  wire _19747_;
  wire _19748_;
  wire _19749_;
  wire _19750_;
  wire _19751_;
  wire _19752_;
  wire _19753_;
  wire _19754_;
  wire _19755_;
  wire _19756_;
  wire _19757_;
  wire _19758_;
  wire _19759_;
  wire _19760_;
  wire _19761_;
  wire _19762_;
  wire _19763_;
  wire _19764_;
  wire _19765_;
  wire _19766_;
  wire _19767_;
  wire _19768_;
  wire _19769_;
  wire _19770_;
  wire _19771_;
  wire _19772_;
  wire _19773_;
  wire _19774_;
  wire _19775_;
  wire _19776_;
  wire _19777_;
  wire _19778_;
  wire _19779_;
  wire _19780_;
  wire _19781_;
  wire _19782_;
  wire _19783_;
  wire _19784_;
  wire _19785_;
  wire _19786_;
  wire _19787_;
  wire _19788_;
  wire _19789_;
  wire _19790_;
  wire _19791_;
  wire _19792_;
  wire _19793_;
  wire _19794_;
  wire _19795_;
  wire _19796_;
  wire _19797_;
  wire _19798_;
  wire _19799_;
  wire _19800_;
  wire _19801_;
  wire _19802_;
  wire _19803_;
  wire _19804_;
  wire _19805_;
  wire _19806_;
  wire _19807_;
  wire _19808_;
  wire _19809_;
  wire _19810_;
  wire _19811_;
  wire _19812_;
  wire _19813_;
  wire _19814_;
  wire _19815_;
  wire _19816_;
  wire _19817_;
  wire _19818_;
  wire _19819_;
  wire _19820_;
  wire _19821_;
  wire _19822_;
  wire _19823_;
  wire _19824_;
  wire _19825_;
  wire _19826_;
  wire _19827_;
  wire _19828_;
  wire _19829_;
  wire _19830_;
  wire _19831_;
  wire _19832_;
  wire _19833_;
  wire _19834_;
  wire _19835_;
  wire _19836_;
  wire _19837_;
  wire _19838_;
  wire _19839_;
  wire _19840_;
  wire _19841_;
  wire _19842_;
  wire _19843_;
  wire _19844_;
  wire _19845_;
  wire _19846_;
  wire _19847_;
  wire _19848_;
  wire _19849_;
  wire _19850_;
  wire _19851_;
  wire _19852_;
  wire _19853_;
  wire _19854_;
  wire _19855_;
  wire _19856_;
  wire _19857_;
  wire _19858_;
  wire _19859_;
  wire _19860_;
  wire _19861_;
  wire _19862_;
  wire _19863_;
  wire _19864_;
  wire _19865_;
  wire _19866_;
  wire _19867_;
  wire _19868_;
  wire _19869_;
  wire _19870_;
  wire _19871_;
  wire _19872_;
  wire _19873_;
  wire _19874_;
  wire _19875_;
  wire _19876_;
  wire _19877_;
  wire _19878_;
  wire _19879_;
  wire _19880_;
  wire _19881_;
  wire _19882_;
  wire _19883_;
  wire _19884_;
  wire _19885_;
  wire _19886_;
  wire _19887_;
  wire _19888_;
  wire _19889_;
  wire _19890_;
  wire _19891_;
  wire _19892_;
  wire _19893_;
  wire _19894_;
  wire _19895_;
  wire _19896_;
  wire _19897_;
  wire _19898_;
  wire _19899_;
  wire _19900_;
  wire _19901_;
  wire _19902_;
  wire _19903_;
  wire _19904_;
  wire _19905_;
  wire _19906_;
  wire _19907_;
  wire _19908_;
  wire _19909_;
  wire _19910_;
  wire _19911_;
  wire _19912_;
  wire _19913_;
  wire _19914_;
  wire _19915_;
  wire _19916_;
  wire _19917_;
  wire _19918_;
  wire _19919_;
  wire _19920_;
  wire _19921_;
  wire _19922_;
  wire _19923_;
  wire _19924_;
  wire _19925_;
  wire _19926_;
  wire _19927_;
  wire _19928_;
  wire _19929_;
  wire _19930_;
  wire _19931_;
  wire _19932_;
  wire _19933_;
  wire _19934_;
  wire _19935_;
  wire _19936_;
  wire _19937_;
  wire _19938_;
  wire _19939_;
  wire _19940_;
  wire _19941_;
  wire _19942_;
  wire _19943_;
  wire _19944_;
  wire _19945_;
  wire _19946_;
  wire _19947_;
  wire _19948_;
  wire _19949_;
  wire _19950_;
  wire _19951_;
  wire _19952_;
  wire _19953_;
  wire _19954_;
  wire _19955_;
  wire _19956_;
  wire _19957_;
  wire _19958_;
  wire _19959_;
  wire _19960_;
  wire _19961_;
  wire _19962_;
  wire _19963_;
  wire _19964_;
  wire _19965_;
  wire _19966_;
  wire _19967_;
  wire _19968_;
  wire _19969_;
  wire _19970_;
  wire _19971_;
  wire _19972_;
  wire _19973_;
  wire _19974_;
  wire _19975_;
  wire _19976_;
  wire _19977_;
  wire _19978_;
  wire _19979_;
  wire _19980_;
  wire _19981_;
  wire _19982_;
  wire _19983_;
  wire _19984_;
  wire _19985_;
  wire _19986_;
  wire _19987_;
  wire _19988_;
  wire _19989_;
  wire _19990_;
  wire _19991_;
  wire _19992_;
  wire _19993_;
  wire _19994_;
  wire _19995_;
  wire _19996_;
  wire _19997_;
  wire _19998_;
  wire _19999_;
  wire _20000_;
  wire _20001_;
  wire _20002_;
  wire _20003_;
  wire _20004_;
  wire _20005_;
  wire _20006_;
  wire _20007_;
  wire _20008_;
  wire _20009_;
  wire _20010_;
  wire _20011_;
  wire _20012_;
  wire _20013_;
  wire _20014_;
  wire _20015_;
  wire _20016_;
  wire _20017_;
  wire _20018_;
  wire _20019_;
  wire _20020_;
  wire _20021_;
  wire _20022_;
  wire _20023_;
  wire _20024_;
  wire _20025_;
  wire _20026_;
  wire _20027_;
  wire _20028_;
  wire _20029_;
  wire _20030_;
  wire _20031_;
  wire _20032_;
  wire _20033_;
  wire _20034_;
  wire _20035_;
  wire _20036_;
  wire _20037_;
  wire _20038_;
  wire _20039_;
  wire _20040_;
  wire _20041_;
  wire _20042_;
  wire _20043_;
  wire _20044_;
  wire _20045_;
  wire _20046_;
  wire _20047_;
  wire _20048_;
  wire _20049_;
  wire _20050_;
  wire _20051_;
  wire _20052_;
  wire _20053_;
  wire _20054_;
  wire _20055_;
  wire _20056_;
  wire _20057_;
  wire _20058_;
  wire _20059_;
  wire _20060_;
  wire _20061_;
  wire _20062_;
  wire _20063_;
  wire _20064_;
  wire _20065_;
  wire _20066_;
  wire _20067_;
  wire _20068_;
  wire _20069_;
  wire _20070_;
  wire _20071_;
  wire _20072_;
  wire _20073_;
  wire _20074_;
  wire _20075_;
  wire _20076_;
  wire _20077_;
  wire _20078_;
  wire _20079_;
  wire _20080_;
  wire _20081_;
  wire _20082_;
  wire _20083_;
  wire _20084_;
  wire _20085_;
  wire _20086_;
  wire _20087_;
  wire _20088_;
  wire _20089_;
  wire _20090_;
  wire _20091_;
  wire _20092_;
  wire _20093_;
  wire _20094_;
  wire _20095_;
  wire _20096_;
  wire _20097_;
  wire _20098_;
  wire _20099_;
  wire _20100_;
  wire _20101_;
  wire _20102_;
  wire _20103_;
  wire _20104_;
  wire _20105_;
  wire _20106_;
  wire _20107_;
  wire _20108_;
  wire _20109_;
  wire _20110_;
  wire _20111_;
  wire _20112_;
  wire _20113_;
  wire _20114_;
  wire _20115_;
  wire _20116_;
  wire _20117_;
  wire _20118_;
  wire _20119_;
  wire _20120_;
  wire _20121_;
  wire _20122_;
  wire _20123_;
  wire _20124_;
  wire _20125_;
  wire _20126_;
  wire _20127_;
  wire _20128_;
  wire _20129_;
  wire _20130_;
  wire _20131_;
  wire _20132_;
  wire _20133_;
  wire _20134_;
  wire _20135_;
  wire _20136_;
  wire _20137_;
  wire _20138_;
  wire _20139_;
  wire _20140_;
  wire _20141_;
  wire _20142_;
  wire _20143_;
  wire _20144_;
  wire _20145_;
  wire _20146_;
  wire _20147_;
  wire _20148_;
  wire _20149_;
  wire _20150_;
  wire _20151_;
  wire _20152_;
  wire _20153_;
  wire _20154_;
  wire _20155_;
  wire _20156_;
  wire _20157_;
  wire _20158_;
  wire _20159_;
  wire _20160_;
  wire _20161_;
  wire _20162_;
  wire _20163_;
  wire _20164_;
  wire _20165_;
  wire _20166_;
  wire _20167_;
  wire _20168_;
  wire _20169_;
  wire _20170_;
  wire _20171_;
  wire _20172_;
  wire _20173_;
  wire _20174_;
  wire _20175_;
  wire _20176_;
  wire _20177_;
  wire _20178_;
  wire _20179_;
  wire _20180_;
  wire _20181_;
  wire _20182_;
  wire _20183_;
  wire _20184_;
  wire _20185_;
  wire _20186_;
  wire _20187_;
  wire _20188_;
  wire _20189_;
  wire _20190_;
  wire _20191_;
  wire _20192_;
  wire _20193_;
  wire _20194_;
  wire _20195_;
  wire _20196_;
  wire _20197_;
  wire _20198_;
  wire _20199_;
  wire _20200_;
  wire _20201_;
  wire _20202_;
  wire _20203_;
  wire _20204_;
  wire _20205_;
  wire _20206_;
  wire _20207_;
  wire _20208_;
  wire _20209_;
  wire _20210_;
  wire _20211_;
  wire _20212_;
  wire _20213_;
  wire _20214_;
  wire _20215_;
  wire _20216_;
  wire _20217_;
  wire _20218_;
  wire _20219_;
  wire _20220_;
  wire _20221_;
  wire _20222_;
  wire _20223_;
  wire _20224_;
  wire _20225_;
  wire _20226_;
  wire _20227_;
  wire _20228_;
  wire _20229_;
  wire _20230_;
  wire _20231_;
  wire _20232_;
  wire _20233_;
  wire _20234_;
  wire _20235_;
  wire _20236_;
  wire _20237_;
  wire _20238_;
  wire _20239_;
  wire _20240_;
  wire _20241_;
  wire _20242_;
  wire _20243_;
  wire _20244_;
  wire _20245_;
  wire _20246_;
  wire _20247_;
  wire _20248_;
  wire _20249_;
  wire _20250_;
  wire _20251_;
  wire _20252_;
  wire _20253_;
  wire _20254_;
  wire _20255_;
  wire _20256_;
  wire _20257_;
  wire _20258_;
  wire _20259_;
  wire _20260_;
  wire _20261_;
  wire _20262_;
  wire _20263_;
  wire _20264_;
  wire _20265_;
  wire _20266_;
  wire _20267_;
  wire _20268_;
  wire _20269_;
  wire _20270_;
  wire _20271_;
  wire _20272_;
  wire _20273_;
  wire _20274_;
  wire _20275_;
  wire _20276_;
  wire _20277_;
  wire _20278_;
  wire _20279_;
  wire _20280_;
  wire _20281_;
  wire _20282_;
  wire _20283_;
  wire _20284_;
  wire _20285_;
  wire _20286_;
  wire _20287_;
  wire _20288_;
  wire _20289_;
  wire _20290_;
  wire _20291_;
  wire _20292_;
  wire _20293_;
  wire _20294_;
  wire _20295_;
  wire _20296_;
  wire _20297_;
  wire _20298_;
  wire _20299_;
  wire _20300_;
  wire _20301_;
  wire _20302_;
  wire _20303_;
  wire _20304_;
  wire _20305_;
  wire _20306_;
  wire _20307_;
  wire _20308_;
  wire _20309_;
  wire _20310_;
  wire _20311_;
  wire _20312_;
  wire _20313_;
  wire _20314_;
  wire _20315_;
  wire _20316_;
  wire _20317_;
  wire _20318_;
  wire _20319_;
  wire _20320_;
  wire _20321_;
  wire _20322_;
  wire _20323_;
  wire _20324_;
  wire _20325_;
  wire _20326_;
  wire _20327_;
  wire _20328_;
  wire _20329_;
  wire _20330_;
  wire _20331_;
  wire _20332_;
  wire _20333_;
  wire _20334_;
  wire _20335_;
  wire _20336_;
  wire _20337_;
  wire _20338_;
  wire _20339_;
  wire _20340_;
  wire _20341_;
  wire _20342_;
  wire _20343_;
  wire _20344_;
  wire _20345_;
  wire _20346_;
  wire _20347_;
  wire _20348_;
  wire _20349_;
  wire _20350_;
  wire _20351_;
  wire _20352_;
  wire _20353_;
  wire _20354_;
  wire _20355_;
  wire _20356_;
  wire _20357_;
  wire _20358_;
  wire _20359_;
  wire _20360_;
  wire _20361_;
  wire _20362_;
  wire _20363_;
  wire _20364_;
  wire _20365_;
  wire _20366_;
  wire _20367_;
  wire _20368_;
  wire _20369_;
  wire _20370_;
  wire _20371_;
  wire _20372_;
  wire _20373_;
  wire _20374_;
  wire _20375_;
  wire _20376_;
  wire _20377_;
  wire _20378_;
  wire _20379_;
  wire _20380_;
  wire _20381_;
  wire _20382_;
  wire _20383_;
  wire _20384_;
  wire _20385_;
  wire _20386_;
  wire _20387_;
  wire _20388_;
  wire _20389_;
  wire _20390_;
  wire _20391_;
  wire _20392_;
  wire _20393_;
  wire _20394_;
  wire _20395_;
  wire _20396_;
  wire _20397_;
  wire _20398_;
  wire _20399_;
  wire _20400_;
  wire _20401_;
  wire _20402_;
  wire _20403_;
  wire _20404_;
  wire _20405_;
  wire _20406_;
  wire _20407_;
  wire _20408_;
  wire _20409_;
  wire _20410_;
  wire _20411_;
  wire _20412_;
  wire _20413_;
  wire _20414_;
  wire _20415_;
  wire _20416_;
  wire _20417_;
  wire _20418_;
  wire _20419_;
  wire _20420_;
  wire _20421_;
  wire _20422_;
  wire _20423_;
  wire _20424_;
  wire _20425_;
  wire _20426_;
  wire _20427_;
  wire _20428_;
  wire _20429_;
  wire _20430_;
  wire _20431_;
  wire _20432_;
  wire _20433_;
  wire _20434_;
  wire _20435_;
  wire _20436_;
  wire _20437_;
  wire _20438_;
  wire _20439_;
  wire _20440_;
  wire _20441_;
  wire _20442_;
  wire _20443_;
  wire _20444_;
  wire _20445_;
  wire _20446_;
  wire _20447_;
  wire _20448_;
  wire _20449_;
  wire _20450_;
  wire _20451_;
  wire _20452_;
  wire _20453_;
  wire _20454_;
  wire _20455_;
  wire _20456_;
  wire _20457_;
  wire _20458_;
  wire _20459_;
  wire _20460_;
  wire _20461_;
  wire _20462_;
  wire _20463_;
  wire _20464_;
  wire _20465_;
  wire _20466_;
  wire _20467_;
  wire _20468_;
  wire _20469_;
  wire _20470_;
  wire _20471_;
  wire _20472_;
  wire _20473_;
  wire _20474_;
  wire _20475_;
  wire _20476_;
  wire _20477_;
  wire _20478_;
  wire _20479_;
  wire _20480_;
  wire _20481_;
  wire _20482_;
  wire _20483_;
  wire _20484_;
  wire _20485_;
  wire _20486_;
  wire _20487_;
  wire _20488_;
  wire _20489_;
  wire _20490_;
  wire _20491_;
  wire _20492_;
  wire _20493_;
  wire _20494_;
  wire _20495_;
  wire _20496_;
  wire _20497_;
  wire _20498_;
  wire _20499_;
  wire _20500_;
  wire _20501_;
  wire _20502_;
  wire _20503_;
  wire _20504_;
  wire _20505_;
  wire _20506_;
  wire _20507_;
  wire _20508_;
  wire _20509_;
  wire _20510_;
  wire _20511_;
  wire _20512_;
  wire _20513_;
  wire _20514_;
  wire _20515_;
  wire _20516_;
  wire _20517_;
  wire _20518_;
  wire _20519_;
  wire _20520_;
  wire _20521_;
  wire _20522_;
  wire _20523_;
  wire _20524_;
  wire _20525_;
  wire _20526_;
  wire _20527_;
  wire _20528_;
  wire _20529_;
  wire _20530_;
  wire _20531_;
  wire _20532_;
  wire _20533_;
  wire _20534_;
  wire _20535_;
  wire _20536_;
  wire _20537_;
  wire _20538_;
  wire _20539_;
  wire _20540_;
  wire _20541_;
  wire _20542_;
  wire _20543_;
  wire _20544_;
  wire _20545_;
  wire _20546_;
  wire _20547_;
  wire _20548_;
  wire _20549_;
  wire _20550_;
  wire _20551_;
  wire _20552_;
  wire _20553_;
  wire _20554_;
  wire _20555_;
  wire _20556_;
  wire _20557_;
  wire _20558_;
  wire _20559_;
  wire _20560_;
  wire _20561_;
  wire _20562_;
  wire _20563_;
  wire _20564_;
  wire _20565_;
  wire _20566_;
  wire _20567_;
  wire _20568_;
  wire _20569_;
  wire _20570_;
  wire _20571_;
  wire _20572_;
  wire _20573_;
  wire _20574_;
  wire _20575_;
  wire _20576_;
  wire _20577_;
  wire _20578_;
  wire _20579_;
  wire _20580_;
  wire _20581_;
  wire _20582_;
  wire _20583_;
  wire _20584_;
  wire _20585_;
  wire _20586_;
  wire _20587_;
  wire _20588_;
  wire _20589_;
  wire _20590_;
  wire _20591_;
  wire _20592_;
  wire _20593_;
  wire _20594_;
  wire _20595_;
  wire _20596_;
  wire _20597_;
  wire _20598_;
  wire _20599_;
  wire _20600_;
  wire _20601_;
  wire _20602_;
  wire _20603_;
  wire _20604_;
  wire _20605_;
  wire _20606_;
  wire _20607_;
  wire _20608_;
  wire _20609_;
  wire _20610_;
  wire _20611_;
  wire _20612_;
  wire _20613_;
  wire _20614_;
  wire _20615_;
  wire _20616_;
  wire _20617_;
  wire _20618_;
  wire _20619_;
  wire _20620_;
  wire _20621_;
  wire _20622_;
  wire _20623_;
  wire _20624_;
  wire _20625_;
  wire _20626_;
  wire _20627_;
  wire _20628_;
  wire _20629_;
  wire _20630_;
  wire _20631_;
  wire _20632_;
  wire _20633_;
  wire _20634_;
  wire _20635_;
  wire _20636_;
  wire _20637_;
  wire _20638_;
  wire _20639_;
  wire _20640_;
  wire _20641_;
  wire _20642_;
  wire _20643_;
  wire _20644_;
  wire _20645_;
  wire _20646_;
  wire _20647_;
  wire _20648_;
  wire _20649_;
  wire _20650_;
  wire _20651_;
  wire _20652_;
  wire _20653_;
  wire _20654_;
  wire _20655_;
  wire _20656_;
  wire _20657_;
  wire _20658_;
  wire _20659_;
  wire _20660_;
  wire _20661_;
  wire _20662_;
  wire _20663_;
  wire _20664_;
  wire _20665_;
  wire _20666_;
  wire _20667_;
  wire _20668_;
  wire _20669_;
  wire _20670_;
  wire _20671_;
  wire _20672_;
  wire _20673_;
  wire _20674_;
  wire _20675_;
  wire _20676_;
  wire _20677_;
  wire _20678_;
  wire _20679_;
  wire _20680_;
  wire _20681_;
  wire _20682_;
  wire _20683_;
  wire _20684_;
  wire _20685_;
  wire _20686_;
  wire _20687_;
  wire _20688_;
  wire _20689_;
  wire _20690_;
  wire _20691_;
  wire _20692_;
  wire _20693_;
  wire _20694_;
  wire _20695_;
  wire _20696_;
  wire _20697_;
  wire _20698_;
  wire _20699_;
  wire _20700_;
  wire _20701_;
  wire _20702_;
  wire _20703_;
  wire _20704_;
  wire _20705_;
  wire _20706_;
  wire _20707_;
  wire _20708_;
  wire _20709_;
  wire _20710_;
  wire _20711_;
  wire _20712_;
  wire _20713_;
  wire _20714_;
  wire _20715_;
  wire _20716_;
  wire _20717_;
  wire _20718_;
  wire _20719_;
  wire _20720_;
  wire _20721_;
  wire _20722_;
  wire _20723_;
  wire _20724_;
  wire _20725_;
  wire _20726_;
  wire _20727_;
  wire _20728_;
  wire _20729_;
  wire _20730_;
  wire _20731_;
  wire _20732_;
  wire _20733_;
  wire _20734_;
  wire _20735_;
  wire _20736_;
  wire _20737_;
  wire _20738_;
  wire _20739_;
  wire _20740_;
  wire _20741_;
  wire _20742_;
  wire _20743_;
  wire _20744_;
  wire _20745_;
  wire _20746_;
  wire _20747_;
  wire _20748_;
  wire _20749_;
  wire _20750_;
  wire _20751_;
  wire _20752_;
  wire _20753_;
  wire _20754_;
  wire _20755_;
  wire _20756_;
  wire _20757_;
  wire _20758_;
  wire _20759_;
  wire _20760_;
  wire _20761_;
  wire _20762_;
  wire _20763_;
  wire _20764_;
  wire _20765_;
  wire _20766_;
  wire _20767_;
  wire _20768_;
  wire _20769_;
  wire _20770_;
  wire _20771_;
  wire _20772_;
  wire _20773_;
  wire _20774_;
  wire _20775_;
  wire _20776_;
  wire _20777_;
  wire _20778_;
  wire _20779_;
  wire _20780_;
  wire _20781_;
  wire _20782_;
  wire _20783_;
  wire _20784_;
  wire _20785_;
  wire _20786_;
  wire _20787_;
  wire _20788_;
  wire _20789_;
  wire _20790_;
  wire _20791_;
  wire _20792_;
  wire _20793_;
  wire _20794_;
  wire _20795_;
  wire _20796_;
  wire _20797_;
  wire _20798_;
  wire _20799_;
  wire _20800_;
  wire _20801_;
  wire _20802_;
  wire _20803_;
  wire _20804_;
  wire _20805_;
  wire _20806_;
  wire _20807_;
  wire _20808_;
  wire _20809_;
  wire _20810_;
  wire _20811_;
  wire _20812_;
  wire _20813_;
  wire _20814_;
  wire _20815_;
  wire _20816_;
  wire _20817_;
  wire _20818_;
  wire _20819_;
  wire _20820_;
  wire _20821_;
  wire _20822_;
  wire _20823_;
  wire _20824_;
  wire _20825_;
  wire _20826_;
  wire _20827_;
  wire _20828_;
  wire _20829_;
  wire _20830_;
  wire _20831_;
  wire _20832_;
  wire _20833_;
  wire _20834_;
  wire _20835_;
  wire _20836_;
  wire _20837_;
  wire _20838_;
  wire _20839_;
  wire _20840_;
  wire _20841_;
  wire _20842_;
  wire _20843_;
  wire _20844_;
  wire _20845_;
  wire _20846_;
  wire _20847_;
  wire _20848_;
  wire _20849_;
  wire _20850_;
  wire _20851_;
  wire _20852_;
  wire _20853_;
  wire _20854_;
  wire _20855_;
  wire _20856_;
  wire _20857_;
  wire _20858_;
  wire _20859_;
  wire _20860_;
  wire _20861_;
  wire _20862_;
  wire _20863_;
  wire _20864_;
  wire _20865_;
  wire _20866_;
  wire _20867_;
  wire _20868_;
  wire _20869_;
  wire _20870_;
  wire _20871_;
  wire _20872_;
  wire _20873_;
  wire _20874_;
  wire _20875_;
  wire _20876_;
  wire _20877_;
  wire _20878_;
  wire _20879_;
  wire _20880_;
  wire _20881_;
  wire _20882_;
  wire _20883_;
  wire _20884_;
  wire _20885_;
  wire _20886_;
  wire _20887_;
  wire _20888_;
  wire _20889_;
  wire _20890_;
  wire _20891_;
  wire _20892_;
  wire _20893_;
  wire _20894_;
  wire _20895_;
  wire _20896_;
  wire _20897_;
  wire _20898_;
  wire _20899_;
  wire _20900_;
  wire _20901_;
  wire _20902_;
  wire _20903_;
  wire _20904_;
  wire _20905_;
  wire _20906_;
  wire _20907_;
  wire _20908_;
  wire _20909_;
  wire _20910_;
  wire _20911_;
  wire _20912_;
  wire _20913_;
  wire _20914_;
  wire _20915_;
  wire _20916_;
  wire _20917_;
  wire _20918_;
  wire _20919_;
  wire _20920_;
  wire _20921_;
  wire _20922_;
  wire _20923_;
  wire _20924_;
  wire _20925_;
  wire _20926_;
  wire _20927_;
  wire _20928_;
  wire _20929_;
  wire _20930_;
  wire _20931_;
  wire _20932_;
  wire _20933_;
  wire _20934_;
  wire _20935_;
  wire _20936_;
  wire _20937_;
  wire _20938_;
  wire _20939_;
  wire _20940_;
  wire _20941_;
  wire _20942_;
  wire _20943_;
  wire _20944_;
  wire _20945_;
  wire _20946_;
  wire _20947_;
  wire _20948_;
  wire _20949_;
  wire _20950_;
  wire _20951_;
  wire _20952_;
  wire _20953_;
  wire _20954_;
  wire _20955_;
  wire _20956_;
  wire _20957_;
  wire _20958_;
  wire _20959_;
  wire _20960_;
  wire _20961_;
  wire _20962_;
  wire _20963_;
  wire _20964_;
  wire _20965_;
  wire _20966_;
  wire _20967_;
  wire _20968_;
  wire _20969_;
  wire _20970_;
  wire _20971_;
  wire _20972_;
  wire _20973_;
  wire _20974_;
  wire _20975_;
  wire _20976_;
  wire _20977_;
  wire _20978_;
  wire _20979_;
  wire _20980_;
  wire _20981_;
  wire _20982_;
  wire _20983_;
  wire _20984_;
  wire _20985_;
  wire _20986_;
  wire _20987_;
  wire _20988_;
  wire _20989_;
  wire _20990_;
  wire _20991_;
  wire _20992_;
  wire _20993_;
  wire _20994_;
  wire _20995_;
  wire _20996_;
  wire _20997_;
  wire _20998_;
  wire _20999_;
  wire _21000_;
  wire _21001_;
  wire _21002_;
  wire _21003_;
  wire _21004_;
  wire _21005_;
  wire _21006_;
  wire _21007_;
  wire _21008_;
  wire _21009_;
  wire _21010_;
  wire _21011_;
  wire _21012_;
  wire _21013_;
  wire _21014_;
  wire _21015_;
  wire _21016_;
  wire _21017_;
  wire _21018_;
  wire _21019_;
  wire _21020_;
  wire _21021_;
  wire _21022_;
  wire _21023_;
  wire _21024_;
  wire _21025_;
  wire _21026_;
  wire _21027_;
  wire _21028_;
  wire _21029_;
  wire _21030_;
  wire _21031_;
  wire _21032_;
  wire _21033_;
  wire _21034_;
  wire _21035_;
  wire _21036_;
  wire _21037_;
  wire _21038_;
  wire _21039_;
  wire _21040_;
  wire _21041_;
  wire _21042_;
  wire _21043_;
  wire _21044_;
  wire _21045_;
  wire _21046_;
  wire _21047_;
  wire _21048_;
  wire _21049_;
  wire _21050_;
  wire _21051_;
  wire _21052_;
  wire _21053_;
  wire _21054_;
  wire _21055_;
  wire _21056_;
  wire _21057_;
  wire _21058_;
  wire _21059_;
  wire _21060_;
  wire _21061_;
  wire _21062_;
  wire _21063_;
  wire _21064_;
  wire _21065_;
  wire _21066_;
  wire _21067_;
  wire _21068_;
  wire _21069_;
  wire _21070_;
  wire _21071_;
  wire _21072_;
  wire _21073_;
  wire _21074_;
  wire _21075_;
  wire _21076_;
  wire _21077_;
  wire _21078_;
  wire _21079_;
  wire _21080_;
  wire _21081_;
  wire _21082_;
  wire _21083_;
  wire _21084_;
  wire _21085_;
  wire _21086_;
  wire _21087_;
  wire _21088_;
  wire _21089_;
  wire _21090_;
  wire _21091_;
  wire _21092_;
  wire _21093_;
  wire _21094_;
  wire _21095_;
  wire _21096_;
  wire _21097_;
  wire _21098_;
  wire _21099_;
  wire _21100_;
  wire _21101_;
  wire _21102_;
  wire _21103_;
  wire _21104_;
  wire _21105_;
  wire _21106_;
  wire _21107_;
  wire _21108_;
  wire _21109_;
  wire _21110_;
  wire _21111_;
  wire _21112_;
  wire _21113_;
  wire _21114_;
  wire _21115_;
  wire _21116_;
  wire _21117_;
  wire _21118_;
  wire _21119_;
  wire _21120_;
  wire _21121_;
  wire _21122_;
  wire _21123_;
  wire _21124_;
  wire _21125_;
  wire _21126_;
  wire _21127_;
  wire _21128_;
  wire _21129_;
  wire _21130_;
  wire _21131_;
  wire _21132_;
  wire _21133_;
  wire _21134_;
  wire _21135_;
  wire _21136_;
  wire _21137_;
  wire _21138_;
  wire _21139_;
  wire _21140_;
  wire _21141_;
  wire _21142_;
  wire _21143_;
  wire _21144_;
  wire _21145_;
  wire _21146_;
  wire _21147_;
  wire _21148_;
  wire _21149_;
  wire _21150_;
  wire _21151_;
  wire _21152_;
  wire _21153_;
  wire _21154_;
  wire _21155_;
  wire _21156_;
  wire _21157_;
  wire _21158_;
  wire _21159_;
  wire _21160_;
  wire _21161_;
  wire _21162_;
  wire _21163_;
  wire _21164_;
  wire _21165_;
  wire _21166_;
  wire _21167_;
  wire _21168_;
  wire _21169_;
  wire _21170_;
  wire _21171_;
  wire _21172_;
  wire _21173_;
  wire _21174_;
  wire _21175_;
  wire _21176_;
  wire _21177_;
  wire _21178_;
  wire _21179_;
  wire _21180_;
  wire _21181_;
  wire _21182_;
  wire _21183_;
  wire _21184_;
  wire _21185_;
  wire _21186_;
  wire _21187_;
  wire _21188_;
  wire _21189_;
  wire _21190_;
  wire _21191_;
  wire _21192_;
  wire _21193_;
  wire _21194_;
  wire _21195_;
  wire _21196_;
  wire _21197_;
  wire _21198_;
  wire _21199_;
  wire _21200_;
  wire _21201_;
  wire _21202_;
  wire _21203_;
  wire _21204_;
  wire _21205_;
  wire _21206_;
  wire _21207_;
  wire _21208_;
  wire _21209_;
  wire _21210_;
  wire _21211_;
  wire _21212_;
  wire _21213_;
  wire _21214_;
  wire _21215_;
  wire _21216_;
  wire _21217_;
  wire _21218_;
  wire _21219_;
  wire _21220_;
  wire _21221_;
  wire _21222_;
  wire _21223_;
  wire _21224_;
  wire _21225_;
  wire _21226_;
  wire _21227_;
  wire _21228_;
  wire _21229_;
  wire _21230_;
  wire _21231_;
  wire _21232_;
  wire _21233_;
  wire _21234_;
  wire _21235_;
  wire _21236_;
  wire _21237_;
  wire _21238_;
  wire _21239_;
  wire _21240_;
  wire _21241_;
  wire _21242_;
  wire _21243_;
  wire _21244_;
  wire _21245_;
  wire _21246_;
  wire _21247_;
  wire _21248_;
  wire _21249_;
  wire _21250_;
  wire _21251_;
  wire _21252_;
  wire _21253_;
  wire _21254_;
  wire _21255_;
  wire _21256_;
  wire _21257_;
  wire _21258_;
  wire _21259_;
  wire _21260_;
  wire _21261_;
  wire _21262_;
  wire _21263_;
  wire _21264_;
  wire _21265_;
  wire _21266_;
  wire _21267_;
  wire _21268_;
  wire _21269_;
  wire _21270_;
  wire _21271_;
  wire _21272_;
  wire _21273_;
  wire _21274_;
  wire _21275_;
  wire _21276_;
  wire _21277_;
  wire _21278_;
  wire _21279_;
  wire _21280_;
  wire _21281_;
  wire _21282_;
  wire _21283_;
  wire _21284_;
  wire _21285_;
  wire _21286_;
  wire _21287_;
  wire _21288_;
  wire _21289_;
  wire _21290_;
  wire _21291_;
  wire _21292_;
  wire _21293_;
  wire _21294_;
  wire _21295_;
  wire _21296_;
  wire _21297_;
  wire _21298_;
  wire _21299_;
  wire _21300_;
  wire _21301_;
  wire _21302_;
  wire _21303_;
  wire _21304_;
  wire _21305_;
  wire _21306_;
  wire _21307_;
  wire _21308_;
  wire _21309_;
  wire _21310_;
  wire _21311_;
  wire _21312_;
  wire _21313_;
  wire _21314_;
  wire _21315_;
  wire _21316_;
  wire _21317_;
  wire _21318_;
  wire _21319_;
  wire _21320_;
  wire _21321_;
  wire _21322_;
  wire _21323_;
  wire _21324_;
  wire _21325_;
  wire _21326_;
  wire _21327_;
  wire _21328_;
  wire _21329_;
  wire _21330_;
  wire _21331_;
  wire _21332_;
  wire _21333_;
  wire _21334_;
  wire _21335_;
  wire _21336_;
  wire _21337_;
  wire _21338_;
  wire _21339_;
  wire _21340_;
  wire _21341_;
  wire _21342_;
  wire _21343_;
  wire _21344_;
  wire _21345_;
  wire _21346_;
  wire _21347_;
  wire _21348_;
  wire _21349_;
  wire _21350_;
  wire _21351_;
  wire _21352_;
  wire _21353_;
  wire _21354_;
  wire _21355_;
  wire _21356_;
  wire _21357_;
  wire _21358_;
  wire _21359_;
  wire _21360_;
  wire _21361_;
  wire _21362_;
  wire _21363_;
  wire _21364_;
  wire _21365_;
  wire _21366_;
  wire _21367_;
  wire _21368_;
  wire _21369_;
  wire _21370_;
  wire _21371_;
  wire _21372_;
  wire _21373_;
  wire _21374_;
  wire _21375_;
  wire _21376_;
  wire _21377_;
  wire _21378_;
  wire _21379_;
  wire _21380_;
  wire _21381_;
  wire _21382_;
  wire _21383_;
  wire _21384_;
  wire _21385_;
  wire _21386_;
  wire _21387_;
  wire _21388_;
  wire _21389_;
  wire _21390_;
  wire _21391_;
  wire _21392_;
  wire _21393_;
  wire _21394_;
  wire _21395_;
  wire _21396_;
  wire _21397_;
  wire _21398_;
  wire _21399_;
  wire _21400_;
  wire _21401_;
  wire _21402_;
  wire _21403_;
  wire _21404_;
  wire _21405_;
  wire _21406_;
  wire _21407_;
  wire _21408_;
  wire _21409_;
  wire _21410_;
  wire _21411_;
  wire _21412_;
  wire _21413_;
  wire _21414_;
  wire _21415_;
  wire _21416_;
  wire _21417_;
  wire _21418_;
  wire _21419_;
  wire _21420_;
  wire _21421_;
  wire _21422_;
  wire _21423_;
  wire _21424_;
  wire _21425_;
  wire _21426_;
  wire _21427_;
  wire _21428_;
  wire _21429_;
  wire _21430_;
  wire _21431_;
  wire _21432_;
  wire _21433_;
  wire _21434_;
  wire _21435_;
  wire _21436_;
  wire _21437_;
  wire _21438_;
  wire _21439_;
  wire _21440_;
  wire _21441_;
  wire _21442_;
  wire _21443_;
  wire _21444_;
  wire _21445_;
  wire _21446_;
  wire _21447_;
  wire _21448_;
  wire _21449_;
  wire _21450_;
  wire _21451_;
  wire _21452_;
  wire _21453_;
  wire _21454_;
  wire _21455_;
  wire _21456_;
  wire _21457_;
  wire _21458_;
  wire _21459_;
  wire _21460_;
  wire _21461_;
  wire _21462_;
  wire _21463_;
  wire _21464_;
  wire _21465_;
  wire _21466_;
  wire _21467_;
  wire _21468_;
  wire _21469_;
  wire _21470_;
  wire _21471_;
  wire _21472_;
  wire _21473_;
  wire _21474_;
  wire _21475_;
  wire _21476_;
  wire _21477_;
  wire _21478_;
  wire _21479_;
  wire _21480_;
  wire _21481_;
  wire _21482_;
  wire _21483_;
  wire _21484_;
  wire _21485_;
  wire _21486_;
  wire _21487_;
  wire _21488_;
  wire _21489_;
  wire _21490_;
  wire _21491_;
  wire _21492_;
  wire _21493_;
  wire _21494_;
  wire _21495_;
  wire _21496_;
  wire _21497_;
  wire _21498_;
  wire _21499_;
  wire _21500_;
  wire _21501_;
  wire _21502_;
  wire _21503_;
  wire _21504_;
  wire _21505_;
  wire _21506_;
  wire _21507_;
  wire _21508_;
  wire _21509_;
  wire _21510_;
  wire _21511_;
  wire _21512_;
  wire _21513_;
  wire _21514_;
  wire _21515_;
  wire _21516_;
  wire _21517_;
  wire _21518_;
  wire _21519_;
  wire _21520_;
  wire _21521_;
  wire _21522_;
  wire _21523_;
  wire _21524_;
  wire _21525_;
  wire _21526_;
  wire _21527_;
  wire _21528_;
  wire _21529_;
  wire _21530_;
  wire _21531_;
  wire _21532_;
  wire _21533_;
  wire _21534_;
  wire _21535_;
  wire _21536_;
  wire _21537_;
  wire _21538_;
  wire _21539_;
  wire _21540_;
  wire _21541_;
  wire _21542_;
  wire _21543_;
  wire _21544_;
  wire _21545_;
  wire _21546_;
  wire _21547_;
  wire _21548_;
  wire _21549_;
  wire _21550_;
  wire _21551_;
  wire _21552_;
  wire _21553_;
  wire _21554_;
  wire _21555_;
  wire _21556_;
  wire _21557_;
  wire _21558_;
  wire _21559_;
  wire _21560_;
  wire _21561_;
  wire _21562_;
  wire _21563_;
  wire _21564_;
  wire _21565_;
  wire _21566_;
  wire _21567_;
  wire _21568_;
  wire _21569_;
  wire _21570_;
  wire _21571_;
  wire _21572_;
  wire _21573_;
  wire _21574_;
  wire _21575_;
  wire _21576_;
  wire _21577_;
  wire _21578_;
  wire _21579_;
  wire _21580_;
  wire _21581_;
  wire _21582_;
  wire _21583_;
  wire _21584_;
  wire _21585_;
  wire _21586_;
  wire _21587_;
  wire _21588_;
  wire _21589_;
  wire _21590_;
  wire _21591_;
  wire _21592_;
  wire _21593_;
  wire _21594_;
  wire _21595_;
  wire _21596_;
  wire _21597_;
  wire _21598_;
  wire _21599_;
  wire _21600_;
  wire _21601_;
  wire _21602_;
  wire _21603_;
  wire _21604_;
  wire _21605_;
  wire _21606_;
  wire _21607_;
  wire _21608_;
  wire _21609_;
  wire _21610_;
  wire _21611_;
  wire _21612_;
  wire _21613_;
  wire _21614_;
  wire _21615_;
  wire _21616_;
  wire _21617_;
  wire _21618_;
  wire _21619_;
  wire _21620_;
  wire _21621_;
  wire _21622_;
  wire _21623_;
  wire _21624_;
  wire _21625_;
  wire _21626_;
  wire _21627_;
  wire _21628_;
  wire _21629_;
  wire _21630_;
  wire _21631_;
  wire _21632_;
  wire _21633_;
  wire _21634_;
  wire _21635_;
  wire _21636_;
  wire _21637_;
  wire _21638_;
  wire _21639_;
  wire _21640_;
  wire _21641_;
  wire _21642_;
  wire _21643_;
  wire _21644_;
  wire _21645_;
  wire _21646_;
  wire _21647_;
  wire _21648_;
  wire _21649_;
  wire _21650_;
  wire _21651_;
  wire _21652_;
  wire _21653_;
  wire _21654_;
  wire _21655_;
  wire _21656_;
  wire _21657_;
  wire _21658_;
  wire _21659_;
  wire _21660_;
  wire _21661_;
  wire _21662_;
  wire _21663_;
  wire _21664_;
  wire _21665_;
  wire _21666_;
  wire _21667_;
  wire _21668_;
  wire _21669_;
  wire _21670_;
  wire _21671_;
  wire _21672_;
  wire _21673_;
  wire _21674_;
  wire _21675_;
  wire _21676_;
  wire _21677_;
  wire _21678_;
  wire _21679_;
  wire _21680_;
  wire _21681_;
  wire _21682_;
  wire _21683_;
  wire _21684_;
  wire _21685_;
  wire _21686_;
  wire _21687_;
  wire _21688_;
  wire _21689_;
  wire _21690_;
  wire _21691_;
  wire _21692_;
  wire _21693_;
  wire _21694_;
  wire _21695_;
  wire _21696_;
  wire _21697_;
  wire _21698_;
  wire _21699_;
  wire _21700_;
  wire _21701_;
  wire _21702_;
  wire _21703_;
  wire _21704_;
  wire _21705_;
  wire _21706_;
  wire _21707_;
  wire _21708_;
  wire _21709_;
  wire _21710_;
  wire _21711_;
  wire _21712_;
  wire _21713_;
  wire _21714_;
  wire _21715_;
  wire _21716_;
  wire _21717_;
  wire _21718_;
  wire _21719_;
  wire _21720_;
  wire _21721_;
  wire _21722_;
  wire _21723_;
  wire _21724_;
  wire _21725_;
  wire _21726_;
  wire _21727_;
  wire _21728_;
  wire _21729_;
  wire _21730_;
  wire _21731_;
  wire _21732_;
  wire _21733_;
  wire _21734_;
  wire _21735_;
  wire _21736_;
  wire _21737_;
  wire _21738_;
  wire _21739_;
  wire _21740_;
  wire _21741_;
  wire _21742_;
  wire _21743_;
  wire _21744_;
  wire _21745_;
  wire _21746_;
  wire _21747_;
  wire _21748_;
  wire _21749_;
  wire _21750_;
  wire _21751_;
  wire _21752_;
  wire _21753_;
  wire _21754_;
  wire _21755_;
  wire _21756_;
  wire _21757_;
  wire _21758_;
  wire _21759_;
  wire _21760_;
  wire _21761_;
  wire _21762_;
  wire _21763_;
  wire _21764_;
  wire _21765_;
  wire _21766_;
  wire _21767_;
  wire _21768_;
  wire _21769_;
  wire _21770_;
  wire _21771_;
  wire _21772_;
  wire _21773_;
  wire _21774_;
  wire _21775_;
  wire _21776_;
  wire _21777_;
  wire _21778_;
  wire _21779_;
  wire _21780_;
  wire _21781_;
  wire _21782_;
  wire _21783_;
  wire _21784_;
  wire _21785_;
  wire _21786_;
  wire _21787_;
  wire _21788_;
  wire _21789_;
  wire _21790_;
  wire _21791_;
  wire _21792_;
  wire _21793_;
  wire _21794_;
  wire _21795_;
  wire _21796_;
  wire _21797_;
  wire _21798_;
  wire _21799_;
  wire _21800_;
  wire _21801_;
  wire _21802_;
  wire _21803_;
  wire _21804_;
  wire _21805_;
  wire _21806_;
  wire _21807_;
  wire _21808_;
  wire _21809_;
  wire _21810_;
  wire _21811_;
  wire _21812_;
  wire _21813_;
  wire _21814_;
  wire _21815_;
  wire _21816_;
  wire _21817_;
  wire _21818_;
  wire _21819_;
  wire _21820_;
  wire _21821_;
  wire _21822_;
  wire _21823_;
  wire _21824_;
  wire _21825_;
  wire _21826_;
  wire _21827_;
  wire _21828_;
  wire _21829_;
  wire _21830_;
  wire _21831_;
  wire _21832_;
  wire _21833_;
  wire _21834_;
  wire _21835_;
  wire _21836_;
  wire _21837_;
  wire _21838_;
  wire _21839_;
  wire _21840_;
  wire _21841_;
  wire _21842_;
  wire _21843_;
  wire _21844_;
  wire _21845_;
  wire _21846_;
  wire _21847_;
  wire _21848_;
  wire _21849_;
  wire _21850_;
  wire _21851_;
  wire _21852_;
  wire _21853_;
  wire _21854_;
  wire _21855_;
  wire _21856_;
  wire _21857_;
  wire _21858_;
  wire _21859_;
  wire _21860_;
  wire _21861_;
  wire _21862_;
  wire _21863_;
  wire _21864_;
  wire _21865_;
  wire _21866_;
  wire _21867_;
  wire _21868_;
  wire _21869_;
  wire _21870_;
  wire _21871_;
  wire _21872_;
  wire _21873_;
  wire _21874_;
  wire _21875_;
  wire _21876_;
  wire _21877_;
  wire _21878_;
  wire _21879_;
  wire _21880_;
  wire _21881_;
  wire _21882_;
  wire _21883_;
  wire _21884_;
  wire _21885_;
  wire _21886_;
  wire _21887_;
  wire _21888_;
  wire _21889_;
  wire _21890_;
  wire _21891_;
  wire _21892_;
  wire _21893_;
  wire _21894_;
  wire _21895_;
  wire _21896_;
  wire _21897_;
  wire _21898_;
  wire _21899_;
  wire _21900_;
  wire _21901_;
  wire _21902_;
  wire _21903_;
  wire _21904_;
  wire _21905_;
  wire _21906_;
  wire _21907_;
  wire _21908_;
  wire _21909_;
  wire _21910_;
  wire _21911_;
  wire _21912_;
  wire _21913_;
  wire _21914_;
  wire _21915_;
  wire _21916_;
  wire _21917_;
  wire _21918_;
  wire _21919_;
  wire _21920_;
  wire _21921_;
  wire _21922_;
  wire _21923_;
  wire _21924_;
  wire _21925_;
  wire _21926_;
  wire _21927_;
  wire _21928_;
  wire _21929_;
  wire _21930_;
  wire _21931_;
  wire _21932_;
  wire _21933_;
  wire _21934_;
  wire _21935_;
  wire _21936_;
  wire _21937_;
  wire _21938_;
  wire _21939_;
  wire _21940_;
  wire _21941_;
  wire _21942_;
  wire _21943_;
  wire _21944_;
  wire _21945_;
  wire _21946_;
  wire _21947_;
  wire _21948_;
  wire _21949_;
  wire _21950_;
  wire _21951_;
  wire _21952_;
  wire _21953_;
  wire _21954_;
  wire _21955_;
  wire _21956_;
  wire _21957_;
  wire _21958_;
  wire _21959_;
  wire _21960_;
  wire _21961_;
  wire _21962_;
  wire _21963_;
  wire _21964_;
  wire _21965_;
  wire _21966_;
  wire _21967_;
  wire _21968_;
  wire _21969_;
  wire _21970_;
  wire _21971_;
  wire _21972_;
  wire _21973_;
  wire _21974_;
  wire _21975_;
  wire _21976_;
  wire _21977_;
  wire _21978_;
  wire _21979_;
  wire _21980_;
  wire _21981_;
  wire _21982_;
  wire _21983_;
  wire _21984_;
  wire _21985_;
  wire _21986_;
  wire _21987_;
  wire _21988_;
  wire _21989_;
  wire _21990_;
  wire _21991_;
  wire _21992_;
  wire _21993_;
  wire _21994_;
  wire _21995_;
  wire _21996_;
  wire _21997_;
  wire _21998_;
  wire _21999_;
  wire _22000_;
  wire _22001_;
  wire _22002_;
  wire _22003_;
  wire _22004_;
  wire _22005_;
  wire _22006_;
  wire _22007_;
  wire _22008_;
  wire _22009_;
  wire _22010_;
  wire _22011_;
  wire _22012_;
  wire _22013_;
  wire _22014_;
  wire _22015_;
  wire _22016_;
  wire _22017_;
  wire _22018_;
  wire _22019_;
  wire _22020_;
  wire _22021_;
  wire _22022_;
  wire _22023_;
  wire _22024_;
  wire _22025_;
  wire _22026_;
  wire _22027_;
  wire _22028_;
  wire _22029_;
  wire _22030_;
  wire _22031_;
  wire _22032_;
  wire _22033_;
  wire _22034_;
  wire _22035_;
  wire _22036_;
  wire _22037_;
  wire _22038_;
  wire _22039_;
  wire _22040_;
  wire _22041_;
  wire _22042_;
  wire _22043_;
  wire _22044_;
  wire _22045_;
  wire _22046_;
  wire _22047_;
  wire _22048_;
  wire _22049_;
  wire _22050_;
  wire _22051_;
  wire _22052_;
  wire _22053_;
  wire _22054_;
  wire _22055_;
  wire _22056_;
  wire _22057_;
  wire _22058_;
  wire _22059_;
  wire _22060_;
  wire _22061_;
  wire _22062_;
  wire _22063_;
  wire _22064_;
  wire _22065_;
  wire _22066_;
  wire _22067_;
  wire _22068_;
  wire _22069_;
  wire _22070_;
  wire _22071_;
  wire _22072_;
  wire _22073_;
  wire _22074_;
  wire _22075_;
  wire _22076_;
  wire _22077_;
  wire _22078_;
  wire _22079_;
  wire _22080_;
  wire _22081_;
  wire _22082_;
  wire _22083_;
  wire _22084_;
  wire _22085_;
  wire _22086_;
  wire _22087_;
  wire _22088_;
  wire _22089_;
  wire _22090_;
  wire _22091_;
  wire _22092_;
  wire _22093_;
  wire _22094_;
  wire _22095_;
  wire _22096_;
  wire _22097_;
  wire _22098_;
  wire _22099_;
  wire _22100_;
  wire _22101_;
  wire _22102_;
  wire _22103_;
  wire _22104_;
  wire _22105_;
  wire _22106_;
  wire _22107_;
  wire _22108_;
  wire _22109_;
  wire _22110_;
  wire _22111_;
  wire _22112_;
  wire _22113_;
  wire _22114_;
  wire _22115_;
  wire _22116_;
  wire _22117_;
  wire _22118_;
  wire _22119_;
  wire _22120_;
  wire _22121_;
  wire _22122_;
  wire _22123_;
  wire _22124_;
  wire _22125_;
  wire _22126_;
  wire _22127_;
  wire _22128_;
  wire _22129_;
  wire _22130_;
  wire _22131_;
  wire _22132_;
  wire _22133_;
  wire _22134_;
  wire _22135_;
  wire _22136_;
  wire _22137_;
  wire _22138_;
  wire _22139_;
  wire _22140_;
  wire _22141_;
  wire _22142_;
  wire _22143_;
  wire _22144_;
  wire _22145_;
  wire _22146_;
  wire _22147_;
  wire _22148_;
  wire _22149_;
  wire _22150_;
  wire _22151_;
  wire _22152_;
  wire _22153_;
  wire _22154_;
  wire _22155_;
  wire _22156_;
  wire _22157_;
  wire _22158_;
  wire _22159_;
  wire _22160_;
  wire _22161_;
  wire _22162_;
  wire _22163_;
  wire _22164_;
  wire _22165_;
  wire _22166_;
  wire _22167_;
  wire _22168_;
  wire _22169_;
  wire _22170_;
  wire _22171_;
  wire _22172_;
  wire _22173_;
  wire _22174_;
  wire _22175_;
  wire _22176_;
  wire _22177_;
  wire _22178_;
  wire _22179_;
  wire _22180_;
  wire _22181_;
  wire _22182_;
  wire _22183_;
  wire _22184_;
  wire _22185_;
  wire _22186_;
  wire _22187_;
  wire _22188_;
  wire _22189_;
  wire _22190_;
  wire _22191_;
  wire _22192_;
  wire _22193_;
  wire _22194_;
  wire _22195_;
  wire _22196_;
  wire _22197_;
  wire _22198_;
  wire _22199_;
  wire _22200_;
  wire _22201_;
  wire _22202_;
  wire _22203_;
  wire _22204_;
  wire _22205_;
  wire _22206_;
  wire _22207_;
  wire _22208_;
  wire _22209_;
  wire _22210_;
  wire _22211_;
  wire _22212_;
  wire _22213_;
  wire _22214_;
  wire _22215_;
  wire _22216_;
  wire _22217_;
  wire _22218_;
  wire _22219_;
  wire _22220_;
  wire _22221_;
  wire _22222_;
  wire _22223_;
  wire _22224_;
  wire _22225_;
  wire _22226_;
  wire _22227_;
  wire _22228_;
  wire _22229_;
  wire _22230_;
  wire _22231_;
  wire _22232_;
  wire _22233_;
  wire _22234_;
  wire _22235_;
  wire _22236_;
  wire _22237_;
  wire _22238_;
  wire _22239_;
  wire _22240_;
  wire _22241_;
  wire _22242_;
  wire _22243_;
  wire _22244_;
  wire _22245_;
  wire _22246_;
  wire _22247_;
  wire _22248_;
  wire _22249_;
  wire _22250_;
  wire _22251_;
  wire _22252_;
  wire _22253_;
  wire _22254_;
  wire _22255_;
  wire _22256_;
  wire _22257_;
  wire _22258_;
  wire _22259_;
  wire _22260_;
  wire _22261_;
  wire _22262_;
  wire _22263_;
  wire _22264_;
  wire _22265_;
  wire _22266_;
  wire _22267_;
  wire _22268_;
  wire _22269_;
  wire _22270_;
  wire _22271_;
  wire _22272_;
  wire _22273_;
  wire _22274_;
  wire _22275_;
  wire _22276_;
  wire _22277_;
  wire _22278_;
  wire _22279_;
  wire _22280_;
  wire _22281_;
  wire _22282_;
  wire _22283_;
  wire _22284_;
  wire _22285_;
  wire _22286_;
  wire _22287_;
  wire _22288_;
  wire _22289_;
  wire _22290_;
  wire _22291_;
  wire _22292_;
  wire _22293_;
  wire _22294_;
  wire _22295_;
  wire _22296_;
  wire _22297_;
  wire _22298_;
  wire _22299_;
  wire _22300_;
  wire _22301_;
  wire _22302_;
  wire _22303_;
  wire _22304_;
  wire _22305_;
  wire _22306_;
  wire _22307_;
  wire _22308_;
  wire _22309_;
  wire _22310_;
  wire _22311_;
  wire _22312_;
  wire _22313_;
  wire _22314_;
  wire _22315_;
  wire _22316_;
  wire _22317_;
  wire _22318_;
  wire _22319_;
  wire _22320_;
  wire _22321_;
  wire _22322_;
  wire _22323_;
  wire _22324_;
  wire _22325_;
  wire _22326_;
  wire _22327_;
  wire _22328_;
  wire _22329_;
  wire _22330_;
  wire _22331_;
  wire _22332_;
  wire _22333_;
  wire _22334_;
  wire _22335_;
  wire _22336_;
  wire _22337_;
  wire _22338_;
  wire _22339_;
  wire _22340_;
  wire _22341_;
  wire _22342_;
  wire _22343_;
  wire _22344_;
  wire _22345_;
  wire _22346_;
  wire _22347_;
  wire _22348_;
  wire _22349_;
  wire _22350_;
  wire _22351_;
  wire _22352_;
  wire _22353_;
  wire _22354_;
  wire _22355_;
  wire _22356_;
  wire _22357_;
  wire _22358_;
  wire _22359_;
  wire _22360_;
  wire _22361_;
  wire _22362_;
  wire _22363_;
  wire _22364_;
  wire _22365_;
  wire _22366_;
  wire _22367_;
  wire _22368_;
  wire _22369_;
  wire _22370_;
  wire _22371_;
  wire _22372_;
  wire _22373_;
  wire _22374_;
  wire _22375_;
  wire _22376_;
  wire _22377_;
  wire _22378_;
  wire _22379_;
  wire _22380_;
  wire _22381_;
  wire _22382_;
  wire _22383_;
  wire _22384_;
  wire _22385_;
  wire _22386_;
  wire _22387_;
  wire _22388_;
  wire _22389_;
  wire _22390_;
  wire _22391_;
  wire _22392_;
  wire _22393_;
  wire _22394_;
  wire _22395_;
  wire _22396_;
  wire _22397_;
  wire _22398_;
  wire _22399_;
  wire _22400_;
  wire _22401_;
  wire _22402_;
  wire _22403_;
  wire _22404_;
  wire _22405_;
  wire _22406_;
  wire _22407_;
  wire _22408_;
  wire _22409_;
  wire _22410_;
  wire _22411_;
  wire _22412_;
  wire _22413_;
  wire _22414_;
  wire _22415_;
  wire _22416_;
  wire _22417_;
  wire _22418_;
  wire _22419_;
  wire _22420_;
  wire _22421_;
  wire _22422_;
  wire _22423_;
  wire _22424_;
  wire _22425_;
  wire _22426_;
  wire _22427_;
  wire _22428_;
  wire _22429_;
  wire _22430_;
  wire _22431_;
  wire _22432_;
  wire _22433_;
  wire _22434_;
  wire _22435_;
  wire _22436_;
  wire _22437_;
  wire _22438_;
  wire _22439_;
  wire _22440_;
  wire _22441_;
  wire _22442_;
  wire _22443_;
  wire _22444_;
  wire _22445_;
  wire _22446_;
  wire _22447_;
  wire _22448_;
  wire _22449_;
  wire _22450_;
  wire _22451_;
  wire _22452_;
  wire _22453_;
  wire _22454_;
  wire _22455_;
  wire _22456_;
  wire _22457_;
  wire _22458_;
  wire _22459_;
  wire _22460_;
  wire _22461_;
  wire _22462_;
  wire _22463_;
  wire _22464_;
  wire _22465_;
  wire _22466_;
  wire _22467_;
  wire _22468_;
  wire _22469_;
  wire _22470_;
  wire _22471_;
  wire _22472_;
  wire _22473_;
  wire _22474_;
  wire _22475_;
  wire _22476_;
  wire _22477_;
  wire _22478_;
  wire _22479_;
  wire _22480_;
  wire _22481_;
  wire _22482_;
  wire _22483_;
  wire _22484_;
  wire _22485_;
  wire _22486_;
  wire _22487_;
  wire _22488_;
  wire _22489_;
  wire _22490_;
  wire _22491_;
  wire _22492_;
  wire _22493_;
  wire _22494_;
  wire _22495_;
  wire _22496_;
  wire _22497_;
  wire _22498_;
  wire _22499_;
  wire _22500_;
  wire _22501_;
  wire _22502_;
  wire _22503_;
  wire _22504_;
  wire _22505_;
  wire _22506_;
  wire _22507_;
  wire _22508_;
  wire _22509_;
  wire _22510_;
  wire _22511_;
  wire _22512_;
  wire _22513_;
  wire _22514_;
  wire _22515_;
  wire _22516_;
  wire _22517_;
  wire _22518_;
  wire _22519_;
  wire _22520_;
  wire _22521_;
  wire _22522_;
  wire _22523_;
  wire _22524_;
  wire _22525_;
  wire _22526_;
  wire _22527_;
  wire _22528_;
  wire _22529_;
  wire _22530_;
  wire _22531_;
  wire _22532_;
  wire _22533_;
  wire _22534_;
  wire _22535_;
  wire _22536_;
  wire _22537_;
  wire _22538_;
  wire _22539_;
  wire _22540_;
  wire _22541_;
  wire _22542_;
  wire _22543_;
  wire _22544_;
  wire _22545_;
  wire _22546_;
  wire _22547_;
  wire _22548_;
  wire _22549_;
  wire _22550_;
  wire _22551_;
  wire _22552_;
  wire _22553_;
  wire _22554_;
  wire _22555_;
  wire _22556_;
  wire _22557_;
  wire _22558_;
  wire _22559_;
  wire _22560_;
  wire _22561_;
  wire _22562_;
  wire _22563_;
  wire _22564_;
  wire _22565_;
  wire _22566_;
  wire _22567_;
  wire _22568_;
  wire _22569_;
  wire _22570_;
  wire _22571_;
  wire _22572_;
  wire _22573_;
  wire _22574_;
  wire _22575_;
  wire _22576_;
  wire _22577_;
  wire _22578_;
  wire _22579_;
  wire _22580_;
  wire _22581_;
  wire _22582_;
  wire _22583_;
  wire _22584_;
  wire _22585_;
  wire _22586_;
  wire _22587_;
  wire _22588_;
  wire _22589_;
  wire _22590_;
  wire _22591_;
  wire _22592_;
  wire _22593_;
  wire _22594_;
  wire _22595_;
  wire _22596_;
  wire _22597_;
  wire _22598_;
  wire _22599_;
  wire _22600_;
  wire _22601_;
  wire _22602_;
  wire _22603_;
  wire _22604_;
  wire _22605_;
  wire _22606_;
  wire _22607_;
  wire _22608_;
  wire _22609_;
  wire _22610_;
  wire _22611_;
  wire _22612_;
  wire _22613_;
  wire _22614_;
  wire _22615_;
  wire _22616_;
  wire _22617_;
  wire _22618_;
  wire _22619_;
  wire _22620_;
  wire _22621_;
  wire _22622_;
  wire _22623_;
  wire _22624_;
  wire _22625_;
  wire _22626_;
  wire _22627_;
  wire _22628_;
  wire _22629_;
  wire _22630_;
  wire _22631_;
  wire _22632_;
  wire _22633_;
  wire _22634_;
  wire _22635_;
  wire _22636_;
  wire _22637_;
  wire _22638_;
  wire _22639_;
  wire _22640_;
  wire _22641_;
  wire _22642_;
  wire _22643_;
  wire _22644_;
  wire _22645_;
  wire _22646_;
  wire _22647_;
  wire _22648_;
  wire _22649_;
  wire _22650_;
  wire _22651_;
  wire _22652_;
  wire _22653_;
  wire _22654_;
  wire _22655_;
  wire _22656_;
  wire _22657_;
  wire _22658_;
  wire _22659_;
  wire _22660_;
  wire _22661_;
  wire _22662_;
  wire _22663_;
  wire _22664_;
  wire _22665_;
  wire _22666_;
  wire _22667_;
  wire _22668_;
  wire _22669_;
  wire _22670_;
  wire _22671_;
  wire _22672_;
  wire _22673_;
  wire _22674_;
  wire _22675_;
  wire _22676_;
  wire _22677_;
  wire _22678_;
  wire _22679_;
  wire _22680_;
  wire _22681_;
  wire _22682_;
  wire _22683_;
  wire _22684_;
  wire _22685_;
  wire _22686_;
  wire _22687_;
  wire _22688_;
  wire _22689_;
  wire _22690_;
  wire _22691_;
  wire _22692_;
  wire _22693_;
  wire _22694_;
  wire _22695_;
  wire _22696_;
  wire _22697_;
  wire _22698_;
  wire _22699_;
  wire _22700_;
  wire _22701_;
  wire _22702_;
  wire _22703_;
  wire _22704_;
  wire _22705_;
  wire _22706_;
  wire _22707_;
  wire _22708_;
  wire _22709_;
  wire _22710_;
  wire _22711_;
  wire _22712_;
  wire _22713_;
  wire _22714_;
  wire _22715_;
  wire _22716_;
  wire _22717_;
  wire _22718_;
  wire _22719_;
  wire _22720_;
  wire _22721_;
  wire _22722_;
  wire _22723_;
  wire _22724_;
  wire _22725_;
  wire _22726_;
  wire _22727_;
  wire _22728_;
  wire _22729_;
  wire _22730_;
  wire _22731_;
  wire _22732_;
  wire _22733_;
  wire _22734_;
  wire _22735_;
  wire _22736_;
  wire _22737_;
  wire _22738_;
  wire _22739_;
  wire _22740_;
  wire _22741_;
  wire _22742_;
  wire _22743_;
  wire _22744_;
  wire _22745_;
  wire _22746_;
  wire _22747_;
  wire _22748_;
  wire _22749_;
  wire _22750_;
  wire _22751_;
  wire _22752_;
  wire _22753_;
  wire _22754_;
  wire _22755_;
  wire _22756_;
  wire _22757_;
  wire _22758_;
  wire _22759_;
  wire _22760_;
  wire _22761_;
  wire _22762_;
  wire _22763_;
  wire _22764_;
  wire _22765_;
  wire _22766_;
  wire _22767_;
  wire _22768_;
  wire _22769_;
  wire _22770_;
  wire _22771_;
  wire _22772_;
  wire _22773_;
  wire _22774_;
  wire _22775_;
  wire _22776_;
  wire _22777_;
  wire _22778_;
  wire _22779_;
  wire _22780_;
  wire _22781_;
  wire _22782_;
  wire _22783_;
  wire _22784_;
  wire _22785_;
  wire _22786_;
  wire _22787_;
  wire _22788_;
  wire _22789_;
  wire _22790_;
  wire _22791_;
  wire _22792_;
  wire _22793_;
  wire _22794_;
  wire _22795_;
  wire _22796_;
  wire _22797_;
  wire _22798_;
  wire _22799_;
  wire _22800_;
  wire _22801_;
  wire _22802_;
  wire _22803_;
  wire _22804_;
  wire _22805_;
  wire _22806_;
  wire _22807_;
  wire _22808_;
  wire _22809_;
  wire _22810_;
  wire _22811_;
  wire _22812_;
  wire _22813_;
  wire _22814_;
  wire _22815_;
  wire _22816_;
  wire _22817_;
  wire _22818_;
  wire _22819_;
  wire _22820_;
  wire _22821_;
  wire _22822_;
  wire _22823_;
  wire _22824_;
  wire _22825_;
  wire _22826_;
  wire _22827_;
  wire _22828_;
  wire _22829_;
  wire _22830_;
  wire _22831_;
  wire _22832_;
  wire _22833_;
  wire _22834_;
  wire _22835_;
  wire _22836_;
  wire _22837_;
  wire _22838_;
  wire _22839_;
  wire _22840_;
  wire _22841_;
  wire _22842_;
  wire _22843_;
  wire _22844_;
  wire _22845_;
  wire _22846_;
  wire _22847_;
  wire _22848_;
  wire _22849_;
  wire _22850_;
  wire _22851_;
  wire _22852_;
  wire _22853_;
  wire _22854_;
  wire _22855_;
  wire _22856_;
  wire _22857_;
  wire _22858_;
  wire _22859_;
  wire _22860_;
  wire _22861_;
  wire _22862_;
  wire _22863_;
  wire _22864_;
  wire _22865_;
  wire _22866_;
  wire _22867_;
  wire _22868_;
  wire _22869_;
  wire _22870_;
  wire _22871_;
  wire _22872_;
  wire _22873_;
  wire _22874_;
  wire _22875_;
  wire _22876_;
  wire _22877_;
  wire _22878_;
  wire _22879_;
  wire _22880_;
  wire _22881_;
  wire _22882_;
  wire _22883_;
  wire _22884_;
  wire _22885_;
  wire _22886_;
  wire _22887_;
  wire _22888_;
  wire _22889_;
  wire _22890_;
  wire _22891_;
  wire _22892_;
  wire _22893_;
  wire _22894_;
  wire _22895_;
  wire _22896_;
  wire _22897_;
  wire _22898_;
  wire _22899_;
  wire _22900_;
  wire _22901_;
  wire _22902_;
  wire _22903_;
  wire _22904_;
  wire _22905_;
  wire _22906_;
  wire _22907_;
  wire _22908_;
  wire _22909_;
  wire _22910_;
  wire _22911_;
  wire _22912_;
  wire _22913_;
  wire _22914_;
  wire _22915_;
  wire _22916_;
  wire _22917_;
  wire _22918_;
  wire _22919_;
  wire _22920_;
  wire _22921_;
  wire _22922_;
  wire _22923_;
  wire _22924_;
  wire _22925_;
  wire _22926_;
  wire _22927_;
  wire _22928_;
  wire _22929_;
  wire _22930_;
  wire _22931_;
  wire _22932_;
  wire _22933_;
  wire _22934_;
  wire _22935_;
  wire _22936_;
  wire _22937_;
  wire _22938_;
  wire _22939_;
  wire _22940_;
  wire _22941_;
  wire _22942_;
  wire _22943_;
  wire _22944_;
  wire _22945_;
  wire _22946_;
  wire _22947_;
  wire _22948_;
  wire _22949_;
  wire _22950_;
  wire _22951_;
  wire _22952_;
  wire _22953_;
  wire _22954_;
  wire _22955_;
  wire _22956_;
  wire _22957_;
  wire _22958_;
  wire _22959_;
  wire _22960_;
  wire _22961_;
  wire _22962_;
  wire _22963_;
  wire _22964_;
  wire _22965_;
  wire _22966_;
  wire _22967_;
  wire _22968_;
  wire _22969_;
  wire _22970_;
  wire _22971_;
  wire _22972_;
  wire _22973_;
  wire _22974_;
  wire _22975_;
  wire _22976_;
  wire _22977_;
  wire _22978_;
  wire _22979_;
  wire _22980_;
  wire _22981_;
  wire _22982_;
  wire _22983_;
  wire _22984_;
  wire _22985_;
  wire _22986_;
  wire _22987_;
  wire _22988_;
  wire _22989_;
  wire _22990_;
  wire _22991_;
  wire _22992_;
  wire _22993_;
  wire _22994_;
  wire _22995_;
  wire _22996_;
  wire _22997_;
  wire _22998_;
  wire _22999_;
  wire _23000_;
  wire _23001_;
  wire _23002_;
  wire _23003_;
  wire _23004_;
  wire _23005_;
  wire _23006_;
  wire _23007_;
  wire _23008_;
  wire _23009_;
  wire _23010_;
  wire _23011_;
  wire _23012_;
  wire _23013_;
  wire _23014_;
  wire _23015_;
  wire _23016_;
  wire _23017_;
  wire _23018_;
  wire _23019_;
  wire _23020_;
  wire _23021_;
  wire _23022_;
  wire _23023_;
  wire _23024_;
  wire _23025_;
  wire _23026_;
  wire _23027_;
  wire _23028_;
  wire _23029_;
  wire _23030_;
  wire _23031_;
  wire _23032_;
  wire _23033_;
  wire _23034_;
  wire _23035_;
  wire _23036_;
  wire _23037_;
  wire _23038_;
  wire _23039_;
  wire _23040_;
  wire _23041_;
  wire _23042_;
  wire _23043_;
  wire _23044_;
  wire _23045_;
  wire _23046_;
  wire _23047_;
  wire _23048_;
  wire _23049_;
  wire _23050_;
  wire _23051_;
  wire _23052_;
  wire _23053_;
  wire _23054_;
  wire _23055_;
  wire _23056_;
  wire _23057_;
  wire _23058_;
  wire _23059_;
  wire _23060_;
  wire _23061_;
  wire _23062_;
  wire _23063_;
  wire _23064_;
  wire _23065_;
  wire _23066_;
  wire _23067_;
  wire _23068_;
  wire _23069_;
  wire _23070_;
  wire _23071_;
  wire _23072_;
  wire _23073_;
  wire _23074_;
  wire _23075_;
  wire _23076_;
  wire _23077_;
  wire _23078_;
  wire _23079_;
  wire _23080_;
  wire _23081_;
  wire _23082_;
  wire _23083_;
  wire _23084_;
  wire _23085_;
  wire _23086_;
  wire _23087_;
  wire _23088_;
  wire _23089_;
  wire _23090_;
  wire _23091_;
  wire _23092_;
  wire _23093_;
  wire _23094_;
  wire _23095_;
  wire _23096_;
  wire _23097_;
  wire _23098_;
  wire _23099_;
  wire _23100_;
  wire _23101_;
  wire _23102_;
  wire _23103_;
  wire _23104_;
  wire _23105_;
  wire _23106_;
  wire _23107_;
  wire _23108_;
  wire _23109_;
  wire _23110_;
  wire _23111_;
  wire _23112_;
  wire _23113_;
  wire _23114_;
  wire _23115_;
  wire _23116_;
  wire _23117_;
  wire _23118_;
  wire _23119_;
  wire _23120_;
  wire _23121_;
  wire _23122_;
  wire _23123_;
  wire _23124_;
  wire _23125_;
  wire _23126_;
  wire _23127_;
  wire _23128_;
  wire _23129_;
  wire _23130_;
  wire _23131_;
  wire _23132_;
  wire _23133_;
  wire _23134_;
  wire _23135_;
  wire _23136_;
  wire _23137_;
  wire _23138_;
  wire _23139_;
  wire _23140_;
  wire _23141_;
  wire _23142_;
  wire _23143_;
  wire _23144_;
  wire _23145_;
  wire _23146_;
  wire _23147_;
  wire _23148_;
  wire _23149_;
  wire _23150_;
  wire _23151_;
  wire _23152_;
  wire _23153_;
  wire _23154_;
  wire _23155_;
  wire _23156_;
  wire _23157_;
  wire _23158_;
  wire _23159_;
  wire _23160_;
  wire _23161_;
  wire _23162_;
  wire _23163_;
  wire _23164_;
  wire _23165_;
  wire _23166_;
  wire _23167_;
  wire _23168_;
  wire _23169_;
  wire _23170_;
  wire _23171_;
  wire _23172_;
  wire _23173_;
  wire _23174_;
  wire _23175_;
  wire _23176_;
  wire _23177_;
  wire _23178_;
  wire _23179_;
  wire _23180_;
  wire _23181_;
  wire _23182_;
  wire _23183_;
  wire _23184_;
  wire _23185_;
  wire _23186_;
  wire _23187_;
  wire _23188_;
  wire _23189_;
  wire _23190_;
  wire _23191_;
  wire _23192_;
  wire _23193_;
  wire _23194_;
  wire _23195_;
  wire _23196_;
  wire _23197_;
  wire _23198_;
  wire _23199_;
  wire _23200_;
  wire _23201_;
  wire _23202_;
  wire _23203_;
  wire _23204_;
  wire _23205_;
  wire _23206_;
  wire _23207_;
  wire _23208_;
  wire _23209_;
  wire _23210_;
  wire _23211_;
  wire _23212_;
  wire _23213_;
  wire _23214_;
  wire _23215_;
  wire _23216_;
  wire _23217_;
  wire _23218_;
  wire _23219_;
  wire _23220_;
  wire _23221_;
  wire _23222_;
  wire _23223_;
  wire _23224_;
  wire _23225_;
  wire _23226_;
  wire _23227_;
  wire _23228_;
  wire _23229_;
  wire _23230_;
  wire _23231_;
  wire _23232_;
  wire _23233_;
  wire _23234_;
  wire _23235_;
  wire _23236_;
  wire _23237_;
  wire _23238_;
  wire _23239_;
  wire _23240_;
  wire _23241_;
  wire _23242_;
  wire _23243_;
  wire _23244_;
  wire _23245_;
  wire _23246_;
  wire _23247_;
  wire _23248_;
  wire _23249_;
  wire _23250_;
  wire _23251_;
  wire _23252_;
  wire _23253_;
  wire _23254_;
  wire _23255_;
  wire _23256_;
  wire _23257_;
  wire _23258_;
  wire _23259_;
  wire _23260_;
  wire _23261_;
  wire _23262_;
  wire _23263_;
  wire _23264_;
  wire _23265_;
  wire _23266_;
  wire _23267_;
  wire _23268_;
  wire _23269_;
  wire _23270_;
  wire _23271_;
  wire _23272_;
  wire _23273_;
  wire _23274_;
  wire _23275_;
  wire _23276_;
  wire _23277_;
  wire _23278_;
  wire _23279_;
  wire _23280_;
  wire _23281_;
  wire _23282_;
  wire _23283_;
  wire _23284_;
  wire _23285_;
  wire _23286_;
  wire _23287_;
  wire _23288_;
  wire _23289_;
  wire _23290_;
  wire _23291_;
  wire _23292_;
  wire _23293_;
  wire _23294_;
  wire _23295_;
  wire _23296_;
  wire _23297_;
  wire _23298_;
  wire _23299_;
  wire _23300_;
  wire _23301_;
  wire _23302_;
  wire _23303_;
  wire _23304_;
  wire _23305_;
  wire _23306_;
  wire _23307_;
  wire _23308_;
  wire _23309_;
  wire _23310_;
  wire _23311_;
  wire _23312_;
  wire _23313_;
  wire _23314_;
  wire _23315_;
  wire _23316_;
  wire _23317_;
  wire _23318_;
  wire _23319_;
  wire _23320_;
  wire _23321_;
  wire _23322_;
  wire _23323_;
  wire _23324_;
  wire _23325_;
  wire _23326_;
  wire _23327_;
  wire _23328_;
  wire _23329_;
  wire _23330_;
  wire _23331_;
  wire _23332_;
  wire _23333_;
  wire _23334_;
  wire _23335_;
  wire _23336_;
  wire _23337_;
  wire _23338_;
  wire _23339_;
  wire _23340_;
  wire _23341_;
  wire _23342_;
  wire _23343_;
  wire _23344_;
  wire _23345_;
  wire _23346_;
  wire _23347_;
  wire _23348_;
  wire _23349_;
  wire _23350_;
  wire _23351_;
  wire _23352_;
  wire _23353_;
  wire _23354_;
  wire _23355_;
  wire _23356_;
  wire _23357_;
  wire _23358_;
  wire _23359_;
  wire _23360_;
  wire _23361_;
  wire _23362_;
  wire _23363_;
  wire _23364_;
  wire _23365_;
  wire _23366_;
  wire _23367_;
  wire _23368_;
  wire _23369_;
  wire _23370_;
  wire _23371_;
  wire _23372_;
  wire _23373_;
  wire _23374_;
  wire _23375_;
  wire _23376_;
  wire _23377_;
  wire _23378_;
  wire _23379_;
  wire _23380_;
  wire _23381_;
  wire _23382_;
  wire _23383_;
  wire _23384_;
  wire _23385_;
  wire _23386_;
  wire _23387_;
  wire _23388_;
  wire _23389_;
  wire _23390_;
  wire _23391_;
  wire _23392_;
  wire _23393_;
  wire _23394_;
  wire _23395_;
  wire _23396_;
  wire _23397_;
  wire _23398_;
  wire _23399_;
  wire _23400_;
  wire _23401_;
  wire _23402_;
  wire _23403_;
  wire _23404_;
  wire _23405_;
  wire _23406_;
  wire _23407_;
  wire _23408_;
  wire _23409_;
  wire _23410_;
  wire _23411_;
  wire _23412_;
  wire _23413_;
  wire _23414_;
  wire _23415_;
  wire _23416_;
  wire _23417_;
  wire _23418_;
  wire _23419_;
  wire _23420_;
  wire _23421_;
  wire _23422_;
  wire _23423_;
  wire _23424_;
  wire _23425_;
  wire _23426_;
  wire _23427_;
  wire _23428_;
  wire _23429_;
  wire _23430_;
  wire _23431_;
  wire _23432_;
  wire _23433_;
  wire _23434_;
  wire _23435_;
  wire _23436_;
  wire _23437_;
  wire _23438_;
  wire _23439_;
  wire _23440_;
  wire _23441_;
  wire _23442_;
  wire _23443_;
  wire _23444_;
  wire _23445_;
  wire _23446_;
  wire _23447_;
  wire _23448_;
  wire _23449_;
  wire _23450_;
  wire _23451_;
  wire _23452_;
  wire _23453_;
  wire _23454_;
  wire _23455_;
  wire _23456_;
  wire _23457_;
  wire _23458_;
  wire _23459_;
  wire _23460_;
  wire _23461_;
  wire _23462_;
  wire _23463_;
  wire _23464_;
  wire _23465_;
  wire _23466_;
  wire _23467_;
  wire _23468_;
  wire _23469_;
  wire _23470_;
  wire _23471_;
  wire _23472_;
  wire _23473_;
  wire _23474_;
  wire _23475_;
  wire _23476_;
  wire _23477_;
  wire _23478_;
  wire _23479_;
  wire _23480_;
  wire _23481_;
  wire _23482_;
  wire _23483_;
  wire _23484_;
  wire _23485_;
  wire _23486_;
  wire _23487_;
  wire _23488_;
  wire _23489_;
  wire _23490_;
  wire _23491_;
  wire _23492_;
  wire _23493_;
  wire _23494_;
  wire _23495_;
  wire _23496_;
  wire _23497_;
  wire _23498_;
  wire _23499_;
  wire _23500_;
  wire _23501_;
  wire _23502_;
  wire _23503_;
  wire _23504_;
  wire _23505_;
  wire _23506_;
  wire _23507_;
  wire _23508_;
  wire _23509_;
  wire _23510_;
  wire _23511_;
  wire _23512_;
  wire _23513_;
  wire _23514_;
  wire _23515_;
  wire _23516_;
  wire _23517_;
  wire _23518_;
  wire _23519_;
  wire _23520_;
  wire _23521_;
  wire _23522_;
  wire _23523_;
  wire _23524_;
  wire _23525_;
  wire _23526_;
  wire _23527_;
  wire _23528_;
  wire _23529_;
  wire _23530_;
  wire _23531_;
  wire _23532_;
  wire _23533_;
  wire _23534_;
  wire _23535_;
  wire _23536_;
  wire _23537_;
  wire _23538_;
  wire _23539_;
  wire _23540_;
  wire _23541_;
  wire _23542_;
  wire _23543_;
  wire _23544_;
  wire _23545_;
  wire _23546_;
  wire _23547_;
  wire _23548_;
  wire _23549_;
  wire _23550_;
  wire _23551_;
  wire _23552_;
  wire _23553_;
  wire _23554_;
  wire _23555_;
  wire _23556_;
  wire _23557_;
  wire _23558_;
  wire _23559_;
  wire _23560_;
  wire _23561_;
  wire _23562_;
  wire _23563_;
  wire _23564_;
  wire _23565_;
  wire _23566_;
  wire _23567_;
  wire _23568_;
  wire _23569_;
  wire _23570_;
  wire _23571_;
  wire _23572_;
  wire _23573_;
  wire _23574_;
  wire _23575_;
  wire _23576_;
  wire _23577_;
  wire _23578_;
  wire _23579_;
  wire _23580_;
  wire _23581_;
  wire _23582_;
  wire _23583_;
  wire _23584_;
  wire _23585_;
  wire _23586_;
  wire _23587_;
  wire _23588_;
  wire _23589_;
  wire _23590_;
  wire _23591_;
  wire _23592_;
  wire _23593_;
  wire _23594_;
  wire _23595_;
  wire _23596_;
  wire _23597_;
  wire _23598_;
  wire _23599_;
  wire _23600_;
  wire _23601_;
  wire _23602_;
  wire _23603_;
  wire _23604_;
  wire _23605_;
  wire _23606_;
  wire _23607_;
  wire _23608_;
  wire _23609_;
  wire _23610_;
  wire _23611_;
  wire _23612_;
  wire _23613_;
  wire _23614_;
  wire _23615_;
  wire _23616_;
  wire _23617_;
  wire _23618_;
  wire _23619_;
  wire _23620_;
  wire _23621_;
  wire _23622_;
  wire _23623_;
  wire _23624_;
  wire _23625_;
  wire _23626_;
  wire _23627_;
  wire _23628_;
  wire _23629_;
  wire _23630_;
  wire _23631_;
  wire _23632_;
  wire _23633_;
  wire _23634_;
  wire _23635_;
  wire _23636_;
  wire _23637_;
  wire _23638_;
  wire _23639_;
  wire _23640_;
  wire _23641_;
  wire _23642_;
  wire _23643_;
  wire _23644_;
  wire _23645_;
  wire _23646_;
  wire _23647_;
  wire _23648_;
  wire _23649_;
  wire _23650_;
  wire _23651_;
  wire _23652_;
  wire _23653_;
  wire _23654_;
  wire _23655_;
  wire _23656_;
  wire _23657_;
  wire _23658_;
  wire _23659_;
  wire _23660_;
  wire _23661_;
  wire _23662_;
  wire _23663_;
  wire _23664_;
  wire _23665_;
  wire _23666_;
  wire _23667_;
  wire _23668_;
  wire _23669_;
  wire _23670_;
  wire _23671_;
  wire _23672_;
  wire _23673_;
  wire _23674_;
  wire _23675_;
  wire _23676_;
  wire _23677_;
  wire _23678_;
  wire _23679_;
  wire _23680_;
  wire _23681_;
  wire _23682_;
  wire _23683_;
  wire _23684_;
  wire _23685_;
  wire _23686_;
  wire _23687_;
  wire _23688_;
  wire _23689_;
  wire _23690_;
  wire _23691_;
  wire _23692_;
  wire _23693_;
  wire _23694_;
  wire _23695_;
  wire _23696_;
  wire _23697_;
  wire _23698_;
  wire _23699_;
  wire _23700_;
  wire _23701_;
  wire _23702_;
  wire _23703_;
  wire _23704_;
  wire _23705_;
  wire _23706_;
  wire _23707_;
  wire _23708_;
  wire _23709_;
  wire _23710_;
  wire _23711_;
  wire _23712_;
  wire _23713_;
  wire _23714_;
  wire _23715_;
  wire _23716_;
  wire _23717_;
  wire _23718_;
  wire _23719_;
  wire _23720_;
  wire _23721_;
  wire _23722_;
  wire _23723_;
  wire _23724_;
  wire _23725_;
  wire _23726_;
  wire _23727_;
  wire _23728_;
  wire _23729_;
  wire _23730_;
  wire _23731_;
  wire _23732_;
  wire _23733_;
  wire _23734_;
  wire _23735_;
  wire _23736_;
  wire _23737_;
  wire _23738_;
  wire _23739_;
  wire _23740_;
  wire _23741_;
  wire _23742_;
  wire _23743_;
  wire _23744_;
  wire _23745_;
  wire _23746_;
  wire _23747_;
  wire _23748_;
  wire _23749_;
  wire _23750_;
  wire _23751_;
  wire _23752_;
  wire _23753_;
  wire _23754_;
  wire _23755_;
  wire _23756_;
  wire _23757_;
  wire _23758_;
  wire _23759_;
  wire _23760_;
  wire _23761_;
  wire _23762_;
  wire _23763_;
  wire _23764_;
  wire _23765_;
  wire _23766_;
  wire _23767_;
  wire _23768_;
  wire _23769_;
  wire _23770_;
  wire _23771_;
  wire _23772_;
  wire _23773_;
  wire _23774_;
  wire _23775_;
  wire _23776_;
  wire _23777_;
  wire _23778_;
  wire _23779_;
  wire _23780_;
  wire _23781_;
  wire _23782_;
  wire _23783_;
  wire _23784_;
  wire _23785_;
  wire _23786_;
  wire _23787_;
  wire _23788_;
  wire _23789_;
  wire _23790_;
  wire _23791_;
  wire _23792_;
  wire _23793_;
  wire _23794_;
  wire _23795_;
  wire _23796_;
  wire _23797_;
  wire _23798_;
  wire _23799_;
  wire _23800_;
  wire _23801_;
  wire _23802_;
  wire _23803_;
  wire _23804_;
  wire _23805_;
  wire _23806_;
  wire _23807_;
  wire _23808_;
  wire _23809_;
  wire _23810_;
  wire _23811_;
  wire _23812_;
  wire _23813_;
  wire _23814_;
  wire _23815_;
  wire _23816_;
  wire _23817_;
  wire _23818_;
  wire _23819_;
  wire _23820_;
  wire _23821_;
  wire _23822_;
  wire _23823_;
  wire _23824_;
  wire _23825_;
  wire _23826_;
  wire _23827_;
  wire _23828_;
  wire _23829_;
  wire _23830_;
  wire _23831_;
  wire _23832_;
  wire _23833_;
  wire _23834_;
  wire _23835_;
  wire _23836_;
  wire _23837_;
  wire _23838_;
  wire _23839_;
  wire _23840_;
  wire _23841_;
  wire _23842_;
  wire _23843_;
  wire _23844_;
  wire _23845_;
  wire _23846_;
  wire _23847_;
  wire _23848_;
  wire _23849_;
  wire _23850_;
  wire _23851_;
  wire _23852_;
  wire _23853_;
  wire _23854_;
  wire _23855_;
  wire _23856_;
  wire _23857_;
  wire _23858_;
  wire _23859_;
  wire _23860_;
  wire _23861_;
  wire _23862_;
  wire _23863_;
  wire _23864_;
  wire _23865_;
  wire _23866_;
  wire _23867_;
  wire _23868_;
  wire _23869_;
  wire _23870_;
  wire _23871_;
  wire _23872_;
  wire _23873_;
  wire _23874_;
  wire _23875_;
  wire _23876_;
  wire _23877_;
  wire _23878_;
  wire _23879_;
  wire _23880_;
  wire _23881_;
  wire _23882_;
  wire _23883_;
  wire _23884_;
  wire _23885_;
  wire _23886_;
  wire _23887_;
  wire _23888_;
  wire _23889_;
  wire _23890_;
  wire _23891_;
  wire _23892_;
  wire _23893_;
  wire _23894_;
  wire _23895_;
  wire _23896_;
  wire _23897_;
  wire _23898_;
  wire _23899_;
  wire _23900_;
  wire _23901_;
  wire _23902_;
  wire _23903_;
  wire _23904_;
  wire _23905_;
  wire _23906_;
  wire _23907_;
  wire _23908_;
  wire _23909_;
  wire _23910_;
  wire _23911_;
  wire _23912_;
  wire _23913_;
  wire _23914_;
  wire _23915_;
  wire _23916_;
  wire _23917_;
  wire _23918_;
  wire _23919_;
  wire _23920_;
  wire _23921_;
  wire _23922_;
  wire _23923_;
  wire _23924_;
  wire _23925_;
  wire _23926_;
  wire _23927_;
  wire _23928_;
  wire _23929_;
  wire _23930_;
  wire _23931_;
  wire _23932_;
  wire _23933_;
  wire _23934_;
  wire _23935_;
  wire _23936_;
  wire _23937_;
  wire _23938_;
  wire _23939_;
  wire _23940_;
  wire _23941_;
  wire _23942_;
  wire _23943_;
  wire _23944_;
  wire _23945_;
  wire _23946_;
  wire _23947_;
  wire _23948_;
  wire _23949_;
  wire _23950_;
  wire _23951_;
  wire _23952_;
  wire _23953_;
  wire _23954_;
  wire _23955_;
  wire _23956_;
  wire _23957_;
  wire _23958_;
  wire _23959_;
  wire _23960_;
  wire _23961_;
  wire _23962_;
  wire _23963_;
  wire _23964_;
  wire _23965_;
  wire _23966_;
  wire _23967_;
  wire _23968_;
  wire _23969_;
  wire _23970_;
  wire _23971_;
  wire _23972_;
  wire _23973_;
  wire _23974_;
  wire _23975_;
  wire _23976_;
  wire _23977_;
  wire _23978_;
  wire _23979_;
  wire _23980_;
  wire _23981_;
  wire _23982_;
  wire _23983_;
  wire _23984_;
  wire _23985_;
  wire _23986_;
  wire _23987_;
  wire _23988_;
  wire _23989_;
  wire _23990_;
  wire _23991_;
  wire _23992_;
  wire _23993_;
  wire _23994_;
  wire _23995_;
  wire _23996_;
  wire _23997_;
  wire _23998_;
  wire _23999_;
  wire _24000_;
  wire _24001_;
  wire _24002_;
  wire _24003_;
  wire _24004_;
  wire _24005_;
  wire _24006_;
  wire _24007_;
  wire _24008_;
  wire _24009_;
  wire _24010_;
  wire _24011_;
  wire _24012_;
  wire _24013_;
  wire _24014_;
  wire _24015_;
  wire _24016_;
  wire _24017_;
  wire _24018_;
  wire _24019_;
  wire _24020_;
  wire _24021_;
  wire _24022_;
  wire _24023_;
  wire _24024_;
  wire _24025_;
  wire _24026_;
  wire _24027_;
  wire _24028_;
  wire _24029_;
  wire _24030_;
  wire _24031_;
  wire _24032_;
  wire _24033_;
  wire _24034_;
  wire _24035_;
  wire _24036_;
  wire _24037_;
  wire _24038_;
  wire _24039_;
  wire _24040_;
  wire _24041_;
  wire _24042_;
  wire _24043_;
  wire _24044_;
  wire _24045_;
  wire _24046_;
  wire _24047_;
  wire _24048_;
  wire _24049_;
  wire _24050_;
  wire _24051_;
  wire _24052_;
  wire _24053_;
  wire _24054_;
  wire _24055_;
  wire _24056_;
  wire _24057_;
  wire _24058_;
  wire _24059_;
  wire _24060_;
  wire _24061_;
  wire _24062_;
  wire _24063_;
  wire _24064_;
  wire _24065_;
  wire _24066_;
  wire _24067_;
  wire _24068_;
  wire _24069_;
  wire _24070_;
  wire _24071_;
  wire _24072_;
  wire _24073_;
  wire _24074_;
  wire _24075_;
  wire _24076_;
  wire _24077_;
  wire _24078_;
  wire _24079_;
  wire _24080_;
  wire _24081_;
  wire _24082_;
  wire _24083_;
  wire _24084_;
  wire _24085_;
  wire _24086_;
  wire _24087_;
  wire _24088_;
  wire _24089_;
  wire _24090_;
  wire _24091_;
  wire _24092_;
  wire _24093_;
  wire _24094_;
  wire _24095_;
  wire _24096_;
  wire _24097_;
  wire _24098_;
  wire _24099_;
  wire _24100_;
  wire _24101_;
  wire _24102_;
  wire _24103_;
  wire _24104_;
  wire _24105_;
  wire _24106_;
  wire _24107_;
  wire _24108_;
  wire _24109_;
  wire _24110_;
  wire _24111_;
  wire _24112_;
  wire _24113_;
  wire _24114_;
  wire _24115_;
  wire _24116_;
  wire _24117_;
  wire _24118_;
  wire _24119_;
  wire _24120_;
  wire _24121_;
  wire _24122_;
  wire _24123_;
  wire _24124_;
  wire _24125_;
  wire _24126_;
  wire _24127_;
  wire _24128_;
  wire _24129_;
  wire _24130_;
  wire _24131_;
  wire _24132_;
  wire _24133_;
  wire _24134_;
  wire _24135_;
  wire _24136_;
  wire _24137_;
  wire _24138_;
  wire _24139_;
  wire _24140_;
  wire _24141_;
  wire _24142_;
  wire _24143_;
  wire _24144_;
  wire _24145_;
  wire _24146_;
  wire _24147_;
  wire _24148_;
  wire _24149_;
  wire _24150_;
  wire _24151_;
  wire _24152_;
  wire _24153_;
  wire _24154_;
  wire _24155_;
  wire _24156_;
  wire _24157_;
  wire _24158_;
  wire _24159_;
  wire _24160_;
  wire _24161_;
  wire _24162_;
  wire _24163_;
  wire _24164_;
  wire _24165_;
  wire _24166_;
  wire _24167_;
  wire _24168_;
  wire _24169_;
  wire _24170_;
  wire _24171_;
  wire _24172_;
  wire _24173_;
  wire _24174_;
  wire _24175_;
  wire _24176_;
  wire _24177_;
  wire _24178_;
  wire _24179_;
  wire _24180_;
  wire _24181_;
  wire _24182_;
  wire _24183_;
  wire _24184_;
  wire _24185_;
  wire _24186_;
  wire _24187_;
  wire _24188_;
  wire _24189_;
  wire _24190_;
  wire _24191_;
  wire _24192_;
  wire _24193_;
  wire _24194_;
  wire _24195_;
  wire _24196_;
  wire _24197_;
  wire _24198_;
  wire _24199_;
  wire _24200_;
  wire _24201_;
  wire _24202_;
  wire _24203_;
  wire _24204_;
  wire _24205_;
  wire _24206_;
  wire _24207_;
  wire _24208_;
  wire _24209_;
  wire _24210_;
  wire _24211_;
  wire _24212_;
  wire _24213_;
  wire _24214_;
  wire _24215_;
  wire _24216_;
  wire _24217_;
  wire _24218_;
  wire _24219_;
  wire _24220_;
  wire _24221_;
  wire _24222_;
  wire _24223_;
  wire _24224_;
  wire _24225_;
  wire _24226_;
  wire _24227_;
  wire _24228_;
  wire _24229_;
  wire _24230_;
  wire _24231_;
  wire _24232_;
  wire _24233_;
  wire _24234_;
  wire _24235_;
  wire _24236_;
  wire _24237_;
  wire _24238_;
  wire _24239_;
  wire _24240_;
  wire _24241_;
  wire _24242_;
  wire _24243_;
  wire _24244_;
  wire _24245_;
  wire _24246_;
  wire _24247_;
  wire _24248_;
  wire _24249_;
  wire _24250_;
  wire _24251_;
  wire _24252_;
  wire _24253_;
  wire _24254_;
  wire _24255_;
  wire _24256_;
  wire _24257_;
  wire _24258_;
  wire _24259_;
  wire _24260_;
  wire _24261_;
  wire _24262_;
  wire _24263_;
  wire _24264_;
  wire _24265_;
  wire _24266_;
  wire _24267_;
  wire _24268_;
  wire _24269_;
  wire _24270_;
  wire _24271_;
  wire _24272_;
  wire _24273_;
  wire _24274_;
  wire _24275_;
  wire _24276_;
  wire _24277_;
  wire _24278_;
  wire _24279_;
  wire _24280_;
  wire _24281_;
  wire _24282_;
  wire _24283_;
  wire _24284_;
  wire _24285_;
  wire _24286_;
  wire _24287_;
  wire _24288_;
  wire _24289_;
  wire _24290_;
  wire _24291_;
  wire _24292_;
  wire _24293_;
  wire _24294_;
  wire _24295_;
  wire _24296_;
  wire _24297_;
  wire _24298_;
  wire _24299_;
  wire _24300_;
  wire _24301_;
  wire _24302_;
  wire _24303_;
  wire _24304_;
  wire _24305_;
  wire _24306_;
  wire _24307_;
  wire _24308_;
  wire _24309_;
  wire _24310_;
  wire _24311_;
  wire _24312_;
  wire _24313_;
  wire _24314_;
  wire _24315_;
  wire _24316_;
  wire _24317_;
  wire _24318_;
  wire _24319_;
  wire _24320_;
  wire _24321_;
  wire _24322_;
  wire _24323_;
  wire _24324_;
  wire _24325_;
  wire _24326_;
  wire _24327_;
  wire _24328_;
  wire _24329_;
  wire _24330_;
  wire _24331_;
  wire _24332_;
  wire _24333_;
  wire _24334_;
  wire _24335_;
  wire _24336_;
  wire _24337_;
  wire _24338_;
  wire _24339_;
  wire _24340_;
  wire _24341_;
  wire _24342_;
  wire _24343_;
  wire _24344_;
  wire _24345_;
  wire _24346_;
  wire _24347_;
  wire _24348_;
  wire _24349_;
  wire _24350_;
  wire _24351_;
  wire _24352_;
  wire _24353_;
  wire _24354_;
  wire _24355_;
  wire _24356_;
  wire _24357_;
  wire _24358_;
  wire _24359_;
  wire _24360_;
  wire _24361_;
  wire _24362_;
  wire _24363_;
  wire _24364_;
  wire _24365_;
  wire _24366_;
  wire _24367_;
  wire _24368_;
  wire _24369_;
  wire _24370_;
  wire _24371_;
  wire _24372_;
  wire _24373_;
  wire _24374_;
  wire _24375_;
  wire _24376_;
  wire _24377_;
  wire _24378_;
  wire _24379_;
  wire _24380_;
  wire _24381_;
  wire _24382_;
  wire _24383_;
  wire _24384_;
  wire _24385_;
  wire _24386_;
  wire _24387_;
  wire _24388_;
  wire _24389_;
  wire _24390_;
  wire _24391_;
  wire _24392_;
  wire _24393_;
  wire _24394_;
  wire _24395_;
  wire _24396_;
  wire _24397_;
  wire _24398_;
  wire _24399_;
  wire _24400_;
  wire _24401_;
  wire _24402_;
  wire _24403_;
  wire _24404_;
  wire _24405_;
  wire _24406_;
  wire _24407_;
  wire _24408_;
  wire _24409_;
  wire _24410_;
  wire _24411_;
  wire _24412_;
  wire _24413_;
  wire _24414_;
  wire _24415_;
  wire _24416_;
  wire _24417_;
  wire _24418_;
  wire _24419_;
  wire _24420_;
  wire _24421_;
  wire _24422_;
  wire _24423_;
  wire _24424_;
  wire _24425_;
  wire _24426_;
  wire _24427_;
  wire _24428_;
  wire _24429_;
  wire _24430_;
  wire _24431_;
  wire _24432_;
  wire _24433_;
  wire _24434_;
  wire _24435_;
  wire _24436_;
  wire _24437_;
  wire _24438_;
  wire _24439_;
  wire _24440_;
  wire _24441_;
  wire _24442_;
  wire _24443_;
  wire _24444_;
  wire _24445_;
  wire _24446_;
  wire _24447_;
  wire _24448_;
  wire _24449_;
  wire _24450_;
  wire _24451_;
  wire _24452_;
  wire _24453_;
  wire _24454_;
  wire _24455_;
  wire _24456_;
  wire _24457_;
  wire _24458_;
  wire _24459_;
  wire _24460_;
  wire _24461_;
  wire _24462_;
  wire _24463_;
  wire _24464_;
  wire _24465_;
  wire _24466_;
  wire _24467_;
  wire _24468_;
  wire _24469_;
  wire _24470_;
  wire _24471_;
  wire _24472_;
  wire _24473_;
  wire _24474_;
  wire _24475_;
  wire _24476_;
  wire _24477_;
  wire _24478_;
  wire _24479_;
  wire _24480_;
  wire _24481_;
  wire _24482_;
  wire _24483_;
  wire _24484_;
  wire _24485_;
  wire _24486_;
  wire _24487_;
  wire _24488_;
  wire _24489_;
  wire _24490_;
  wire _24491_;
  wire _24492_;
  wire _24493_;
  wire _24494_;
  wire _24495_;
  wire _24496_;
  wire _24497_;
  wire _24498_;
  wire _24499_;
  wire _24500_;
  wire _24501_;
  wire _24502_;
  wire _24503_;
  wire _24504_;
  wire _24505_;
  wire _24506_;
  wire _24507_;
  wire _24508_;
  wire _24509_;
  wire _24510_;
  wire _24511_;
  wire _24512_;
  wire _24513_;
  wire _24514_;
  wire _24515_;
  wire _24516_;
  wire _24517_;
  wire _24518_;
  wire _24519_;
  wire _24520_;
  wire _24521_;
  wire _24522_;
  wire _24523_;
  wire _24524_;
  wire _24525_;
  wire _24526_;
  wire _24527_;
  wire _24528_;
  wire _24529_;
  wire _24530_;
  wire _24531_;
  wire _24532_;
  wire _24533_;
  wire _24534_;
  wire _24535_;
  wire _24536_;
  wire _24537_;
  wire _24538_;
  wire _24539_;
  wire _24540_;
  wire _24541_;
  wire _24542_;
  wire _24543_;
  wire _24544_;
  wire _24545_;
  wire _24546_;
  wire _24547_;
  wire _24548_;
  wire _24549_;
  wire _24550_;
  wire _24551_;
  wire _24552_;
  wire _24553_;
  wire _24554_;
  wire _24555_;
  wire _24556_;
  wire _24557_;
  wire _24558_;
  wire _24559_;
  wire _24560_;
  wire _24561_;
  wire _24562_;
  wire _24563_;
  wire _24564_;
  wire _24565_;
  wire _24566_;
  wire _24567_;
  wire _24568_;
  wire _24569_;
  wire _24570_;
  wire _24571_;
  wire _24572_;
  wire _24573_;
  wire _24574_;
  wire _24575_;
  wire _24576_;
  wire _24577_;
  wire _24578_;
  wire _24579_;
  wire _24580_;
  wire _24581_;
  wire _24582_;
  wire _24583_;
  wire _24584_;
  wire _24585_;
  wire _24586_;
  wire _24587_;
  wire _24588_;
  wire _24589_;
  wire _24590_;
  wire _24591_;
  wire _24592_;
  wire _24593_;
  wire _24594_;
  wire _24595_;
  wire _24596_;
  wire _24597_;
  wire _24598_;
  wire _24599_;
  wire _24600_;
  wire _24601_;
  wire _24602_;
  wire _24603_;
  wire _24604_;
  wire _24605_;
  wire _24606_;
  wire _24607_;
  wire _24608_;
  wire _24609_;
  wire _24610_;
  wire _24611_;
  wire _24612_;
  wire _24613_;
  wire _24614_;
  wire _24615_;
  wire _24616_;
  wire _24617_;
  wire _24618_;
  wire _24619_;
  wire _24620_;
  wire _24621_;
  wire _24622_;
  wire _24623_;
  wire _24624_;
  wire _24625_;
  wire _24626_;
  wire _24627_;
  wire _24628_;
  wire _24629_;
  wire _24630_;
  wire _24631_;
  wire _24632_;
  wire _24633_;
  wire _24634_;
  wire _24635_;
  wire _24636_;
  wire _24637_;
  wire _24638_;
  wire _24639_;
  wire _24640_;
  wire _24641_;
  wire _24642_;
  wire _24643_;
  wire _24644_;
  wire _24645_;
  wire _24646_;
  wire _24647_;
  wire _24648_;
  wire _24649_;
  wire _24650_;
  wire _24651_;
  wire _24652_;
  wire _24653_;
  wire _24654_;
  wire _24655_;
  wire _24656_;
  wire _24657_;
  wire _24658_;
  wire _24659_;
  wire _24660_;
  wire _24661_;
  wire _24662_;
  wire _24663_;
  wire _24664_;
  wire _24665_;
  wire _24666_;
  wire _24667_;
  wire _24668_;
  wire _24669_;
  wire _24670_;
  wire _24671_;
  wire _24672_;
  wire _24673_;
  wire _24674_;
  wire _24675_;
  wire _24676_;
  wire _24677_;
  wire _24678_;
  wire _24679_;
  wire _24680_;
  wire _24681_;
  wire _24682_;
  wire _24683_;
  wire _24684_;
  wire _24685_;
  wire _24686_;
  wire _24687_;
  wire _24688_;
  wire _24689_;
  wire _24690_;
  wire _24691_;
  wire _24692_;
  wire _24693_;
  wire _24694_;
  wire _24695_;
  wire _24696_;
  wire _24697_;
  wire _24698_;
  wire _24699_;
  wire _24700_;
  wire _24701_;
  wire _24702_;
  wire _24703_;
  wire _24704_;
  wire _24705_;
  wire _24706_;
  wire _24707_;
  wire _24708_;
  wire _24709_;
  wire _24710_;
  wire _24711_;
  wire _24712_;
  wire _24713_;
  wire _24714_;
  wire _24715_;
  wire _24716_;
  wire _24717_;
  wire _24718_;
  wire _24719_;
  wire _24720_;
  wire _24721_;
  wire _24722_;
  wire _24723_;
  wire _24724_;
  wire _24725_;
  wire _24726_;
  wire _24727_;
  wire _24728_;
  wire _24729_;
  wire _24730_;
  wire _24731_;
  wire _24732_;
  wire _24733_;
  wire _24734_;
  wire _24735_;
  wire _24736_;
  wire _24737_;
  wire _24738_;
  wire _24739_;
  wire _24740_;
  wire _24741_;
  wire _24742_;
  wire _24743_;
  wire _24744_;
  wire _24745_;
  wire _24746_;
  wire _24747_;
  wire _24748_;
  wire _24749_;
  wire _24750_;
  wire _24751_;
  wire _24752_;
  wire _24753_;
  wire _24754_;
  wire _24755_;
  wire _24756_;
  wire _24757_;
  wire _24758_;
  wire _24759_;
  wire _24760_;
  wire _24761_;
  wire _24762_;
  wire _24763_;
  wire _24764_;
  wire _24765_;
  wire _24766_;
  wire _24767_;
  wire _24768_;
  wire _24769_;
  wire _24770_;
  wire _24771_;
  wire _24772_;
  wire _24773_;
  wire _24774_;
  wire _24775_;
  wire _24776_;
  wire _24777_;
  wire _24778_;
  wire _24779_;
  wire _24780_;
  wire _24781_;
  wire _24782_;
  wire _24783_;
  wire _24784_;
  wire _24785_;
  wire _24786_;
  wire _24787_;
  wire _24788_;
  wire _24789_;
  wire _24790_;
  wire _24791_;
  wire _24792_;
  wire _24793_;
  wire _24794_;
  wire _24795_;
  wire _24796_;
  wire _24797_;
  wire _24798_;
  wire _24799_;
  wire _24800_;
  wire _24801_;
  wire _24802_;
  wire _24803_;
  wire _24804_;
  wire _24805_;
  wire _24806_;
  wire _24807_;
  wire _24808_;
  wire _24809_;
  wire _24810_;
  wire _24811_;
  wire _24812_;
  wire _24813_;
  wire _24814_;
  wire _24815_;
  wire _24816_;
  wire _24817_;
  wire _24818_;
  wire _24819_;
  wire _24820_;
  wire _24821_;
  wire _24822_;
  wire _24823_;
  wire _24824_;
  wire _24825_;
  wire _24826_;
  wire _24827_;
  wire _24828_;
  wire _24829_;
  wire _24830_;
  wire _24831_;
  wire _24832_;
  wire _24833_;
  wire _24834_;
  wire _24835_;
  wire _24836_;
  wire _24837_;
  wire _24838_;
  wire _24839_;
  wire _24840_;
  wire _24841_;
  wire _24842_;
  wire _24843_;
  wire _24844_;
  wire _24845_;
  wire _24846_;
  wire _24847_;
  wire _24848_;
  wire _24849_;
  wire _24850_;
  wire _24851_;
  wire _24852_;
  wire _24853_;
  wire _24854_;
  wire _24855_;
  wire _24856_;
  wire _24857_;
  wire _24858_;
  wire _24859_;
  wire _24860_;
  wire _24861_;
  wire _24862_;
  wire _24863_;
  wire _24864_;
  wire _24865_;
  wire _24866_;
  wire _24867_;
  wire _24868_;
  wire _24869_;
  wire _24870_;
  wire _24871_;
  wire _24872_;
  wire _24873_;
  wire _24874_;
  wire _24875_;
  wire _24876_;
  wire _24877_;
  wire _24878_;
  wire _24879_;
  wire _24880_;
  wire _24881_;
  wire _24882_;
  wire _24883_;
  wire _24884_;
  wire _24885_;
  wire _24886_;
  wire _24887_;
  wire _24888_;
  wire _24889_;
  wire _24890_;
  wire _24891_;
  wire _24892_;
  wire _24893_;
  wire _24894_;
  wire _24895_;
  wire _24896_;
  wire _24897_;
  wire _24898_;
  wire _24899_;
  wire _24900_;
  wire _24901_;
  wire _24902_;
  wire _24903_;
  wire _24904_;
  wire _24905_;
  wire _24906_;
  wire _24907_;
  wire _24908_;
  wire _24909_;
  wire _24910_;
  wire _24911_;
  wire _24912_;
  wire _24913_;
  wire _24914_;
  wire _24915_;
  wire _24916_;
  wire _24917_;
  wire _24918_;
  wire _24919_;
  wire _24920_;
  wire _24921_;
  wire _24922_;
  wire _24923_;
  wire _24924_;
  wire _24925_;
  wire _24926_;
  wire _24927_;
  wire _24928_;
  wire _24929_;
  wire _24930_;
  wire _24931_;
  wire _24932_;
  wire _24933_;
  wire _24934_;
  wire _24935_;
  wire _24936_;
  wire _24937_;
  wire _24938_;
  wire _24939_;
  wire _24940_;
  wire _24941_;
  wire _24942_;
  wire _24943_;
  wire _24944_;
  wire _24945_;
  wire _24946_;
  wire _24947_;
  wire _24948_;
  wire _24949_;
  wire _24950_;
  wire _24951_;
  wire _24952_;
  wire _24953_;
  wire _24954_;
  wire _24955_;
  wire _24956_;
  wire _24957_;
  wire _24958_;
  wire _24959_;
  wire _24960_;
  wire _24961_;
  wire _24962_;
  wire _24963_;
  wire _24964_;
  wire _24965_;
  wire _24966_;
  wire _24967_;
  wire _24968_;
  wire _24969_;
  wire _24970_;
  wire _24971_;
  wire _24972_;
  wire _24973_;
  wire _24974_;
  wire _24975_;
  wire _24976_;
  wire _24977_;
  wire _24978_;
  wire _24979_;
  wire _24980_;
  wire _24981_;
  wire _24982_;
  wire _24983_;
  wire _24984_;
  wire _24985_;
  wire _24986_;
  wire _24987_;
  wire _24988_;
  wire _24989_;
  wire _24990_;
  wire _24991_;
  wire _24992_;
  wire _24993_;
  wire _24994_;
  wire _24995_;
  wire _24996_;
  wire _24997_;
  wire _24998_;
  wire _24999_;
  wire _25000_;
  wire _25001_;
  wire _25002_;
  wire _25003_;
  wire _25004_;
  wire _25005_;
  wire _25006_;
  wire _25007_;
  wire _25008_;
  wire _25009_;
  wire _25010_;
  wire _25011_;
  wire _25012_;
  wire _25013_;
  wire _25014_;
  wire _25015_;
  wire _25016_;
  wire _25017_;
  wire _25018_;
  wire _25019_;
  wire _25020_;
  wire _25021_;
  wire _25022_;
  wire _25023_;
  wire _25024_;
  wire _25025_;
  wire _25026_;
  wire _25027_;
  wire _25028_;
  wire _25029_;
  wire _25030_;
  wire _25031_;
  wire _25032_;
  wire _25033_;
  wire _25034_;
  wire _25035_;
  wire _25036_;
  wire _25037_;
  wire _25038_;
  wire _25039_;
  wire _25040_;
  wire _25041_;
  wire _25042_;
  wire _25043_;
  wire _25044_;
  wire _25045_;
  wire _25046_;
  wire _25047_;
  wire _25048_;
  wire _25049_;
  wire _25050_;
  wire _25051_;
  wire _25052_;
  wire _25053_;
  wire _25054_;
  wire _25055_;
  wire _25056_;
  wire _25057_;
  wire _25058_;
  wire _25059_;
  wire _25060_;
  wire _25061_;
  wire _25062_;
  wire _25063_;
  wire _25064_;
  wire _25065_;
  wire _25066_;
  wire _25067_;
  wire _25068_;
  wire _25069_;
  wire _25070_;
  wire _25071_;
  wire _25072_;
  wire _25073_;
  wire _25074_;
  wire _25075_;
  wire _25076_;
  wire _25077_;
  wire _25078_;
  wire _25079_;
  wire _25080_;
  wire _25081_;
  wire _25082_;
  wire _25083_;
  wire _25084_;
  wire _25085_;
  wire _25086_;
  wire _25087_;
  wire _25088_;
  wire _25089_;
  wire _25090_;
  wire _25091_;
  wire _25092_;
  wire _25093_;
  wire _25094_;
  wire _25095_;
  wire _25096_;
  wire _25097_;
  wire _25098_;
  wire _25099_;
  wire _25100_;
  wire _25101_;
  wire _25102_;
  wire _25103_;
  wire _25104_;
  wire _25105_;
  wire _25106_;
  wire _25107_;
  wire _25108_;
  wire _25109_;
  wire _25110_;
  wire _25111_;
  wire _25112_;
  wire _25113_;
  wire _25114_;
  wire _25115_;
  wire _25116_;
  wire _25117_;
  wire _25118_;
  wire _25119_;
  wire _25120_;
  wire _25121_;
  wire _25122_;
  wire _25123_;
  wire _25124_;
  wire _25125_;
  wire _25126_;
  wire _25127_;
  wire _25128_;
  wire _25129_;
  wire _25130_;
  wire _25131_;
  wire _25132_;
  wire _25133_;
  wire _25134_;
  wire _25135_;
  wire _25136_;
  wire _25137_;
  wire _25138_;
  wire _25139_;
  wire _25140_;
  wire _25141_;
  wire _25142_;
  wire _25143_;
  wire _25144_;
  wire _25145_;
  wire _25146_;
  wire _25147_;
  wire _25148_;
  wire _25149_;
  wire _25150_;
  wire _25151_;
  wire _25152_;
  wire _25153_;
  wire _25154_;
  wire _25155_;
  wire _25156_;
  wire _25157_;
  wire _25158_;
  wire _25159_;
  wire _25160_;
  wire _25161_;
  wire _25162_;
  wire _25163_;
  wire _25164_;
  wire _25165_;
  wire _25166_;
  wire _25167_;
  wire _25168_;
  wire _25169_;
  wire _25170_;
  wire _25171_;
  wire _25172_;
  wire _25173_;
  wire _25174_;
  wire _25175_;
  wire _25176_;
  wire _25177_;
  wire _25178_;
  wire _25179_;
  wire _25180_;
  wire _25181_;
  wire _25182_;
  wire _25183_;
  wire _25184_;
  wire _25185_;
  wire _25186_;
  wire _25187_;
  wire _25188_;
  wire _25189_;
  wire _25190_;
  wire _25191_;
  wire _25192_;
  wire _25193_;
  wire _25194_;
  wire _25195_;
  wire _25196_;
  wire _25197_;
  wire _25198_;
  wire _25199_;
  wire _25200_;
  wire _25201_;
  wire _25202_;
  wire _25203_;
  wire _25204_;
  wire _25205_;
  wire _25206_;
  wire _25207_;
  wire _25208_;
  wire _25209_;
  wire _25210_;
  wire _25211_;
  wire _25212_;
  wire _25213_;
  wire _25214_;
  wire _25215_;
  wire _25216_;
  wire _25217_;
  wire _25218_;
  wire _25219_;
  wire _25220_;
  wire _25221_;
  wire _25222_;
  wire _25223_;
  wire _25224_;
  wire _25225_;
  wire _25226_;
  wire _25227_;
  wire _25228_;
  wire _25229_;
  wire _25230_;
  wire _25231_;
  wire _25232_;
  wire _25233_;
  wire _25234_;
  wire _25235_;
  wire _25236_;
  wire _25237_;
  wire _25238_;
  wire _25239_;
  wire _25240_;
  wire _25241_;
  wire _25242_;
  wire _25243_;
  wire _25244_;
  wire _25245_;
  wire _25246_;
  wire _25247_;
  wire _25248_;
  wire _25249_;
  wire _25250_;
  wire _25251_;
  wire _25252_;
  wire _25253_;
  wire _25254_;
  wire _25255_;
  wire _25256_;
  wire _25257_;
  wire _25258_;
  wire _25259_;
  wire _25260_;
  wire _25261_;
  wire _25262_;
  wire _25263_;
  wire _25264_;
  wire _25265_;
  wire _25266_;
  wire _25267_;
  wire _25268_;
  wire _25269_;
  wire _25270_;
  wire _25271_;
  wire _25272_;
  wire _25273_;
  wire _25274_;
  wire _25275_;
  wire _25276_;
  wire _25277_;
  wire _25278_;
  wire _25279_;
  wire _25280_;
  wire _25281_;
  wire _25282_;
  wire _25283_;
  wire _25284_;
  wire _25285_;
  wire _25286_;
  wire _25287_;
  wire _25288_;
  wire _25289_;
  wire _25290_;
  wire _25291_;
  wire _25292_;
  wire _25293_;
  wire _25294_;
  wire _25295_;
  wire _25296_;
  wire _25297_;
  wire _25298_;
  wire _25299_;
  wire _25300_;
  wire _25301_;
  wire _25302_;
  wire _25303_;
  wire _25304_;
  wire _25305_;
  wire _25306_;
  wire _25307_;
  wire _25308_;
  wire _25309_;
  wire _25310_;
  wire _25311_;
  wire _25312_;
  wire _25313_;
  wire _25314_;
  wire _25315_;
  wire _25316_;
  wire _25317_;
  wire _25318_;
  wire _25319_;
  wire _25320_;
  wire _25321_;
  wire _25322_;
  wire _25323_;
  wire _25324_;
  wire _25325_;
  wire _25326_;
  wire _25327_;
  wire _25328_;
  wire _25329_;
  wire _25330_;
  wire _25331_;
  wire _25332_;
  wire _25333_;
  wire _25334_;
  wire _25335_;
  wire _25336_;
  wire _25337_;
  wire _25338_;
  wire _25339_;
  wire _25340_;
  wire _25341_;
  wire _25342_;
  wire _25343_;
  wire _25344_;
  wire _25345_;
  wire _25346_;
  wire _25347_;
  wire _25348_;
  wire _25349_;
  wire _25350_;
  wire _25351_;
  wire _25352_;
  wire _25353_;
  wire _25354_;
  wire _25355_;
  wire _25356_;
  wire _25357_;
  wire _25358_;
  wire _25359_;
  wire _25360_;
  wire _25361_;
  wire _25362_;
  wire _25363_;
  wire _25364_;
  wire _25365_;
  wire _25366_;
  wire _25367_;
  wire _25368_;
  wire _25369_;
  wire _25370_;
  wire _25371_;
  wire _25372_;
  wire _25373_;
  wire _25374_;
  wire _25375_;
  wire _25376_;
  wire _25377_;
  wire _25378_;
  wire _25379_;
  wire _25380_;
  wire _25381_;
  wire _25382_;
  wire _25383_;
  wire _25384_;
  wire _25385_;
  wire _25386_;
  wire _25387_;
  wire _25388_;
  wire _25389_;
  wire _25390_;
  wire _25391_;
  wire _25392_;
  wire _25393_;
  wire _25394_;
  wire _25395_;
  wire _25396_;
  wire _25397_;
  wire _25398_;
  wire _25399_;
  wire _25400_;
  wire _25401_;
  wire _25402_;
  wire _25403_;
  wire _25404_;
  wire _25405_;
  wire _25406_;
  wire _25407_;
  wire _25408_;
  wire _25409_;
  wire _25410_;
  wire _25411_;
  wire _25412_;
  wire _25413_;
  wire _25414_;
  wire _25415_;
  wire _25416_;
  wire _25417_;
  wire _25418_;
  wire _25419_;
  wire _25420_;
  wire _25421_;
  wire _25422_;
  wire _25423_;
  wire _25424_;
  wire _25425_;
  wire _25426_;
  wire _25427_;
  wire _25428_;
  wire _25429_;
  wire _25430_;
  wire _25431_;
  wire _25432_;
  wire _25433_;
  wire _25434_;
  wire _25435_;
  wire _25436_;
  wire _25437_;
  wire _25438_;
  wire _25439_;
  wire _25440_;
  wire _25441_;
  wire _25442_;
  wire _25443_;
  wire _25444_;
  wire _25445_;
  wire _25446_;
  wire _25447_;
  wire _25448_;
  wire _25449_;
  wire _25450_;
  wire _25451_;
  wire _25452_;
  wire _25453_;
  wire _25454_;
  wire _25455_;
  wire _25456_;
  wire _25457_;
  wire _25458_;
  wire _25459_;
  wire _25460_;
  wire _25461_;
  wire _25462_;
  wire _25463_;
  wire _25464_;
  wire _25465_;
  wire _25466_;
  wire _25467_;
  wire _25468_;
  wire _25469_;
  wire _25470_;
  wire _25471_;
  wire _25472_;
  wire _25473_;
  wire _25474_;
  wire _25475_;
  wire _25476_;
  wire _25477_;
  wire _25478_;
  wire _25479_;
  wire _25480_;
  wire _25481_;
  wire _25482_;
  wire _25483_;
  wire _25484_;
  wire _25485_;
  wire _25486_;
  wire _25487_;
  wire _25488_;
  wire _25489_;
  wire _25490_;
  wire _25491_;
  wire _25492_;
  wire _25493_;
  wire _25494_;
  wire _25495_;
  wire _25496_;
  wire _25497_;
  wire _25498_;
  wire _25499_;
  wire _25500_;
  wire _25501_;
  wire _25502_;
  wire _25503_;
  wire _25504_;
  wire _25505_;
  wire _25506_;
  wire _25507_;
  wire _25508_;
  wire _25509_;
  wire _25510_;
  wire _25511_;
  wire _25512_;
  wire _25513_;
  wire _25514_;
  wire _25515_;
  wire _25516_;
  wire _25517_;
  wire _25518_;
  wire _25519_;
  wire _25520_;
  wire _25521_;
  wire _25522_;
  wire _25523_;
  wire _25524_;
  wire _25525_;
  wire _25526_;
  wire _25527_;
  wire _25528_;
  wire _25529_;
  wire _25530_;
  wire _25531_;
  wire _25532_;
  wire _25533_;
  wire _25534_;
  wire _25535_;
  wire _25536_;
  wire _25537_;
  wire _25538_;
  wire _25539_;
  wire _25540_;
  wire _25541_;
  wire _25542_;
  wire _25543_;
  wire _25544_;
  wire _25545_;
  wire _25546_;
  wire _25547_;
  wire _25548_;
  wire _25549_;
  wire _25550_;
  wire _25551_;
  wire _25552_;
  wire _25553_;
  wire _25554_;
  wire _25555_;
  wire _25556_;
  wire _25557_;
  wire _25558_;
  wire _25559_;
  wire _25560_;
  wire _25561_;
  wire _25562_;
  wire _25563_;
  wire _25564_;
  wire _25565_;
  wire _25566_;
  wire _25567_;
  wire _25568_;
  wire _25569_;
  wire _25570_;
  wire _25571_;
  wire _25572_;
  wire _25573_;
  wire _25574_;
  wire _25575_;
  wire _25576_;
  wire _25577_;
  wire _25578_;
  wire _25579_;
  wire _25580_;
  wire _25581_;
  wire _25582_;
  wire _25583_;
  wire _25584_;
  wire _25585_;
  wire _25586_;
  wire _25587_;
  wire _25588_;
  wire _25589_;
  wire _25590_;
  wire _25591_;
  wire _25592_;
  wire _25593_;
  wire _25594_;
  wire _25595_;
  wire _25596_;
  wire _25597_;
  wire _25598_;
  wire _25599_;
  wire _25600_;
  wire _25601_;
  wire _25602_;
  wire _25603_;
  wire _25604_;
  wire _25605_;
  wire _25606_;
  wire _25607_;
  wire _25608_;
  wire _25609_;
  wire _25610_;
  wire _25611_;
  wire _25612_;
  wire _25613_;
  wire _25614_;
  wire _25615_;
  wire _25616_;
  wire _25617_;
  wire _25618_;
  wire _25619_;
  wire _25620_;
  wire _25621_;
  wire _25622_;
  wire _25623_;
  wire _25624_;
  wire _25625_;
  wire _25626_;
  wire _25627_;
  wire _25628_;
  wire _25629_;
  wire _25630_;
  wire _25631_;
  wire _25632_;
  wire _25633_;
  wire _25634_;
  wire _25635_;
  wire _25636_;
  wire _25637_;
  wire _25638_;
  wire _25639_;
  wire _25640_;
  wire _25641_;
  wire _25642_;
  wire _25643_;
  wire _25644_;
  wire _25645_;
  wire _25646_;
  wire _25647_;
  wire _25648_;
  wire _25649_;
  wire _25650_;
  wire _25651_;
  wire _25652_;
  wire _25653_;
  wire _25654_;
  wire _25655_;
  wire _25656_;
  wire _25657_;
  wire _25658_;
  wire _25659_;
  wire _25660_;
  wire _25661_;
  wire _25662_;
  wire _25663_;
  wire _25664_;
  wire _25665_;
  wire _25666_;
  wire _25667_;
  wire _25668_;
  wire _25669_;
  wire _25670_;
  wire _25671_;
  wire _25672_;
  wire _25673_;
  wire _25674_;
  wire _25675_;
  wire _25676_;
  wire _25677_;
  wire _25678_;
  wire _25679_;
  wire _25680_;
  wire _25681_;
  wire _25682_;
  wire _25683_;
  wire _25684_;
  wire _25685_;
  wire _25686_;
  wire _25687_;
  wire _25688_;
  wire _25689_;
  wire _25690_;
  wire _25691_;
  wire _25692_;
  wire _25693_;
  wire _25694_;
  wire _25695_;
  wire _25696_;
  wire _25697_;
  wire _25698_;
  wire _25699_;
  wire _25700_;
  wire _25701_;
  wire _25702_;
  wire _25703_;
  wire _25704_;
  wire _25705_;
  wire _25706_;
  wire _25707_;
  wire _25708_;
  wire _25709_;
  wire _25710_;
  wire _25711_;
  wire _25712_;
  wire _25713_;
  wire _25714_;
  wire _25715_;
  wire _25716_;
  wire _25717_;
  wire _25718_;
  wire _25719_;
  wire _25720_;
  wire _25721_;
  wire _25722_;
  wire _25723_;
  wire _25724_;
  wire _25725_;
  wire _25726_;
  wire _25727_;
  wire _25728_;
  wire _25729_;
  wire _25730_;
  wire _25731_;
  wire _25732_;
  wire _25733_;
  wire _25734_;
  wire _25735_;
  wire _25736_;
  wire _25737_;
  wire _25738_;
  wire _25739_;
  wire _25740_;
  wire _25741_;
  wire _25742_;
  wire _25743_;
  wire _25744_;
  wire _25745_;
  wire _25746_;
  wire _25747_;
  wire _25748_;
  wire _25749_;
  wire _25750_;
  wire _25751_;
  wire _25752_;
  wire _25753_;
  wire _25754_;
  wire _25755_;
  wire _25756_;
  wire _25757_;
  wire _25758_;
  wire _25759_;
  wire _25760_;
  wire _25761_;
  wire _25762_;
  wire _25763_;
  wire _25764_;
  wire _25765_;
  wire _25766_;
  wire _25767_;
  wire _25768_;
  wire _25769_;
  wire _25770_;
  wire _25771_;
  wire _25772_;
  wire _25773_;
  wire _25774_;
  wire _25775_;
  wire _25776_;
  wire _25777_;
  wire _25778_;
  wire _25779_;
  wire _25780_;
  wire _25781_;
  wire _25782_;
  wire _25783_;
  wire _25784_;
  wire _25785_;
  wire _25786_;
  wire _25787_;
  wire _25788_;
  wire _25789_;
  wire _25790_;
  wire _25791_;
  wire _25792_;
  wire _25793_;
  wire _25794_;
  wire _25795_;
  wire _25796_;
  wire _25797_;
  wire _25798_;
  wire _25799_;
  wire _25800_;
  wire _25801_;
  wire _25802_;
  wire _25803_;
  wire _25804_;
  wire _25805_;
  wire _25806_;
  wire _25807_;
  wire _25808_;
  wire _25809_;
  wire _25810_;
  wire _25811_;
  wire _25812_;
  wire _25813_;
  wire _25814_;
  wire _25815_;
  wire _25816_;
  wire _25817_;
  wire _25818_;
  wire _25819_;
  wire _25820_;
  wire _25821_;
  wire _25822_;
  wire _25823_;
  wire _25824_;
  wire _25825_;
  wire _25826_;
  wire _25827_;
  wire _25828_;
  wire _25829_;
  wire _25830_;
  wire _25831_;
  wire _25832_;
  wire _25833_;
  wire _25834_;
  wire _25835_;
  wire _25836_;
  wire _25837_;
  wire _25838_;
  wire _25839_;
  wire _25840_;
  wire _25841_;
  wire _25842_;
  wire _25843_;
  wire _25844_;
  wire _25845_;
  wire _25846_;
  wire _25847_;
  wire _25848_;
  wire _25849_;
  wire _25850_;
  wire _25851_;
  wire _25852_;
  wire _25853_;
  wire _25854_;
  wire _25855_;
  wire _25856_;
  wire _25857_;
  wire _25858_;
  wire _25859_;
  wire _25860_;
  wire _25861_;
  wire _25862_;
  wire _25863_;
  wire _25864_;
  wire _25865_;
  wire _25866_;
  wire _25867_;
  wire _25868_;
  wire _25869_;
  wire _25870_;
  wire _25871_;
  wire _25872_;
  wire _25873_;
  wire _25874_;
  wire _25875_;
  wire _25876_;
  wire _25877_;
  wire _25878_;
  wire _25879_;
  wire _25880_;
  wire _25881_;
  wire _25882_;
  wire _25883_;
  wire _25884_;
  wire _25885_;
  wire _25886_;
  wire _25887_;
  wire _25888_;
  wire _25889_;
  wire _25890_;
  wire _25891_;
  wire _25892_;
  wire _25893_;
  wire _25894_;
  wire _25895_;
  wire _25896_;
  wire _25897_;
  wire _25898_;
  wire _25899_;
  wire _25900_;
  wire _25901_;
  wire _25902_;
  wire _25903_;
  wire _25904_;
  wire _25905_;
  wire _25906_;
  wire _25907_;
  wire _25908_;
  wire _25909_;
  wire _25910_;
  wire _25911_;
  wire _25912_;
  wire _25913_;
  wire _25914_;
  wire _25915_;
  wire _25916_;
  wire _25917_;
  wire _25918_;
  wire _25919_;
  wire _25920_;
  wire _25921_;
  wire _25922_;
  wire _25923_;
  wire _25924_;
  wire _25925_;
  wire _25926_;
  wire _25927_;
  wire _25928_;
  wire _25929_;
  wire _25930_;
  wire _25931_;
  wire _25932_;
  wire _25933_;
  wire _25934_;
  wire _25935_;
  wire _25936_;
  wire _25937_;
  wire _25938_;
  wire _25939_;
  wire _25940_;
  wire _25941_;
  wire _25942_;
  wire _25943_;
  wire _25944_;
  wire _25945_;
  wire _25946_;
  wire _25947_;
  wire _25948_;
  wire _25949_;
  wire _25950_;
  wire _25951_;
  wire _25952_;
  wire _25953_;
  wire _25954_;
  wire _25955_;
  wire _25956_;
  wire _25957_;
  wire _25958_;
  wire _25959_;
  wire _25960_;
  wire _25961_;
  wire _25962_;
  wire _25963_;
  wire _25964_;
  wire _25965_;
  wire _25966_;
  wire _25967_;
  wire _25968_;
  wire _25969_;
  wire _25970_;
  wire _25971_;
  wire _25972_;
  wire _25973_;
  wire _25974_;
  wire _25975_;
  wire _25976_;
  wire _25977_;
  wire _25978_;
  wire _25979_;
  wire _25980_;
  wire _25981_;
  wire _25982_;
  wire _25983_;
  wire _25984_;
  wire _25985_;
  wire _25986_;
  wire _25987_;
  wire _25988_;
  wire _25989_;
  wire _25990_;
  wire _25991_;
  wire _25992_;
  wire _25993_;
  wire _25994_;
  wire _25995_;
  wire _25996_;
  wire _25997_;
  wire _25998_;
  wire _25999_;
  wire _26000_;
  wire _26001_;
  wire _26002_;
  wire _26003_;
  wire _26004_;
  wire _26005_;
  wire _26006_;
  wire _26007_;
  wire _26008_;
  wire _26009_;
  wire _26010_;
  wire _26011_;
  wire _26012_;
  wire _26013_;
  wire _26014_;
  wire _26015_;
  wire _26016_;
  wire _26017_;
  wire _26018_;
  wire _26019_;
  wire _26020_;
  wire _26021_;
  wire _26022_;
  wire _26023_;
  wire _26024_;
  wire _26025_;
  wire _26026_;
  wire _26027_;
  wire _26028_;
  wire _26029_;
  wire _26030_;
  wire _26031_;
  wire _26032_;
  wire _26033_;
  wire _26034_;
  wire _26035_;
  wire _26036_;
  wire _26037_;
  wire _26038_;
  wire _26039_;
  wire _26040_;
  wire _26041_;
  wire _26042_;
  wire _26043_;
  wire _26044_;
  wire _26045_;
  wire _26046_;
  wire _26047_;
  wire _26048_;
  wire _26049_;
  wire _26050_;
  wire _26051_;
  wire _26052_;
  wire _26053_;
  wire _26054_;
  wire _26055_;
  wire _26056_;
  wire _26057_;
  wire _26058_;
  wire _26059_;
  wire _26060_;
  wire _26061_;
  wire _26062_;
  wire _26063_;
  wire _26064_;
  wire _26065_;
  wire _26066_;
  wire _26067_;
  wire _26068_;
  wire _26069_;
  wire _26070_;
  wire _26071_;
  wire _26072_;
  wire _26073_;
  wire _26074_;
  wire _26075_;
  wire _26076_;
  wire _26077_;
  wire _26078_;
  wire _26079_;
  wire _26080_;
  wire _26081_;
  wire _26082_;
  wire _26083_;
  wire _26084_;
  wire _26085_;
  wire _26086_;
  wire _26087_;
  wire _26088_;
  wire _26089_;
  wire _26090_;
  wire _26091_;
  wire _26092_;
  wire _26093_;
  wire _26094_;
  wire _26095_;
  wire _26096_;
  wire _26097_;
  wire _26098_;
  wire _26099_;
  wire _26100_;
  wire _26101_;
  wire _26102_;
  wire _26103_;
  wire _26104_;
  wire _26105_;
  wire _26106_;
  wire _26107_;
  wire _26108_;
  wire _26109_;
  wire _26110_;
  wire _26111_;
  wire _26112_;
  wire _26113_;
  wire _26114_;
  wire _26115_;
  wire _26116_;
  wire _26117_;
  wire _26118_;
  wire _26119_;
  wire _26120_;
  wire _26121_;
  wire _26122_;
  wire _26123_;
  wire _26124_;
  wire _26125_;
  wire _26126_;
  wire _26127_;
  wire _26128_;
  wire _26129_;
  wire _26130_;
  wire _26131_;
  wire _26132_;
  wire _26133_;
  wire _26134_;
  wire _26135_;
  wire _26136_;
  wire _26137_;
  wire _26138_;
  wire _26139_;
  wire _26140_;
  wire _26141_;
  wire _26142_;
  wire _26143_;
  wire _26144_;
  wire _26145_;
  wire _26146_;
  wire _26147_;
  wire _26148_;
  wire _26149_;
  wire _26150_;
  wire _26151_;
  wire _26152_;
  wire _26153_;
  wire _26154_;
  wire _26155_;
  wire _26156_;
  wire _26157_;
  wire _26158_;
  wire _26159_;
  wire _26160_;
  wire _26161_;
  wire _26162_;
  wire _26163_;
  wire _26164_;
  wire _26165_;
  wire _26166_;
  wire _26167_;
  wire _26168_;
  wire _26169_;
  wire _26170_;
  wire _26171_;
  wire _26172_;
  wire _26173_;
  wire _26174_;
  wire _26175_;
  wire _26176_;
  wire _26177_;
  wire _26178_;
  wire _26179_;
  wire _26180_;
  wire _26181_;
  wire _26182_;
  wire _26183_;
  wire _26184_;
  wire _26185_;
  wire _26186_;
  wire _26187_;
  wire _26188_;
  wire _26189_;
  wire _26190_;
  wire _26191_;
  wire _26192_;
  wire _26193_;
  wire _26194_;
  wire _26195_;
  wire _26196_;
  wire _26197_;
  wire _26198_;
  wire _26199_;
  wire _26200_;
  wire _26201_;
  wire _26202_;
  wire _26203_;
  wire _26204_;
  wire _26205_;
  wire _26206_;
  wire _26207_;
  wire _26208_;
  wire _26209_;
  wire _26210_;
  wire _26211_;
  wire _26212_;
  wire _26213_;
  wire _26214_;
  wire _26215_;
  wire _26216_;
  wire _26217_;
  wire _26218_;
  wire _26219_;
  wire _26220_;
  wire _26221_;
  wire _26222_;
  wire _26223_;
  wire _26224_;
  wire _26225_;
  wire _26226_;
  wire _26227_;
  wire _26228_;
  wire _26229_;
  wire _26230_;
  wire _26231_;
  wire _26232_;
  wire _26233_;
  wire _26234_;
  wire _26235_;
  wire _26236_;
  wire _26237_;
  wire _26238_;
  wire _26239_;
  wire _26240_;
  wire _26241_;
  wire _26242_;
  wire _26243_;
  wire _26244_;
  wire _26245_;
  wire _26246_;
  wire _26247_;
  wire _26248_;
  wire _26249_;
  wire _26250_;
  wire _26251_;
  wire _26252_;
  wire _26253_;
  wire _26254_;
  wire _26255_;
  wire _26256_;
  wire _26257_;
  wire _26258_;
  wire _26259_;
  wire _26260_;
  wire _26261_;
  wire _26262_;
  wire _26263_;
  wire _26264_;
  wire _26265_;
  wire _26266_;
  wire _26267_;
  wire _26268_;
  wire _26269_;
  wire _26270_;
  wire _26271_;
  wire _26272_;
  wire _26273_;
  wire _26274_;
  wire _26275_;
  wire _26276_;
  wire _26277_;
  wire _26278_;
  wire _26279_;
  wire _26280_;
  wire _26281_;
  wire _26282_;
  wire _26283_;
  wire _26284_;
  wire _26285_;
  wire _26286_;
  wire _26287_;
  wire _26288_;
  wire _26289_;
  wire _26290_;
  wire _26291_;
  wire _26292_;
  wire _26293_;
  wire _26294_;
  wire _26295_;
  wire _26296_;
  wire _26297_;
  wire _26298_;
  wire _26299_;
  wire _26300_;
  wire _26301_;
  wire _26302_;
  wire _26303_;
  wire _26304_;
  wire _26305_;
  wire _26306_;
  wire _26307_;
  wire _26308_;
  wire _26309_;
  wire _26310_;
  wire _26311_;
  wire _26312_;
  wire _26313_;
  wire _26314_;
  wire _26315_;
  wire _26316_;
  wire _26317_;
  wire _26318_;
  wire _26319_;
  wire _26320_;
  wire _26321_;
  wire _26322_;
  wire _26323_;
  wire _26324_;
  wire _26325_;
  wire _26326_;
  wire _26327_;
  wire _26328_;
  wire _26329_;
  wire _26330_;
  wire _26331_;
  wire _26332_;
  wire _26333_;
  wire _26334_;
  wire _26335_;
  wire _26336_;
  wire _26337_;
  wire _26338_;
  wire _26339_;
  wire _26340_;
  wire _26341_;
  wire _26342_;
  wire _26343_;
  wire _26344_;
  wire _26345_;
  wire _26346_;
  wire _26347_;
  wire _26348_;
  wire _26349_;
  wire _26350_;
  wire _26351_;
  wire _26352_;
  wire _26353_;
  wire _26354_;
  wire _26355_;
  wire _26356_;
  wire _26357_;
  wire _26358_;
  wire _26359_;
  wire _26360_;
  wire _26361_;
  wire _26362_;
  wire _26363_;
  wire _26364_;
  wire _26365_;
  wire _26366_;
  wire _26367_;
  wire _26368_;
  wire _26369_;
  wire _26370_;
  wire _26371_;
  wire _26372_;
  wire _26373_;
  wire _26374_;
  wire _26375_;
  wire _26376_;
  wire _26377_;
  wire _26378_;
  wire _26379_;
  wire _26380_;
  wire _26381_;
  wire _26382_;
  wire _26383_;
  wire _26384_;
  wire _26385_;
  wire _26386_;
  wire _26387_;
  wire _26388_;
  wire _26389_;
  wire _26390_;
  wire _26391_;
  wire _26392_;
  wire _26393_;
  wire _26394_;
  wire _26395_;
  wire _26396_;
  wire _26397_;
  wire _26398_;
  wire _26399_;
  wire _26400_;
  wire _26401_;
  wire _26402_;
  wire _26403_;
  wire _26404_;
  wire _26405_;
  wire _26406_;
  wire _26407_;
  wire _26408_;
  wire _26409_;
  wire _26410_;
  wire _26411_;
  wire _26412_;
  wire _26413_;
  wire _26414_;
  wire _26415_;
  wire _26416_;
  wire _26417_;
  wire _26418_;
  wire _26419_;
  wire _26420_;
  wire _26421_;
  wire _26422_;
  wire _26423_;
  wire _26424_;
  wire _26425_;
  wire _26426_;
  wire _26427_;
  wire _26428_;
  wire _26429_;
  wire _26430_;
  wire _26431_;
  wire _26432_;
  wire _26433_;
  wire _26434_;
  wire _26435_;
  wire _26436_;
  wire _26437_;
  wire _26438_;
  wire _26439_;
  wire _26440_;
  wire _26441_;
  wire _26442_;
  wire _26443_;
  wire _26444_;
  wire _26445_;
  wire _26446_;
  wire _26447_;
  wire _26448_;
  wire _26449_;
  wire _26450_;
  wire _26451_;
  wire _26452_;
  wire _26453_;
  wire _26454_;
  wire _26455_;
  wire _26456_;
  wire _26457_;
  wire _26458_;
  wire _26459_;
  wire _26460_;
  wire _26461_;
  wire _26462_;
  wire _26463_;
  wire _26464_;
  wire _26465_;
  wire _26466_;
  wire _26467_;
  wire _26468_;
  wire _26469_;
  wire _26470_;
  wire _26471_;
  wire _26472_;
  wire _26473_;
  wire _26474_;
  wire _26475_;
  wire _26476_;
  wire _26477_;
  wire _26478_;
  wire _26479_;
  wire _26480_;
  wire _26481_;
  wire _26482_;
  wire _26483_;
  wire _26484_;
  wire _26485_;
  wire _26486_;
  wire _26487_;
  wire _26488_;
  wire _26489_;
  wire _26490_;
  wire _26491_;
  wire _26492_;
  wire _26493_;
  wire _26494_;
  wire _26495_;
  wire _26496_;
  wire _26497_;
  wire _26498_;
  wire _26499_;
  wire _26500_;
  wire _26501_;
  wire _26502_;
  wire _26503_;
  wire _26504_;
  wire _26505_;
  wire _26506_;
  wire _26507_;
  wire _26508_;
  wire _26509_;
  wire _26510_;
  wire _26511_;
  wire _26512_;
  wire _26513_;
  wire _26514_;
  wire _26515_;
  wire _26516_;
  wire _26517_;
  wire _26518_;
  wire _26519_;
  wire _26520_;
  wire _26521_;
  wire _26522_;
  wire _26523_;
  wire _26524_;
  wire _26525_;
  wire _26526_;
  wire _26527_;
  wire _26528_;
  wire _26529_;
  wire _26530_;
  wire _26531_;
  wire _26532_;
  wire _26533_;
  wire _26534_;
  wire _26535_;
  wire _26536_;
  wire _26537_;
  wire _26538_;
  wire _26539_;
  wire _26540_;
  wire _26541_;
  wire _26542_;
  wire _26543_;
  wire _26544_;
  wire _26545_;
  wire _26546_;
  wire _26547_;
  wire _26548_;
  wire _26549_;
  wire _26550_;
  wire _26551_;
  wire _26552_;
  wire _26553_;
  wire _26554_;
  wire _26555_;
  wire _26556_;
  wire _26557_;
  wire _26558_;
  wire _26559_;
  wire _26560_;
  wire _26561_;
  wire _26562_;
  wire _26563_;
  wire _26564_;
  wire _26565_;
  wire _26566_;
  wire _26567_;
  wire _26568_;
  wire _26569_;
  wire _26570_;
  wire _26571_;
  wire _26572_;
  wire _26573_;
  wire _26574_;
  wire _26575_;
  wire _26576_;
  wire _26577_;
  wire _26578_;
  wire _26579_;
  wire _26580_;
  wire _26581_;
  wire _26582_;
  wire _26583_;
  wire _26584_;
  wire _26585_;
  wire _26586_;
  wire _26587_;
  wire _26588_;
  wire _26589_;
  wire _26590_;
  wire _26591_;
  wire _26592_;
  wire _26593_;
  wire _26594_;
  wire _26595_;
  wire _26596_;
  wire _26597_;
  wire _26598_;
  wire _26599_;
  wire _26600_;
  wire _26601_;
  wire _26602_;
  wire _26603_;
  wire _26604_;
  wire _26605_;
  wire _26606_;
  wire _26607_;
  wire _26608_;
  wire _26609_;
  wire _26610_;
  wire _26611_;
  wire _26612_;
  wire _26613_;
  wire _26614_;
  wire _26615_;
  wire _26616_;
  wire _26617_;
  wire _26618_;
  wire _26619_;
  wire _26620_;
  wire _26621_;
  wire _26622_;
  wire _26623_;
  wire _26624_;
  wire _26625_;
  wire _26626_;
  wire _26627_;
  wire _26628_;
  wire _26629_;
  wire _26630_;
  wire _26631_;
  wire _26632_;
  wire _26633_;
  wire _26634_;
  wire _26635_;
  wire _26636_;
  wire _26637_;
  wire _26638_;
  wire _26639_;
  wire _26640_;
  wire _26641_;
  wire _26642_;
  wire _26643_;
  wire _26644_;
  wire _26645_;
  wire _26646_;
  wire _26647_;
  wire _26648_;
  wire _26649_;
  wire _26650_;
  wire _26651_;
  wire _26652_;
  wire _26653_;
  wire _26654_;
  wire _26655_;
  wire _26656_;
  wire _26657_;
  wire _26658_;
  wire _26659_;
  wire _26660_;
  wire _26661_;
  wire _26662_;
  wire _26663_;
  wire _26664_;
  wire _26665_;
  wire _26666_;
  wire _26667_;
  wire _26668_;
  wire _26669_;
  wire _26670_;
  wire _26671_;
  wire _26672_;
  wire _26673_;
  wire _26674_;
  wire _26675_;
  wire _26676_;
  wire _26677_;
  wire _26678_;
  wire _26679_;
  wire _26680_;
  wire _26681_;
  wire _26682_;
  wire _26683_;
  wire _26684_;
  wire _26685_;
  wire _26686_;
  wire _26687_;
  wire _26688_;
  wire _26689_;
  wire _26690_;
  wire _26691_;
  wire _26692_;
  wire _26693_;
  wire _26694_;
  wire _26695_;
  wire _26696_;
  wire _26697_;
  wire _26698_;
  wire _26699_;
  wire _26700_;
  wire _26701_;
  wire _26702_;
  wire _26703_;
  wire _26704_;
  wire _26705_;
  wire _26706_;
  wire _26707_;
  wire _26708_;
  wire _26709_;
  wire _26710_;
  wire _26711_;
  wire _26712_;
  wire _26713_;
  wire _26714_;
  wire _26715_;
  wire _26716_;
  wire _26717_;
  wire _26718_;
  wire _26719_;
  wire _26720_;
  wire _26721_;
  wire _26722_;
  wire _26723_;
  wire _26724_;
  wire _26725_;
  wire _26726_;
  wire _26727_;
  wire _26728_;
  wire _26729_;
  wire _26730_;
  wire _26731_;
  wire _26732_;
  wire _26733_;
  wire _26734_;
  wire _26735_;
  wire _26736_;
  wire _26737_;
  wire _26738_;
  wire _26739_;
  wire _26740_;
  wire _26741_;
  wire _26742_;
  wire _26743_;
  wire _26744_;
  wire _26745_;
  wire _26746_;
  wire _26747_;
  wire _26748_;
  wire _26749_;
  wire _26750_;
  wire _26751_;
  wire _26752_;
  wire _26753_;
  wire _26754_;
  wire _26755_;
  wire _26756_;
  wire _26757_;
  wire _26758_;
  wire _26759_;
  wire _26760_;
  wire _26761_;
  wire _26762_;
  wire _26763_;
  wire _26764_;
  wire _26765_;
  wire _26766_;
  wire _26767_;
  wire _26768_;
  wire _26769_;
  wire _26770_;
  wire _26771_;
  wire _26772_;
  wire _26773_;
  wire _26774_;
  wire _26775_;
  wire _26776_;
  wire _26777_;
  wire _26778_;
  wire _26779_;
  wire _26780_;
  wire _26781_;
  wire _26782_;
  wire _26783_;
  wire _26784_;
  wire _26785_;
  wire _26786_;
  wire _26787_;
  wire _26788_;
  wire _26789_;
  wire _26790_;
  wire _26791_;
  wire _26792_;
  wire _26793_;
  wire _26794_;
  wire _26795_;
  wire _26796_;
  wire _26797_;
  wire _26798_;
  wire _26799_;
  wire _26800_;
  wire _26801_;
  wire _26802_;
  wire _26803_;
  wire _26804_;
  wire _26805_;
  wire _26806_;
  wire _26807_;
  wire _26808_;
  wire _26809_;
  wire _26810_;
  wire _26811_;
  wire _26812_;
  wire _26813_;
  wire _26814_;
  wire _26815_;
  wire _26816_;
  wire _26817_;
  wire _26818_;
  wire _26819_;
  wire _26820_;
  wire _26821_;
  wire _26822_;
  wire _26823_;
  wire _26824_;
  wire _26825_;
  wire _26826_;
  wire _26827_;
  wire _26828_;
  wire _26829_;
  wire _26830_;
  wire _26831_;
  wire _26832_;
  wire _26833_;
  wire _26834_;
  wire _26835_;
  wire _26836_;
  wire _26837_;
  wire _26838_;
  wire _26839_;
  wire _26840_;
  wire _26841_;
  wire _26842_;
  wire _26843_;
  wire _26844_;
  wire _26845_;
  wire _26846_;
  wire _26847_;
  wire _26848_;
  wire _26849_;
  wire _26850_;
  wire _26851_;
  wire _26852_;
  wire _26853_;
  wire _26854_;
  wire _26855_;
  wire _26856_;
  wire _26857_;
  wire _26858_;
  wire _26859_;
  wire _26860_;
  wire _26861_;
  wire _26862_;
  wire _26863_;
  wire _26864_;
  wire _26865_;
  wire _26866_;
  wire _26867_;
  wire _26868_;
  wire _26869_;
  wire _26870_;
  wire _26871_;
  wire _26872_;
  wire _26873_;
  wire _26874_;
  wire _26875_;
  wire _26876_;
  wire _26877_;
  wire _26878_;
  wire _26879_;
  wire _26880_;
  wire _26881_;
  wire _26882_;
  wire _26883_;
  wire _26884_;
  wire _26885_;
  wire _26886_;
  wire _26887_;
  wire _26888_;
  wire _26889_;
  wire _26890_;
  wire _26891_;
  wire _26892_;
  wire _26893_;
  wire _26894_;
  wire _26895_;
  wire _26896_;
  wire _26897_;
  wire _26898_;
  wire _26899_;
  wire _26900_;
  wire _26901_;
  wire _26902_;
  wire _26903_;
  wire _26904_;
  wire _26905_;
  wire _26906_;
  wire _26907_;
  wire _26908_;
  wire _26909_;
  wire _26910_;
  wire _26911_;
  wire _26912_;
  wire _26913_;
  wire _26914_;
  wire _26915_;
  wire _26916_;
  wire _26917_;
  wire _26918_;
  wire _26919_;
  wire _26920_;
  wire _26921_;
  wire _26922_;
  wire _26923_;
  wire _26924_;
  wire _26925_;
  wire _26926_;
  wire _26927_;
  wire _26928_;
  wire _26929_;
  wire _26930_;
  wire _26931_;
  wire _26932_;
  wire _26933_;
  wire _26934_;
  wire _26935_;
  wire _26936_;
  wire _26937_;
  wire _26938_;
  wire _26939_;
  wire _26940_;
  wire _26941_;
  wire _26942_;
  wire _26943_;
  wire _26944_;
  wire _26945_;
  wire _26946_;
  wire _26947_;
  wire _26948_;
  wire _26949_;
  wire _26950_;
  wire _26951_;
  wire _26952_;
  wire _26953_;
  wire _26954_;
  wire _26955_;
  wire _26956_;
  wire _26957_;
  wire _26958_;
  wire _26959_;
  wire _26960_;
  wire _26961_;
  wire _26962_;
  wire _26963_;
  wire _26964_;
  wire _26965_;
  wire _26966_;
  wire _26967_;
  wire _26968_;
  wire _26969_;
  wire _26970_;
  wire _26971_;
  wire _26972_;
  wire _26973_;
  wire _26974_;
  wire _26975_;
  wire _26976_;
  wire _26977_;
  wire _26978_;
  wire _26979_;
  wire _26980_;
  wire _26981_;
  wire _26982_;
  wire _26983_;
  wire _26984_;
  wire _26985_;
  wire _26986_;
  wire _26987_;
  wire _26988_;
  wire _26989_;
  wire _26990_;
  wire _26991_;
  wire _26992_;
  wire _26993_;
  wire _26994_;
  wire _26995_;
  wire _26996_;
  wire _26997_;
  wire _26998_;
  wire _26999_;
  wire _27000_;
  wire _27001_;
  wire _27002_;
  wire _27003_;
  wire _27004_;
  wire _27005_;
  wire _27006_;
  wire _27007_;
  wire _27008_;
  wire _27009_;
  wire _27010_;
  wire _27011_;
  wire _27012_;
  wire _27013_;
  wire _27014_;
  wire _27015_;
  wire _27016_;
  wire _27017_;
  wire _27018_;
  wire _27019_;
  wire _27020_;
  wire _27021_;
  wire _27022_;
  wire _27023_;
  wire _27024_;
  wire _27025_;
  wire _27026_;
  wire _27027_;
  wire _27028_;
  wire _27029_;
  wire _27030_;
  wire _27031_;
  wire _27032_;
  wire _27033_;
  wire _27034_;
  wire _27035_;
  wire _27036_;
  wire _27037_;
  wire _27038_;
  wire _27039_;
  wire _27040_;
  wire _27041_;
  wire _27042_;
  wire _27043_;
  wire _27044_;
  wire _27045_;
  wire _27046_;
  wire _27047_;
  wire _27048_;
  wire _27049_;
  wire _27050_;
  wire _27051_;
  wire _27052_;
  wire _27053_;
  wire _27054_;
  wire _27055_;
  wire _27056_;
  wire _27057_;
  wire _27058_;
  wire _27059_;
  wire _27060_;
  wire _27061_;
  wire _27062_;
  wire _27063_;
  wire _27064_;
  wire _27065_;
  wire _27066_;
  wire _27067_;
  wire _27068_;
  wire _27069_;
  wire _27070_;
  wire _27071_;
  wire _27072_;
  wire _27073_;
  wire _27074_;
  wire _27075_;
  wire _27076_;
  wire _27077_;
  wire _27078_;
  wire _27079_;
  wire _27080_;
  wire _27081_;
  wire _27082_;
  wire _27083_;
  wire _27084_;
  wire _27085_;
  wire _27086_;
  wire _27087_;
  wire _27088_;
  wire _27089_;
  wire _27090_;
  wire _27091_;
  wire _27092_;
  wire _27093_;
  wire _27094_;
  wire _27095_;
  wire _27096_;
  wire _27097_;
  wire _27098_;
  wire _27099_;
  wire _27100_;
  wire _27101_;
  wire _27102_;
  wire _27103_;
  wire _27104_;
  wire _27105_;
  wire _27106_;
  wire _27107_;
  wire _27108_;
  wire _27109_;
  wire _27110_;
  wire _27111_;
  wire _27112_;
  wire _27113_;
  wire _27114_;
  wire _27115_;
  wire _27116_;
  wire _27117_;
  wire _27118_;
  wire _27119_;
  wire _27120_;
  wire _27121_;
  wire _27122_;
  wire _27123_;
  wire _27124_;
  wire _27125_;
  wire _27126_;
  wire _27127_;
  wire _27128_;
  wire _27129_;
  wire _27130_;
  wire _27131_;
  wire _27132_;
  wire _27133_;
  wire _27134_;
  wire _27135_;
  wire _27136_;
  wire _27137_;
  wire _27138_;
  wire _27139_;
  wire _27140_;
  wire _27141_;
  wire _27142_;
  wire _27143_;
  wire _27144_;
  wire _27145_;
  wire _27146_;
  wire _27147_;
  wire _27148_;
  wire _27149_;
  wire _27150_;
  wire _27151_;
  wire _27152_;
  wire _27153_;
  wire _27154_;
  wire _27155_;
  wire _27156_;
  wire _27157_;
  wire _27158_;
  wire _27159_;
  wire _27160_;
  wire _27161_;
  wire _27162_;
  wire _27163_;
  wire _27164_;
  wire _27165_;
  wire _27166_;
  wire _27167_;
  wire _27168_;
  wire _27169_;
  wire _27170_;
  wire _27171_;
  wire _27172_;
  wire _27173_;
  wire _27174_;
  wire _27175_;
  wire _27176_;
  wire _27177_;
  wire _27178_;
  wire _27179_;
  wire _27180_;
  wire _27181_;
  wire _27182_;
  wire _27183_;
  wire _27184_;
  wire _27185_;
  wire _27186_;
  wire _27187_;
  wire _27188_;
  wire _27189_;
  wire _27190_;
  wire _27191_;
  wire _27192_;
  wire _27193_;
  wire _27194_;
  wire _27195_;
  wire _27196_;
  wire _27197_;
  wire _27198_;
  wire _27199_;
  wire _27200_;
  wire _27201_;
  wire _27202_;
  wire _27203_;
  wire _27204_;
  wire _27205_;
  wire _27206_;
  wire _27207_;
  wire _27208_;
  wire _27209_;
  wire _27210_;
  wire _27211_;
  wire _27212_;
  wire _27213_;
  wire _27214_;
  wire _27215_;
  wire _27216_;
  wire _27217_;
  wire _27218_;
  wire _27219_;
  wire _27220_;
  wire _27221_;
  wire _27222_;
  wire _27223_;
  wire _27224_;
  wire _27225_;
  wire _27226_;
  wire _27227_;
  wire _27228_;
  wire _27229_;
  wire _27230_;
  wire _27231_;
  wire _27232_;
  wire _27233_;
  wire _27234_;
  wire _27235_;
  wire _27236_;
  wire _27237_;
  wire _27238_;
  wire _27239_;
  wire _27240_;
  wire _27241_;
  wire _27242_;
  wire _27243_;
  wire _27244_;
  wire _27245_;
  wire _27246_;
  wire _27247_;
  wire _27248_;
  wire _27249_;
  wire _27250_;
  wire _27251_;
  wire _27252_;
  wire _27253_;
  wire _27254_;
  wire _27255_;
  wire _27256_;
  wire _27257_;
  wire _27258_;
  wire _27259_;
  wire _27260_;
  wire _27261_;
  wire _27262_;
  wire _27263_;
  wire _27264_;
  wire _27265_;
  wire _27266_;
  wire _27267_;
  wire _27268_;
  wire _27269_;
  wire _27270_;
  wire _27271_;
  wire _27272_;
  wire _27273_;
  wire _27274_;
  wire _27275_;
  wire _27276_;
  wire _27277_;
  wire _27278_;
  wire _27279_;
  wire _27280_;
  wire _27281_;
  wire _27282_;
  wire _27283_;
  wire _27284_;
  wire _27285_;
  wire _27286_;
  wire _27287_;
  wire _27288_;
  wire _27289_;
  wire _27290_;
  wire _27291_;
  wire _27292_;
  wire _27293_;
  wire _27294_;
  wire _27295_;
  wire _27296_;
  wire _27297_;
  wire _27298_;
  wire _27299_;
  wire _27300_;
  wire _27301_;
  wire _27302_;
  wire _27303_;
  wire _27304_;
  wire _27305_;
  wire _27306_;
  wire _27307_;
  wire _27308_;
  wire _27309_;
  wire _27310_;
  wire _27311_;
  wire _27312_;
  wire _27313_;
  wire _27314_;
  wire _27315_;
  wire _27316_;
  wire _27317_;
  wire _27318_;
  wire _27319_;
  wire _27320_;
  wire _27321_;
  wire _27322_;
  wire _27323_;
  wire _27324_;
  wire _27325_;
  wire _27326_;
  wire _27327_;
  wire _27328_;
  wire _27329_;
  wire _27330_;
  wire _27331_;
  wire _27332_;
  wire _27333_;
  wire _27334_;
  wire _27335_;
  wire _27336_;
  wire _27337_;
  wire _27338_;
  wire _27339_;
  wire _27340_;
  wire _27341_;
  wire _27342_;
  wire _27343_;
  wire _27344_;
  wire _27345_;
  wire _27346_;
  wire _27347_;
  wire _27348_;
  wire _27349_;
  wire _27350_;
  wire _27351_;
  wire _27352_;
  wire _27353_;
  wire _27354_;
  wire _27355_;
  wire _27356_;
  wire _27357_;
  wire _27358_;
  wire _27359_;
  wire _27360_;
  wire _27361_;
  wire _27362_;
  wire _27363_;
  wire _27364_;
  wire _27365_;
  wire _27366_;
  wire _27367_;
  wire _27368_;
  wire _27369_;
  wire _27370_;
  wire _27371_;
  wire _27372_;
  wire _27373_;
  wire _27374_;
  wire _27375_;
  wire _27376_;
  wire _27377_;
  wire _27378_;
  wire _27379_;
  wire _27380_;
  wire _27381_;
  wire _27382_;
  wire _27383_;
  wire _27384_;
  wire _27385_;
  wire _27386_;
  wire _27387_;
  wire _27388_;
  wire _27389_;
  wire _27390_;
  wire _27391_;
  wire _27392_;
  wire _27393_;
  wire _27394_;
  wire _27395_;
  wire _27396_;
  wire _27397_;
  wire _27398_;
  wire _27399_;
  wire _27400_;
  wire _27401_;
  wire _27402_;
  wire _27403_;
  wire _27404_;
  wire _27405_;
  wire _27406_;
  wire _27407_;
  wire _27408_;
  wire _27409_;
  wire _27410_;
  wire _27411_;
  wire _27412_;
  wire _27413_;
  wire _27414_;
  wire _27415_;
  wire _27416_;
  wire _27417_;
  wire _27418_;
  wire _27419_;
  wire _27420_;
  wire _27421_;
  wire _27422_;
  wire _27423_;
  wire _27424_;
  wire _27425_;
  wire _27426_;
  wire _27427_;
  wire _27428_;
  wire _27429_;
  wire _27430_;
  wire _27431_;
  wire _27432_;
  wire _27433_;
  wire _27434_;
  wire _27435_;
  wire _27436_;
  wire _27437_;
  wire _27438_;
  wire _27439_;
  wire _27440_;
  wire _27441_;
  wire _27442_;
  wire _27443_;
  wire _27444_;
  wire _27445_;
  wire _27446_;
  wire _27447_;
  wire _27448_;
  wire _27449_;
  wire _27450_;
  wire _27451_;
  wire _27452_;
  wire _27453_;
  wire _27454_;
  wire _27455_;
  wire _27456_;
  wire _27457_;
  wire _27458_;
  wire _27459_;
  wire _27460_;
  wire _27461_;
  wire _27462_;
  wire _27463_;
  wire _27464_;
  wire _27465_;
  wire _27466_;
  wire _27467_;
  wire _27468_;
  wire _27469_;
  wire _27470_;
  wire _27471_;
  wire _27472_;
  wire _27473_;
  wire _27474_;
  wire _27475_;
  wire _27476_;
  wire _27477_;
  wire _27478_;
  wire _27479_;
  wire _27480_;
  wire _27481_;
  wire _27482_;
  wire _27483_;
  wire _27484_;
  wire _27485_;
  wire _27486_;
  wire _27487_;
  wire _27488_;
  wire _27489_;
  wire _27490_;
  wire _27491_;
  wire _27492_;
  wire _27493_;
  wire _27494_;
  wire _27495_;
  wire _27496_;
  wire _27497_;
  wire _27498_;
  wire _27499_;
  wire _27500_;
  wire _27501_;
  wire _27502_;
  wire _27503_;
  wire _27504_;
  wire _27505_;
  wire _27506_;
  wire _27507_;
  wire _27508_;
  wire _27509_;
  wire _27510_;
  wire _27511_;
  wire _27512_;
  wire _27513_;
  wire _27514_;
  wire _27515_;
  wire _27516_;
  wire _27517_;
  wire _27518_;
  wire _27519_;
  wire _27520_;
  wire _27521_;
  wire _27522_;
  wire _27523_;
  wire _27524_;
  wire _27525_;
  wire _27526_;
  wire _27527_;
  wire _27528_;
  wire _27529_;
  wire _27530_;
  wire _27531_;
  wire _27532_;
  wire _27533_;
  wire _27534_;
  wire _27535_;
  wire _27536_;
  wire _27537_;
  wire _27538_;
  wire _27539_;
  wire _27540_;
  wire _27541_;
  wire _27542_;
  wire _27543_;
  wire _27544_;
  wire _27545_;
  wire _27546_;
  wire _27547_;
  wire _27548_;
  wire _27549_;
  wire _27550_;
  wire _27551_;
  wire _27552_;
  wire _27553_;
  wire _27554_;
  wire _27555_;
  wire _27556_;
  wire _27557_;
  wire _27558_;
  wire _27559_;
  wire _27560_;
  wire _27561_;
  wire _27562_;
  wire _27563_;
  wire _27564_;
  wire _27565_;
  wire _27566_;
  wire _27567_;
  wire _27568_;
  wire _27569_;
  wire _27570_;
  wire _27571_;
  wire _27572_;
  wire _27573_;
  wire _27574_;
  wire _27575_;
  wire _27576_;
  wire _27577_;
  wire _27578_;
  wire _27579_;
  wire _27580_;
  wire _27581_;
  wire _27582_;
  wire _27583_;
  wire _27584_;
  wire _27585_;
  wire _27586_;
  wire _27587_;
  wire _27588_;
  wire _27589_;
  wire _27590_;
  wire _27591_;
  wire _27592_;
  wire _27593_;
  wire _27594_;
  wire _27595_;
  wire _27596_;
  wire _27597_;
  wire _27598_;
  wire _27599_;
  wire _27600_;
  wire _27601_;
  wire _27602_;
  wire _27603_;
  wire _27604_;
  wire _27605_;
  wire _27606_;
  wire _27607_;
  wire _27608_;
  wire _27609_;
  wire _27610_;
  wire _27611_;
  wire _27612_;
  wire _27613_;
  wire _27614_;
  wire _27615_;
  wire _27616_;
  wire _27617_;
  wire _27618_;
  wire _27619_;
  wire _27620_;
  wire _27621_;
  wire _27622_;
  wire _27623_;
  wire _27624_;
  wire _27625_;
  wire _27626_;
  wire _27627_;
  wire _27628_;
  wire _27629_;
  wire _27630_;
  wire _27631_;
  wire _27632_;
  wire _27633_;
  wire _27634_;
  wire _27635_;
  wire _27636_;
  wire _27637_;
  wire _27638_;
  wire _27639_;
  wire _27640_;
  wire _27641_;
  wire _27642_;
  wire _27643_;
  wire _27644_;
  wire _27645_;
  wire _27646_;
  wire _27647_;
  wire _27648_;
  wire _27649_;
  wire _27650_;
  wire _27651_;
  wire _27652_;
  wire _27653_;
  wire _27654_;
  wire _27655_;
  wire _27656_;
  wire _27657_;
  wire _27658_;
  wire _27659_;
  wire _27660_;
  wire _27661_;
  wire _27662_;
  wire _27663_;
  wire _27664_;
  wire _27665_;
  wire _27666_;
  wire _27667_;
  wire _27668_;
  wire _27669_;
  wire _27670_;
  wire _27671_;
  wire _27672_;
  wire _27673_;
  wire _27674_;
  wire _27675_;
  wire _27676_;
  wire _27677_;
  wire _27678_;
  wire _27679_;
  wire _27680_;
  wire _27681_;
  wire _27682_;
  wire _27683_;
  wire _27684_;
  wire _27685_;
  wire _27686_;
  wire _27687_;
  wire _27688_;
  wire _27689_;
  wire _27690_;
  wire _27691_;
  wire _27692_;
  wire _27693_;
  wire _27694_;
  wire _27695_;
  wire _27696_;
  wire _27697_;
  wire _27698_;
  wire _27699_;
  wire _27700_;
  wire _27701_;
  wire _27702_;
  wire _27703_;
  wire _27704_;
  wire _27705_;
  wire _27706_;
  wire _27707_;
  wire _27708_;
  wire _27709_;
  wire _27710_;
  wire _27711_;
  wire _27712_;
  wire _27713_;
  wire _27714_;
  wire _27715_;
  wire _27716_;
  wire _27717_;
  wire _27718_;
  wire _27719_;
  wire _27720_;
  wire _27721_;
  wire _27722_;
  wire _27723_;
  wire _27724_;
  wire _27725_;
  wire _27726_;
  wire _27727_;
  wire _27728_;
  wire _27729_;
  wire _27730_;
  wire _27731_;
  wire _27732_;
  wire _27733_;
  wire _27734_;
  wire _27735_;
  wire _27736_;
  wire _27737_;
  wire _27738_;
  wire _27739_;
  wire _27740_;
  wire _27741_;
  wire _27742_;
  wire _27743_;
  wire _27744_;
  wire _27745_;
  wire _27746_;
  wire _27747_;
  wire _27748_;
  wire _27749_;
  wire _27750_;
  wire _27751_;
  wire _27752_;
  wire _27753_;
  wire _27754_;
  wire _27755_;
  wire _27756_;
  wire _27757_;
  wire _27758_;
  wire _27759_;
  wire _27760_;
  wire _27761_;
  wire _27762_;
  wire _27763_;
  wire _27764_;
  wire _27765_;
  wire _27766_;
  wire _27767_;
  wire _27768_;
  wire _27769_;
  wire _27770_;
  wire _27771_;
  wire _27772_;
  wire _27773_;
  wire _27774_;
  wire _27775_;
  wire _27776_;
  wire _27777_;
  wire _27778_;
  wire _27779_;
  wire _27780_;
  wire _27781_;
  wire _27782_;
  wire _27783_;
  wire _27784_;
  wire _27785_;
  wire _27786_;
  wire _27787_;
  wire _27788_;
  wire _27789_;
  wire _27790_;
  wire _27791_;
  wire _27792_;
  wire _27793_;
  wire _27794_;
  wire _27795_;
  wire _27796_;
  wire _27797_;
  wire _27798_;
  wire _27799_;
  wire _27800_;
  wire _27801_;
  wire _27802_;
  wire _27803_;
  wire _27804_;
  wire _27805_;
  wire _27806_;
  wire _27807_;
  wire _27808_;
  wire _27809_;
  wire _27810_;
  wire _27811_;
  wire _27812_;
  wire _27813_;
  wire _27814_;
  wire _27815_;
  wire _27816_;
  wire _27817_;
  wire _27818_;
  wire _27819_;
  wire _27820_;
  wire _27821_;
  wire _27822_;
  wire _27823_;
  wire _27824_;
  wire _27825_;
  wire _27826_;
  wire _27827_;
  wire _27828_;
  wire _27829_;
  wire _27830_;
  wire _27831_;
  wire _27832_;
  wire _27833_;
  wire _27834_;
  wire _27835_;
  wire _27836_;
  wire _27837_;
  wire _27838_;
  wire _27839_;
  wire _27840_;
  wire _27841_;
  wire _27842_;
  wire _27843_;
  wire _27844_;
  wire _27845_;
  wire _27846_;
  wire _27847_;
  wire _27848_;
  wire _27849_;
  wire _27850_;
  wire _27851_;
  wire _27852_;
  wire _27853_;
  wire _27854_;
  wire _27855_;
  wire _27856_;
  wire _27857_;
  wire _27858_;
  wire _27859_;
  wire _27860_;
  wire _27861_;
  wire _27862_;
  wire _27863_;
  wire _27864_;
  wire _27865_;
  wire _27866_;
  wire _27867_;
  wire _27868_;
  wire _27869_;
  wire _27870_;
  wire _27871_;
  wire _27872_;
  wire _27873_;
  wire _27874_;
  wire _27875_;
  wire _27876_;
  wire _27877_;
  wire _27878_;
  wire _27879_;
  wire _27880_;
  wire _27881_;
  wire _27882_;
  wire _27883_;
  wire _27884_;
  wire _27885_;
  wire _27886_;
  wire _27887_;
  wire _27888_;
  wire _27889_;
  wire _27890_;
  wire _27891_;
  wire _27892_;
  wire _27893_;
  wire _27894_;
  wire _27895_;
  wire _27896_;
  wire _27897_;
  wire _27898_;
  wire _27899_;
  wire _27900_;
  wire _27901_;
  wire _27902_;
  wire _27903_;
  wire _27904_;
  wire _27905_;
  wire _27906_;
  wire _27907_;
  wire _27908_;
  wire _27909_;
  wire _27910_;
  wire _27911_;
  wire _27912_;
  wire _27913_;
  wire _27914_;
  wire _27915_;
  wire _27916_;
  wire _27917_;
  wire _27918_;
  wire _27919_;
  wire _27920_;
  wire _27921_;
  wire _27922_;
  wire _27923_;
  wire _27924_;
  wire _27925_;
  wire _27926_;
  wire _27927_;
  wire _27928_;
  wire _27929_;
  wire _27930_;
  wire _27931_;
  wire _27932_;
  wire _27933_;
  wire _27934_;
  wire _27935_;
  wire _27936_;
  wire _27937_;
  wire _27938_;
  wire _27939_;
  wire _27940_;
  wire _27941_;
  wire _27942_;
  wire _27943_;
  wire _27944_;
  wire _27945_;
  wire _27946_;
  wire _27947_;
  wire _27948_;
  wire _27949_;
  wire _27950_;
  wire _27951_;
  wire _27952_;
  wire _27953_;
  wire _27954_;
  wire _27955_;
  wire _27956_;
  wire _27957_;
  wire _27958_;
  wire _27959_;
  wire _27960_;
  wire _27961_;
  wire _27962_;
  wire _27963_;
  wire _27964_;
  wire _27965_;
  wire _27966_;
  wire _27967_;
  wire _27968_;
  wire _27969_;
  wire _27970_;
  wire _27971_;
  wire _27972_;
  wire _27973_;
  wire _27974_;
  wire _27975_;
  wire _27976_;
  wire _27977_;
  wire _27978_;
  wire _27979_;
  wire _27980_;
  wire _27981_;
  wire _27982_;
  wire _27983_;
  wire _27984_;
  wire _27985_;
  wire _27986_;
  wire _27987_;
  wire _27988_;
  wire _27989_;
  wire _27990_;
  wire _27991_;
  wire _27992_;
  wire _27993_;
  wire _27994_;
  wire _27995_;
  wire _27996_;
  wire _27997_;
  wire _27998_;
  wire _27999_;
  wire _28000_;
  wire _28001_;
  wire _28002_;
  wire _28003_;
  wire _28004_;
  wire _28005_;
  wire _28006_;
  wire _28007_;
  wire _28008_;
  wire _28009_;
  wire _28010_;
  wire _28011_;
  wire _28012_;
  wire _28013_;
  wire _28014_;
  wire _28015_;
  wire _28016_;
  wire _28017_;
  wire _28018_;
  wire _28019_;
  wire _28020_;
  wire _28021_;
  wire _28022_;
  wire _28023_;
  wire _28024_;
  wire _28025_;
  wire _28026_;
  wire _28027_;
  wire _28028_;
  wire _28029_;
  wire _28030_;
  wire _28031_;
  wire _28032_;
  wire _28033_;
  wire _28034_;
  wire _28035_;
  wire _28036_;
  wire _28037_;
  wire _28038_;
  wire _28039_;
  wire _28040_;
  wire _28041_;
  wire _28042_;
  wire _28043_;
  wire _28044_;
  wire _28045_;
  wire _28046_;
  wire _28047_;
  wire _28048_;
  wire _28049_;
  wire _28050_;
  wire _28051_;
  wire _28052_;
  wire _28053_;
  wire _28054_;
  wire _28055_;
  wire _28056_;
  wire _28057_;
  wire _28058_;
  wire _28059_;
  wire _28060_;
  wire _28061_;
  wire _28062_;
  wire _28063_;
  wire _28064_;
  wire _28065_;
  wire _28066_;
  wire _28067_;
  wire _28068_;
  wire _28069_;
  wire _28070_;
  wire _28071_;
  wire _28072_;
  wire _28073_;
  wire _28074_;
  wire _28075_;
  wire _28076_;
  wire _28077_;
  wire _28078_;
  wire _28079_;
  wire _28080_;
  wire _28081_;
  wire _28082_;
  wire _28083_;
  wire _28084_;
  wire _28085_;
  wire _28086_;
  wire _28087_;
  wire _28088_;
  wire _28089_;
  wire _28090_;
  wire _28091_;
  wire _28092_;
  wire _28093_;
  wire _28094_;
  wire _28095_;
  wire _28096_;
  wire _28097_;
  wire _28098_;
  wire _28099_;
  wire _28100_;
  wire _28101_;
  wire _28102_;
  wire _28103_;
  wire _28104_;
  wire _28105_;
  wire _28106_;
  wire _28107_;
  wire _28108_;
  wire _28109_;
  wire _28110_;
  wire _28111_;
  wire _28112_;
  wire _28113_;
  wire _28114_;
  wire _28115_;
  wire _28116_;
  wire _28117_;
  wire _28118_;
  wire _28119_;
  wire _28120_;
  wire _28121_;
  wire _28122_;
  wire _28123_;
  wire _28124_;
  wire _28125_;
  wire _28126_;
  wire _28127_;
  wire _28128_;
  wire _28129_;
  wire _28130_;
  wire _28131_;
  wire _28132_;
  wire _28133_;
  wire _28134_;
  wire _28135_;
  wire _28136_;
  wire _28137_;
  wire _28138_;
  wire _28139_;
  wire _28140_;
  wire _28141_;
  wire _28142_;
  wire _28143_;
  wire _28144_;
  wire _28145_;
  wire _28146_;
  wire _28147_;
  wire _28148_;
  wire _28149_;
  wire _28150_;
  wire _28151_;
  wire _28152_;
  wire _28153_;
  wire _28154_;
  wire _28155_;
  wire _28156_;
  wire _28157_;
  wire _28158_;
  wire _28159_;
  wire _28160_;
  wire _28161_;
  wire _28162_;
  wire _28163_;
  wire _28164_;
  wire _28165_;
  wire _28166_;
  wire _28167_;
  wire _28168_;
  wire _28169_;
  wire _28170_;
  wire _28171_;
  wire _28172_;
  wire _28173_;
  wire _28174_;
  wire _28175_;
  wire _28176_;
  wire _28177_;
  wire _28178_;
  wire _28179_;
  wire _28180_;
  wire _28181_;
  wire _28182_;
  wire _28183_;
  wire _28184_;
  wire _28185_;
  wire _28186_;
  wire _28187_;
  wire _28188_;
  wire _28189_;
  wire _28190_;
  wire _28191_;
  wire _28192_;
  wire _28193_;
  wire _28194_;
  wire _28195_;
  wire _28196_;
  wire _28197_;
  wire _28198_;
  wire _28199_;
  wire _28200_;
  wire _28201_;
  wire _28202_;
  wire _28203_;
  wire _28204_;
  wire _28205_;
  wire _28206_;
  wire _28207_;
  wire _28208_;
  wire _28209_;
  wire _28210_;
  wire _28211_;
  wire _28212_;
  wire _28213_;
  wire _28214_;
  wire _28215_;
  wire _28216_;
  wire _28217_;
  wire _28218_;
  wire _28219_;
  wire _28220_;
  wire _28221_;
  wire _28222_;
  wire _28223_;
  wire _28224_;
  wire _28225_;
  wire _28226_;
  wire _28227_;
  wire _28228_;
  wire _28229_;
  wire _28230_;
  wire _28231_;
  wire _28232_;
  wire _28233_;
  wire _28234_;
  wire _28235_;
  wire _28236_;
  wire _28237_;
  wire _28238_;
  wire _28239_;
  wire _28240_;
  wire _28241_;
  wire _28242_;
  wire _28243_;
  wire _28244_;
  wire _28245_;
  wire _28246_;
  wire _28247_;
  wire _28248_;
  wire _28249_;
  wire _28250_;
  wire _28251_;
  wire _28252_;
  wire _28253_;
  wire _28254_;
  wire _28255_;
  wire _28256_;
  wire _28257_;
  wire _28258_;
  wire _28259_;
  wire _28260_;
  wire _28261_;
  wire _28262_;
  wire _28263_;
  wire _28264_;
  wire _28265_;
  wire _28266_;
  wire _28267_;
  wire _28268_;
  wire _28269_;
  wire _28270_;
  wire _28271_;
  wire _28272_;
  wire _28273_;
  wire _28274_;
  wire _28275_;
  wire _28276_;
  wire _28277_;
  wire _28278_;
  wire _28279_;
  wire _28280_;
  wire _28281_;
  wire _28282_;
  wire _28283_;
  wire _28284_;
  wire _28285_;
  wire _28286_;
  wire _28287_;
  wire _28288_;
  wire _28289_;
  wire _28290_;
  wire _28291_;
  wire _28292_;
  wire _28293_;
  wire _28294_;
  wire _28295_;
  wire _28296_;
  wire _28297_;
  wire _28298_;
  wire _28299_;
  wire _28300_;
  wire _28301_;
  wire _28302_;
  wire _28303_;
  wire _28304_;
  wire _28305_;
  wire _28306_;
  wire _28307_;
  wire _28308_;
  wire _28309_;
  wire _28310_;
  wire _28311_;
  wire _28312_;
  wire _28313_;
  wire _28314_;
  wire _28315_;
  wire _28316_;
  wire _28317_;
  wire _28318_;
  wire _28319_;
  wire _28320_;
  wire _28321_;
  wire _28322_;
  wire _28323_;
  wire _28324_;
  wire _28325_;
  wire _28326_;
  wire _28327_;
  wire _28328_;
  wire _28329_;
  wire _28330_;
  wire _28331_;
  wire _28332_;
  wire _28333_;
  wire _28334_;
  wire _28335_;
  wire _28336_;
  wire _28337_;
  wire _28338_;
  wire _28339_;
  wire _28340_;
  wire _28341_;
  wire _28342_;
  wire _28343_;
  wire _28344_;
  wire _28345_;
  wire _28346_;
  wire _28347_;
  wire _28348_;
  wire _28349_;
  wire _28350_;
  wire _28351_;
  wire _28352_;
  wire _28353_;
  wire _28354_;
  wire _28355_;
  wire _28356_;
  wire _28357_;
  wire _28358_;
  wire _28359_;
  wire _28360_;
  wire _28361_;
  wire _28362_;
  wire _28363_;
  wire _28364_;
  wire _28365_;
  wire _28366_;
  wire _28367_;
  wire _28368_;
  wire _28369_;
  wire _28370_;
  wire _28371_;
  wire _28372_;
  wire _28373_;
  wire _28374_;
  wire _28375_;
  wire _28376_;
  wire _28377_;
  wire _28378_;
  wire _28379_;
  wire _28380_;
  wire _28381_;
  wire _28382_;
  wire _28383_;
  wire _28384_;
  wire _28385_;
  wire _28386_;
  wire _28387_;
  wire _28388_;
  wire _28389_;
  wire _28390_;
  wire _28391_;
  wire _28392_;
  wire _28393_;
  wire _28394_;
  wire _28395_;
  wire _28396_;
  wire _28397_;
  wire _28398_;
  wire _28399_;
  wire _28400_;
  wire _28401_;
  wire _28402_;
  wire _28403_;
  wire _28404_;
  wire _28405_;
  wire _28406_;
  wire _28407_;
  wire _28408_;
  wire _28409_;
  wire _28410_;
  wire _28411_;
  wire _28412_;
  wire _28413_;
  wire _28414_;
  wire _28415_;
  wire _28416_;
  wire _28417_;
  wire _28418_;
  wire _28419_;
  wire _28420_;
  wire _28421_;
  wire _28422_;
  wire _28423_;
  wire _28424_;
  wire _28425_;
  wire _28426_;
  wire _28427_;
  wire _28428_;
  wire _28429_;
  wire _28430_;
  wire _28431_;
  wire _28432_;
  wire _28433_;
  wire _28434_;
  wire _28435_;
  wire _28436_;
  wire _28437_;
  wire _28438_;
  wire _28439_;
  wire _28440_;
  wire _28441_;
  wire _28442_;
  wire _28443_;
  wire _28444_;
  wire _28445_;
  wire _28446_;
  wire _28447_;
  wire _28448_;
  wire _28449_;
  wire _28450_;
  wire _28451_;
  wire _28452_;
  wire _28453_;
  wire _28454_;
  wire _28455_;
  wire _28456_;
  wire _28457_;
  wire _28458_;
  wire _28459_;
  wire _28460_;
  wire _28461_;
  wire _28462_;
  wire _28463_;
  wire _28464_;
  wire _28465_;
  wire _28466_;
  wire _28467_;
  wire _28468_;
  wire _28469_;
  wire _28470_;
  wire _28471_;
  wire _28472_;
  wire _28473_;
  wire _28474_;
  wire _28475_;
  wire _28476_;
  wire _28477_;
  wire _28478_;
  wire _28479_;
  wire _28480_;
  wire _28481_;
  wire _28482_;
  wire _28483_;
  wire _28484_;
  wire _28485_;
  wire _28486_;
  wire _28487_;
  wire _28488_;
  wire _28489_;
  wire _28490_;
  wire _28491_;
  wire _28492_;
  wire _28493_;
  wire _28494_;
  wire _28495_;
  wire _28496_;
  wire _28497_;
  wire _28498_;
  wire _28499_;
  wire _28500_;
  wire _28501_;
  wire _28502_;
  wire _28503_;
  wire _28504_;
  wire _28505_;
  wire _28506_;
  wire _28507_;
  wire _28508_;
  wire _28509_;
  wire _28510_;
  wire _28511_;
  wire _28512_;
  wire _28513_;
  wire _28514_;
  wire _28515_;
  wire _28516_;
  wire _28517_;
  wire _28518_;
  wire _28519_;
  wire _28520_;
  wire _28521_;
  wire _28522_;
  wire _28523_;
  wire _28524_;
  wire _28525_;
  wire _28526_;
  wire _28527_;
  wire _28528_;
  wire _28529_;
  wire _28530_;
  wire _28531_;
  wire _28532_;
  wire _28533_;
  wire _28534_;
  wire _28535_;
  wire _28536_;
  wire _28537_;
  wire _28538_;
  wire _28539_;
  wire _28540_;
  wire _28541_;
  wire _28542_;
  wire _28543_;
  wire _28544_;
  wire _28545_;
  wire _28546_;
  wire _28547_;
  wire _28548_;
  wire _28549_;
  wire _28550_;
  wire _28551_;
  wire _28552_;
  wire _28553_;
  wire _28554_;
  wire _28555_;
  wire _28556_;
  wire _28557_;
  wire _28558_;
  wire _28559_;
  wire _28560_;
  wire _28561_;
  wire _28562_;
  wire _28563_;
  wire _28564_;
  wire _28565_;
  wire _28566_;
  wire _28567_;
  wire _28568_;
  wire _28569_;
  wire _28570_;
  wire _28571_;
  wire _28572_;
  wire _28573_;
  wire _28574_;
  wire _28575_;
  wire _28576_;
  wire _28577_;
  wire _28578_;
  wire _28579_;
  wire _28580_;
  wire _28581_;
  wire _28582_;
  wire _28583_;
  wire _28584_;
  wire _28585_;
  wire _28586_;
  wire _28587_;
  wire _28588_;
  wire _28589_;
  wire _28590_;
  wire _28591_;
  wire _28592_;
  wire _28593_;
  wire _28594_;
  wire _28595_;
  wire _28596_;
  wire _28597_;
  wire _28598_;
  wire _28599_;
  wire _28600_;
  wire _28601_;
  wire _28602_;
  wire _28603_;
  wire _28604_;
  wire _28605_;
  wire _28606_;
  wire _28607_;
  wire _28608_;
  wire _28609_;
  wire _28610_;
  wire _28611_;
  wire _28612_;
  wire _28613_;
  wire _28614_;
  wire _28615_;
  wire _28616_;
  wire _28617_;
  wire _28618_;
  wire _28619_;
  wire _28620_;
  wire _28621_;
  wire _28622_;
  wire _28623_;
  wire _28624_;
  wire _28625_;
  wire _28626_;
  wire _28627_;
  wire _28628_;
  wire _28629_;
  wire _28630_;
  wire _28631_;
  wire _28632_;
  wire _28633_;
  wire _28634_;
  wire _28635_;
  wire _28636_;
  wire _28637_;
  wire _28638_;
  wire _28639_;
  wire _28640_;
  wire _28641_;
  wire _28642_;
  wire _28643_;
  wire _28644_;
  wire _28645_;
  wire _28646_;
  wire _28647_;
  wire _28648_;
  wire _28649_;
  wire _28650_;
  wire _28651_;
  wire _28652_;
  wire _28653_;
  wire _28654_;
  wire _28655_;
  wire _28656_;
  wire _28657_;
  wire _28658_;
  wire _28659_;
  wire _28660_;
  wire _28661_;
  wire _28662_;
  wire _28663_;
  wire _28664_;
  wire _28665_;
  wire _28666_;
  wire _28667_;
  wire _28668_;
  wire _28669_;
  wire _28670_;
  wire _28671_;
  wire _28672_;
  wire _28673_;
  wire _28674_;
  wire _28675_;
  wire _28676_;
  wire _28677_;
  wire _28678_;
  wire _28679_;
  wire _28680_;
  wire _28681_;
  wire _28682_;
  wire _28683_;
  wire _28684_;
  wire _28685_;
  wire _28686_;
  wire _28687_;
  wire _28688_;
  wire _28689_;
  wire _28690_;
  wire _28691_;
  wire _28692_;
  wire _28693_;
  wire _28694_;
  wire _28695_;
  wire _28696_;
  wire _28697_;
  wire _28698_;
  wire _28699_;
  wire _28700_;
  wire _28701_;
  wire _28702_;
  wire _28703_;
  wire _28704_;
  wire _28705_;
  wire _28706_;
  wire _28707_;
  wire _28708_;
  wire _28709_;
  wire _28710_;
  wire _28711_;
  wire _28712_;
  wire _28713_;
  wire _28714_;
  wire _28715_;
  wire _28716_;
  wire _28717_;
  wire _28718_;
  wire _28719_;
  wire _28720_;
  wire _28721_;
  wire _28722_;
  wire _28723_;
  wire _28724_;
  wire _28725_;
  wire _28726_;
  wire _28727_;
  wire _28728_;
  wire _28729_;
  wire _28730_;
  wire _28731_;
  wire _28732_;
  wire _28733_;
  wire _28734_;
  wire _28735_;
  wire _28736_;
  wire _28737_;
  wire _28738_;
  wire _28739_;
  wire _28740_;
  wire _28741_;
  wire _28742_;
  wire _28743_;
  wire _28744_;
  wire _28745_;
  wire _28746_;
  wire _28747_;
  wire _28748_;
  wire _28749_;
  wire _28750_;
  wire _28751_;
  wire _28752_;
  wire _28753_;
  wire _28754_;
  wire _28755_;
  wire _28756_;
  wire _28757_;
  wire _28758_;
  wire _28759_;
  wire _28760_;
  wire _28761_;
  wire _28762_;
  wire _28763_;
  wire _28764_;
  wire _28765_;
  wire _28766_;
  wire _28767_;
  wire _28768_;
  wire _28769_;
  wire _28770_;
  wire _28771_;
  wire _28772_;
  wire _28773_;
  wire _28774_;
  wire _28775_;
  wire _28776_;
  wire _28777_;
  wire _28778_;
  wire _28779_;
  wire _28780_;
  wire _28781_;
  wire _28782_;
  wire _28783_;
  wire _28784_;
  wire _28785_;
  wire _28786_;
  wire _28787_;
  wire _28788_;
  wire _28789_;
  wire _28790_;
  wire _28791_;
  wire _28792_;
  wire _28793_;
  wire _28794_;
  wire _28795_;
  wire _28796_;
  wire _28797_;
  wire _28798_;
  wire _28799_;
  wire _28800_;
  wire _28801_;
  wire _28802_;
  wire _28803_;
  wire _28804_;
  wire _28805_;
  wire _28806_;
  wire _28807_;
  wire _28808_;
  wire _28809_;
  wire _28810_;
  wire _28811_;
  wire _28812_;
  wire _28813_;
  wire _28814_;
  wire _28815_;
  wire _28816_;
  wire _28817_;
  wire _28818_;
  wire _28819_;
  wire _28820_;
  wire _28821_;
  wire _28822_;
  wire _28823_;
  wire _28824_;
  wire _28825_;
  wire _28826_;
  wire _28827_;
  wire _28828_;
  wire _28829_;
  wire _28830_;
  wire _28831_;
  wire _28832_;
  wire _28833_;
  wire _28834_;
  wire _28835_;
  wire _28836_;
  wire _28837_;
  wire _28838_;
  wire _28839_;
  wire _28840_;
  wire _28841_;
  wire _28842_;
  wire _28843_;
  wire _28844_;
  wire _28845_;
  wire _28846_;
  wire _28847_;
  wire _28848_;
  wire _28849_;
  wire _28850_;
  wire _28851_;
  wire _28852_;
  wire _28853_;
  wire _28854_;
  wire _28855_;
  wire _28856_;
  wire _28857_;
  wire _28858_;
  wire _28859_;
  wire _28860_;
  wire _28861_;
  wire _28862_;
  wire _28863_;
  wire _28864_;
  wire _28865_;
  wire _28866_;
  wire _28867_;
  wire _28868_;
  wire _28869_;
  wire _28870_;
  wire _28871_;
  wire _28872_;
  wire _28873_;
  wire _28874_;
  wire _28875_;
  wire _28876_;
  wire _28877_;
  wire _28878_;
  wire _28879_;
  wire _28880_;
  wire _28881_;
  wire _28882_;
  wire _28883_;
  wire _28884_;
  wire _28885_;
  wire _28886_;
  wire _28887_;
  wire _28888_;
  wire _28889_;
  wire _28890_;
  wire _28891_;
  wire _28892_;
  wire _28893_;
  wire _28894_;
  wire _28895_;
  wire _28896_;
  wire _28897_;
  wire _28898_;
  wire _28899_;
  wire _28900_;
  wire _28901_;
  wire _28902_;
  wire _28903_;
  wire _28904_;
  wire _28905_;
  wire _28906_;
  wire _28907_;
  wire _28908_;
  wire _28909_;
  wire _28910_;
  wire _28911_;
  wire _28912_;
  wire _28913_;
  wire _28914_;
  wire _28915_;
  wire _28916_;
  wire _28917_;
  wire _28918_;
  wire _28919_;
  wire _28920_;
  wire _28921_;
  wire _28922_;
  wire _28923_;
  wire _28924_;
  wire _28925_;
  wire _28926_;
  wire _28927_;
  wire _28928_;
  wire _28929_;
  wire _28930_;
  wire _28931_;
  wire _28932_;
  wire _28933_;
  wire _28934_;
  wire _28935_;
  wire _28936_;
  wire _28937_;
  wire _28938_;
  wire _28939_;
  wire _28940_;
  wire _28941_;
  wire _28942_;
  wire _28943_;
  wire _28944_;
  wire _28945_;
  wire _28946_;
  wire _28947_;
  wire _28948_;
  wire _28949_;
  wire _28950_;
  wire _28951_;
  wire _28952_;
  wire _28953_;
  wire _28954_;
  wire _28955_;
  wire _28956_;
  wire _28957_;
  wire _28958_;
  wire _28959_;
  wire _28960_;
  wire _28961_;
  wire _28962_;
  wire _28963_;
  wire _28964_;
  wire _28965_;
  wire _28966_;
  wire _28967_;
  wire _28968_;
  wire _28969_;
  wire _28970_;
  wire _28971_;
  wire _28972_;
  wire _28973_;
  wire _28974_;
  wire _28975_;
  wire _28976_;
  wire _28977_;
  wire _28978_;
  wire _28979_;
  wire _28980_;
  wire _28981_;
  wire _28982_;
  wire _28983_;
  wire _28984_;
  wire _28985_;
  wire _28986_;
  wire _28987_;
  wire _28988_;
  wire _28989_;
  wire _28990_;
  wire _28991_;
  wire _28992_;
  wire _28993_;
  wire _28994_;
  wire _28995_;
  wire _28996_;
  wire _28997_;
  wire _28998_;
  wire _28999_;
  wire _29000_;
  wire _29001_;
  wire _29002_;
  wire _29003_;
  wire _29004_;
  wire _29005_;
  wire _29006_;
  wire _29007_;
  wire _29008_;
  wire _29009_;
  wire _29010_;
  wire _29011_;
  wire _29012_;
  wire _29013_;
  wire _29014_;
  wire _29015_;
  wire _29016_;
  wire _29017_;
  wire _29018_;
  wire _29019_;
  wire _29020_;
  wire _29021_;
  wire _29022_;
  wire _29023_;
  wire _29024_;
  wire _29025_;
  wire _29026_;
  wire _29027_;
  wire _29028_;
  wire _29029_;
  wire _29030_;
  wire _29031_;
  wire _29032_;
  wire _29033_;
  wire _29034_;
  wire _29035_;
  wire _29036_;
  wire _29037_;
  wire _29038_;
  wire _29039_;
  wire _29040_;
  wire _29041_;
  wire _29042_;
  wire _29043_;
  wire _29044_;
  wire _29045_;
  wire _29046_;
  wire _29047_;
  wire _29048_;
  wire _29049_;
  wire _29050_;
  wire _29051_;
  wire _29052_;
  wire _29053_;
  wire _29054_;
  wire _29055_;
  wire _29056_;
  wire _29057_;
  wire _29058_;
  wire _29059_;
  wire _29060_;
  wire _29061_;
  wire _29062_;
  wire _29063_;
  wire _29064_;
  wire _29065_;
  wire _29066_;
  wire _29067_;
  wire _29068_;
  wire _29069_;
  wire _29070_;
  wire _29071_;
  wire _29072_;
  wire _29073_;
  wire _29074_;
  wire _29075_;
  wire _29076_;
  wire _29077_;
  wire _29078_;
  wire _29079_;
  wire _29080_;
  wire _29081_;
  wire _29082_;
  wire _29083_;
  wire _29084_;
  wire _29085_;
  wire _29086_;
  wire _29087_;
  wire _29088_;
  wire _29089_;
  wire _29090_;
  wire _29091_;
  wire _29092_;
  wire _29093_;
  wire _29094_;
  wire _29095_;
  wire _29096_;
  wire _29097_;
  wire _29098_;
  wire _29099_;
  wire _29100_;
  wire _29101_;
  wire _29102_;
  wire _29103_;
  wire _29104_;
  wire _29105_;
  wire _29106_;
  wire _29107_;
  wire _29108_;
  wire _29109_;
  wire _29110_;
  wire _29111_;
  wire _29112_;
  wire _29113_;
  wire _29114_;
  wire _29115_;
  wire _29116_;
  wire _29117_;
  wire _29118_;
  wire _29119_;
  wire _29120_;
  wire _29121_;
  wire _29122_;
  wire _29123_;
  wire _29124_;
  wire _29125_;
  wire _29126_;
  wire _29127_;
  wire _29128_;
  wire _29129_;
  wire _29130_;
  wire _29131_;
  wire _29132_;
  wire _29133_;
  wire _29134_;
  wire _29135_;
  wire _29136_;
  wire _29137_;
  wire _29138_;
  wire _29139_;
  wire _29140_;
  wire _29141_;
  wire _29142_;
  wire _29143_;
  wire _29144_;
  wire [127:0] _29145_;
  wire [1:0] _29146_;
  wire [63:0] _29147_;
  wire [63:0] _29148_;
  wire [31:0] _29149_;
  wire [31:0] _29150_;
  wire [31:0] _29151_;
  wire [31:0] alu_out;
  wire [31:0] alu_out_q;
  input clk;
  wire clk;
  wire compressed_instr;
  wire [63:0] count_cycle;
  wire [63:0] count_instr;
  wire [7:0] cpu_state;
  wire [31:0] \cpuregs[0] ;
  wire [31:0] \cpuregs[10] ;
  wire [31:0] \cpuregs[11] ;
  wire [31:0] \cpuregs[12] ;
  wire [31:0] \cpuregs[13] ;
  wire [31:0] \cpuregs[14] ;
  wire [31:0] \cpuregs[15] ;
  wire [31:0] \cpuregs[16] ;
  wire [31:0] \cpuregs[17] ;
  wire [31:0] \cpuregs[18] ;
  wire [31:0] \cpuregs[19] ;
  wire [31:0] \cpuregs[1] ;
  wire [31:0] \cpuregs[20] ;
  wire [31:0] \cpuregs[21] ;
  wire [31:0] \cpuregs[22] ;
  wire [31:0] \cpuregs[23] ;
  wire [31:0] \cpuregs[24] ;
  wire [31:0] \cpuregs[25] ;
  wire [31:0] \cpuregs[26] ;
  wire [31:0] \cpuregs[27] ;
  wire [31:0] \cpuregs[28] ;
  wire [31:0] \cpuregs[29] ;
  wire [31:0] \cpuregs[2] ;
  wire [31:0] \cpuregs[30] ;
  wire [31:0] \cpuregs[31] ;
  wire [31:0] \cpuregs[3] ;
  wire [31:0] \cpuregs[4] ;
  wire [31:0] \cpuregs[5] ;
  wire [31:0] \cpuregs[6] ;
  wire [31:0] \cpuregs[7] ;
  wire [31:0] \cpuregs[8] ;
  wire [31:0] \cpuregs[9] ;
  wire [31:0] current_pc;
  wire [31:0] dbg_mem_addr;
  wire dbg_mem_instr;
  wire [31:0] dbg_mem_rdata;
  wire dbg_mem_ready;
  wire dbg_mem_valid;
  wire [31:0] dbg_mem_wdata;
  wire [3:0] dbg_mem_wstrb;
  wire [31:0] decoded_imm;
  wire [31:0] decoded_imm_j;
  wire [4:0] decoded_rd;
  wire [4:0] decoded_rs;
  wire [4:0] decoded_rs1;
  wire [4:0] decoded_rs2;
  wire decoder_pseudo_trigger;
  wire decoder_trigger;
  wire do_waitirq;
  output [31:0] eoi;
  wire [31:0] eoi;
  wire instr_add;
  wire instr_addi;
  wire instr_and;
  wire instr_andi;
  wire instr_auipc;
  wire instr_beq;
  wire instr_bge;
  wire instr_bgeu;
  wire instr_blt;
  wire instr_bltu;
  wire instr_bne;
  wire instr_fence;
  wire instr_getq;
  wire instr_jal;
  wire instr_jalr;
  wire instr_lb;
  wire instr_lbu;
  wire instr_lh;
  wire instr_lhu;
  wire instr_lui;
  wire instr_lw;
  wire instr_maskirq;
  wire instr_or;
  wire instr_ori;
  wire instr_rdcycle;
  wire instr_rdcycleh;
  wire instr_rdinstr;
  wire instr_rdinstrh;
  wire instr_retirq;
  wire instr_sb;
  wire instr_setq;
  wire instr_sh;
  wire instr_sll;
  wire instr_slli;
  wire instr_slt;
  wire instr_slti;
  wire instr_sltiu;
  wire instr_sltu;
  wire instr_sra;
  wire instr_srai;
  wire instr_srl;
  wire instr_srli;
  wire instr_sub;
  wire instr_sw;
  wire instr_timer;
  wire instr_waitirq;
  wire instr_xor;
  wire instr_xori;
  input [31:0] irq;
  wire [31:0] irq;
  wire [31:0] irq_mask;
  wire [31:0] irq_pending;
  wire is_alu_reg_imm;
  wire is_alu_reg_reg;
  wire is_beq_bne_blt_bge_bltu_bgeu;
  wire is_compare;
  wire is_jalr_addi_slti_sltiu_xori_ori_andi;
  wire is_lb_lh_lw_lbu_lhu;
  wire is_lbu_lhu_lw;
  wire is_lui_auipc_jal;
  wire is_lui_auipc_jal_jalr_addi_add_sub;
  wire is_sb_sh_sw;
  wire is_sll_srl_sra;
  wire is_slli_srli_srai;
  wire is_slti_blt_slt;
  wire is_sltiu_bltu_sltu;
  wire latched_branch;
  wire latched_compr;
  wire latched_is_lb;
  wire latched_is_lh;
  wire latched_is_lu;
  wire [4:0] latched_rd;
  wire latched_stalu;
  wire latched_store;
  output [31:0] mem_addr;
  wire [31:0] mem_addr;
  wire mem_do_prefetch;
  wire mem_do_rdata;
  wire mem_do_rinst;
  wire mem_do_wdata;
  output mem_instr;
  wire mem_instr;
  output [31:0] mem_la_addr;
  wire [31:0] mem_la_addr;
  wire mem_la_firstword;
  wire mem_la_firstword_reg;
  wire mem_la_firstword_xfer;
  output mem_la_read;
  wire mem_la_read;
  wire mem_la_secondword;
  wire mem_la_use_prefetched_high_word;
  output [31:0] mem_la_wdata;
  wire [31:0] mem_la_wdata;
  output mem_la_write;
  wire mem_la_write;
  output [3:0] mem_la_wstrb;
  wire [3:0] mem_la_wstrb;
  input [31:0] mem_rdata;
  wire [31:0] mem_rdata;
  wire [31:0] mem_rdata_q;
  input mem_ready;
  wire mem_ready;
  wire [1:0] mem_state;
  output mem_valid;
  wire mem_valid;
  output [31:0] mem_wdata;
  wire [31:0] mem_wdata;
  wire [1:0] mem_wordsize;
  output [3:0] mem_wstrb;
  wire [3:0] mem_wstrb;
  wire [31:0] next_irq_pending;
  wire [31:0] pcpi_div_rd;
  wire pcpi_div_ready;
  wire pcpi_div_wait;
  wire pcpi_div_wr;
  output [31:0] pcpi_insn;
  wire [31:0] pcpi_insn;
  wire [31:0] pcpi_int_rd;
  wire pcpi_int_ready;
  wire pcpi_int_wait;
  wire pcpi_int_wr;
  wire [31:0] pcpi_mul_rd;
  wire pcpi_mul_ready;
  wire pcpi_mul_wait;
  wire pcpi_mul_wr;
  input [31:0] pcpi_rd;
  wire [31:0] pcpi_rd;
  input pcpi_ready;
  wire pcpi_ready;
  output [31:0] pcpi_rs1;
  wire [31:0] pcpi_rs1;
  output [31:0] pcpi_rs2;
  wire [31:0] pcpi_rs2;
  wire pcpi_timeout;
  output pcpi_valid;
  wire pcpi_valid;
  input pcpi_wait;
  wire pcpi_wait;
  input pcpi_wr;
  wire pcpi_wr;
  wire [31:0] reg_next_pc;
  wire [31:0] reg_op1;
  wire [31:0] reg_op2;
  wire [31:0] reg_out;
  wire [31:0] reg_pc;
  wire [4:0] reg_sh;
  input resetn;
  wire resetn;
  wire [31:0] timer;
  output [35:0] trace_data;
  wire [35:0] trace_data;
  output trace_valid;
  wire trace_valid;
  output trap;
  wire trap;
  INV_X1 _29152_ (
    .A(reg_next_pc[0]),
    .ZN(_21037_)
  );
  INV_X1 _29153_ (
    .A(mem_do_wdata),
    .ZN(_21038_)
  );
  INV_X1 _29154_ (
    .A(is_beq_bne_blt_bge_bltu_bgeu),
    .ZN(_21039_)
  );
  INV_X1 _29155_ (
    .A(instr_fence),
    .ZN(_21040_)
  );
  INV_X1 _29156_ (
    .A(instr_and),
    .ZN(_21041_)
  );
  INV_X1 _29157_ (
    .A(instr_or),
    .ZN(_21042_)
  );
  INV_X1 _29158_ (
    .A(instr_sra),
    .ZN(_21043_)
  );
  INV_X1 _29159_ (
    .A(instr_srl),
    .ZN(_21044_)
  );
  INV_X1 _29160_ (
    .A(instr_xor),
    .ZN(_21045_)
  );
  INV_X1 _29161_ (
    .A(instr_sltu),
    .ZN(_21046_)
  );
  INV_X1 _29162_ (
    .A(instr_slt),
    .ZN(_21047_)
  );
  INV_X1 _29163_ (
    .A(instr_sll),
    .ZN(_21048_)
  );
  INV_X1 _29164_ (
    .A(instr_sub),
    .ZN(_21049_)
  );
  INV_X1 _29165_ (
    .A(instr_add),
    .ZN(_21050_)
  );
  INV_X1 _29166_ (
    .A(instr_andi),
    .ZN(_21051_)
  );
  INV_X1 _29167_ (
    .A(instr_ori),
    .ZN(_21052_)
  );
  INV_X1 _29168_ (
    .A(instr_xori),
    .ZN(_21053_)
  );
  INV_X1 _29169_ (
    .A(instr_sltiu),
    .ZN(_21054_)
  );
  INV_X1 _29170_ (
    .A(instr_slti),
    .ZN(_21055_)
  );
  INV_X1 _29171_ (
    .A(instr_addi),
    .ZN(_21056_)
  );
  INV_X1 _29172_ (
    .A(instr_bgeu),
    .ZN(_21057_)
  );
  INV_X1 _29173_ (
    .A(instr_bltu),
    .ZN(_21058_)
  );
  INV_X1 _29174_ (
    .A(instr_bge),
    .ZN(_21059_)
  );
  INV_X1 _29175_ (
    .A(instr_blt),
    .ZN(_21060_)
  );
  INV_X1 _29176_ (
    .A(instr_bne),
    .ZN(_21061_)
  );
  INV_X1 _29177_ (
    .A(instr_beq),
    .ZN(_21062_)
  );
  INV_X1 _29178_ (
    .A(latched_is_lb),
    .ZN(_21063_)
  );
  INV_X1 _29179_ (
    .A(latched_is_lh),
    .ZN(_21064_)
  );
  INV_X1 _29180_ (
    .A(latched_is_lu),
    .ZN(_21065_)
  );
  INV_X1 _29181_ (
    .A(latched_branch),
    .ZN(_21066_)
  );
  INV_X1 _29182_ (
    .A(latched_stalu),
    .ZN(_21067_)
  );
  INV_X1 _29183_ (
    .A(latched_store),
    .ZN(_21068_)
  );
  INV_X1 _29184_ (
    .A(mem_do_rdata),
    .ZN(_21069_)
  );
  INV_X1 _29185_ (
    .A(mem_do_rinst),
    .ZN(_21070_)
  );
  INV_X1 _29186_ (
    .A(mem_do_prefetch),
    .ZN(_21071_)
  );
  INV_X1 _29187_ (
    .A(_00028_),
    .ZN(_21072_)
  );
  INV_X1 _29188_ (
    .A(reg_pc[31]),
    .ZN(_21073_)
  );
  INV_X1 _29189_ (
    .A(reg_pc[30]),
    .ZN(_21074_)
  );
  INV_X1 _29190_ (
    .A(reg_pc[29]),
    .ZN(_21075_)
  );
  INV_X1 _29191_ (
    .A(reg_pc[28]),
    .ZN(_21076_)
  );
  INV_X1 _29192_ (
    .A(reg_pc[27]),
    .ZN(_21077_)
  );
  INV_X1 _29193_ (
    .A(reg_pc[26]),
    .ZN(_21078_)
  );
  INV_X1 _29194_ (
    .A(reg_pc[25]),
    .ZN(_21079_)
  );
  INV_X1 _29195_ (
    .A(reg_pc[24]),
    .ZN(_21080_)
  );
  INV_X1 _29196_ (
    .A(reg_pc[23]),
    .ZN(_21081_)
  );
  INV_X1 _29197_ (
    .A(reg_pc[22]),
    .ZN(_21082_)
  );
  INV_X1 _29198_ (
    .A(reg_pc[21]),
    .ZN(_21083_)
  );
  INV_X1 _29199_ (
    .A(reg_pc[20]),
    .ZN(_21084_)
  );
  INV_X1 _29200_ (
    .A(reg_pc[19]),
    .ZN(_21085_)
  );
  INV_X1 _29201_ (
    .A(reg_pc[18]),
    .ZN(_21086_)
  );
  INV_X1 _29202_ (
    .A(reg_pc[17]),
    .ZN(_21087_)
  );
  INV_X1 _29203_ (
    .A(reg_pc[16]),
    .ZN(_21088_)
  );
  INV_X1 _29204_ (
    .A(reg_pc[15]),
    .ZN(_21089_)
  );
  INV_X1 _29205_ (
    .A(reg_pc[14]),
    .ZN(_21090_)
  );
  INV_X1 _29206_ (
    .A(reg_pc[13]),
    .ZN(_21091_)
  );
  INV_X1 _29207_ (
    .A(reg_pc[12]),
    .ZN(_21092_)
  );
  INV_X1 _29208_ (
    .A(reg_pc[11]),
    .ZN(_21093_)
  );
  INV_X1 _29209_ (
    .A(reg_pc[10]),
    .ZN(_21094_)
  );
  INV_X1 _29210_ (
    .A(reg_pc[9]),
    .ZN(_21095_)
  );
  INV_X1 _29211_ (
    .A(reg_pc[8]),
    .ZN(_21096_)
  );
  INV_X1 _29212_ (
    .A(reg_pc[7]),
    .ZN(_21097_)
  );
  INV_X1 _29213_ (
    .A(reg_pc[6]),
    .ZN(_21098_)
  );
  INV_X1 _29214_ (
    .A(reg_pc[5]),
    .ZN(_21099_)
  );
  INV_X1 _29215_ (
    .A(reg_pc[4]),
    .ZN(_21100_)
  );
  INV_X1 _29216_ (
    .A(reg_pc[3]),
    .ZN(_21101_)
  );
  INV_X1 _29217_ (
    .A(reg_pc[2]),
    .ZN(_21102_)
  );
  INV_X1 _29218_ (
    .A(reg_pc[1]),
    .ZN(_21103_)
  );
  INV_X1 _29219_ (
    .A(count_instr[63]),
    .ZN(_21104_)
  );
  INV_X1 _29220_ (
    .A(count_instr[62]),
    .ZN(_21105_)
  );
  INV_X1 _29221_ (
    .A(count_instr[61]),
    .ZN(_21106_)
  );
  INV_X1 _29222_ (
    .A(count_instr[60]),
    .ZN(_21107_)
  );
  INV_X1 _29223_ (
    .A(count_instr[59]),
    .ZN(_21108_)
  );
  INV_X1 _29224_ (
    .A(count_instr[58]),
    .ZN(_21109_)
  );
  INV_X1 _29225_ (
    .A(count_instr[57]),
    .ZN(_21110_)
  );
  INV_X1 _29226_ (
    .A(count_instr[56]),
    .ZN(_21111_)
  );
  INV_X1 _29227_ (
    .A(count_instr[55]),
    .ZN(_21112_)
  );
  INV_X1 _29228_ (
    .A(count_instr[54]),
    .ZN(_21113_)
  );
  INV_X1 _29229_ (
    .A(count_instr[53]),
    .ZN(_21114_)
  );
  INV_X1 _29230_ (
    .A(count_instr[52]),
    .ZN(_21115_)
  );
  INV_X1 _29231_ (
    .A(count_instr[51]),
    .ZN(_21116_)
  );
  INV_X1 _29232_ (
    .A(count_instr[50]),
    .ZN(_21117_)
  );
  INV_X1 _29233_ (
    .A(count_instr[49]),
    .ZN(_21118_)
  );
  INV_X1 _29234_ (
    .A(count_instr[48]),
    .ZN(_21119_)
  );
  INV_X1 _29235_ (
    .A(count_instr[47]),
    .ZN(_21120_)
  );
  INV_X1 _29236_ (
    .A(count_instr[46]),
    .ZN(_21121_)
  );
  INV_X1 _29237_ (
    .A(count_instr[45]),
    .ZN(_21122_)
  );
  INV_X1 _29238_ (
    .A(count_instr[44]),
    .ZN(_21123_)
  );
  INV_X1 _29239_ (
    .A(count_instr[43]),
    .ZN(_21124_)
  );
  INV_X1 _29240_ (
    .A(count_instr[42]),
    .ZN(_21125_)
  );
  INV_X1 _29241_ (
    .A(count_instr[41]),
    .ZN(_21126_)
  );
  INV_X1 _29242_ (
    .A(count_instr[40]),
    .ZN(_21127_)
  );
  INV_X1 _29243_ (
    .A(count_instr[39]),
    .ZN(_21128_)
  );
  INV_X1 _29244_ (
    .A(count_instr[38]),
    .ZN(_21129_)
  );
  INV_X1 _29245_ (
    .A(count_instr[37]),
    .ZN(_21130_)
  );
  INV_X1 _29246_ (
    .A(count_instr[36]),
    .ZN(_21131_)
  );
  INV_X1 _29247_ (
    .A(count_instr[35]),
    .ZN(_21132_)
  );
  INV_X1 _29248_ (
    .A(count_instr[34]),
    .ZN(_21133_)
  );
  INV_X1 _29249_ (
    .A(count_instr[33]),
    .ZN(_21134_)
  );
  INV_X1 _29250_ (
    .A(count_instr[32]),
    .ZN(_21135_)
  );
  INV_X1 _29251_ (
    .A(count_instr[31]),
    .ZN(_21136_)
  );
  INV_X1 _29252_ (
    .A(count_instr[30]),
    .ZN(_21137_)
  );
  INV_X1 _29253_ (
    .A(count_instr[29]),
    .ZN(_21138_)
  );
  INV_X1 _29254_ (
    .A(count_instr[28]),
    .ZN(_21139_)
  );
  INV_X1 _29255_ (
    .A(count_instr[27]),
    .ZN(_21140_)
  );
  INV_X1 _29256_ (
    .A(count_instr[26]),
    .ZN(_21141_)
  );
  INV_X1 _29257_ (
    .A(count_instr[25]),
    .ZN(_21142_)
  );
  INV_X1 _29258_ (
    .A(count_instr[24]),
    .ZN(_21143_)
  );
  INV_X1 _29259_ (
    .A(count_instr[23]),
    .ZN(_21144_)
  );
  INV_X1 _29260_ (
    .A(count_instr[22]),
    .ZN(_21145_)
  );
  INV_X1 _29261_ (
    .A(count_instr[21]),
    .ZN(_21146_)
  );
  INV_X1 _29262_ (
    .A(count_instr[20]),
    .ZN(_21147_)
  );
  INV_X1 _29263_ (
    .A(count_instr[19]),
    .ZN(_21148_)
  );
  INV_X1 _29264_ (
    .A(count_instr[18]),
    .ZN(_21149_)
  );
  INV_X1 _29265_ (
    .A(count_instr[17]),
    .ZN(_21150_)
  );
  INV_X1 _29266_ (
    .A(count_instr[16]),
    .ZN(_21151_)
  );
  INV_X1 _29267_ (
    .A(count_instr[15]),
    .ZN(_21152_)
  );
  INV_X1 _29268_ (
    .A(count_instr[14]),
    .ZN(_21153_)
  );
  INV_X1 _29269_ (
    .A(count_instr[13]),
    .ZN(_21154_)
  );
  INV_X1 _29270_ (
    .A(count_instr[12]),
    .ZN(_21155_)
  );
  INV_X1 _29271_ (
    .A(count_instr[11]),
    .ZN(_21156_)
  );
  INV_X1 _29272_ (
    .A(count_instr[10]),
    .ZN(_21157_)
  );
  INV_X1 _29273_ (
    .A(count_instr[9]),
    .ZN(_21158_)
  );
  INV_X1 _29274_ (
    .A(count_instr[8]),
    .ZN(_21159_)
  );
  INV_X1 _29275_ (
    .A(count_instr[7]),
    .ZN(_21160_)
  );
  INV_X1 _29276_ (
    .A(count_instr[6]),
    .ZN(_21161_)
  );
  INV_X1 _29277_ (
    .A(count_instr[5]),
    .ZN(_21162_)
  );
  INV_X1 _29278_ (
    .A(count_instr[4]),
    .ZN(_21163_)
  );
  INV_X1 _29279_ (
    .A(count_instr[3]),
    .ZN(_21164_)
  );
  INV_X1 _29280_ (
    .A(count_instr[2]),
    .ZN(_21165_)
  );
  INV_X1 _29281_ (
    .A(count_instr[1]),
    .ZN(_21166_)
  );
  INV_X1 _29282_ (
    .A(_29148_[0]),
    .ZN(_21167_)
  );
  INV_X1 _29283_ (
    .A(reg_op1[0]),
    .ZN(_21168_)
  );
  INV_X1 _29284_ (
    .A(reg_op1[2]),
    .ZN(_21169_)
  );
  INV_X1 _29285_ (
    .A(reg_op1[3]),
    .ZN(_21170_)
  );
  INV_X1 _29286_ (
    .A(reg_op1[4]),
    .ZN(_21171_)
  );
  INV_X1 _29287_ (
    .A(reg_op1[5]),
    .ZN(_21172_)
  );
  INV_X1 _29288_ (
    .A(reg_op1[6]),
    .ZN(_21173_)
  );
  INV_X1 _29289_ (
    .A(reg_op1[7]),
    .ZN(_21174_)
  );
  INV_X1 _29290_ (
    .A(reg_op1[8]),
    .ZN(_21175_)
  );
  INV_X1 _29291_ (
    .A(reg_op1[9]),
    .ZN(_21176_)
  );
  INV_X1 _29292_ (
    .A(reg_op1[10]),
    .ZN(_21177_)
  );
  INV_X1 _29293_ (
    .A(reg_op1[11]),
    .ZN(_21178_)
  );
  INV_X1 _29294_ (
    .A(reg_op1[12]),
    .ZN(_21179_)
  );
  INV_X1 _29295_ (
    .A(reg_op1[13]),
    .ZN(_21180_)
  );
  INV_X1 _29296_ (
    .A(reg_op1[14]),
    .ZN(_21181_)
  );
  INV_X1 _29297_ (
    .A(reg_op1[15]),
    .ZN(_21182_)
  );
  INV_X1 _29298_ (
    .A(reg_op1[16]),
    .ZN(_21183_)
  );
  INV_X1 _29299_ (
    .A(reg_op1[17]),
    .ZN(_21184_)
  );
  INV_X1 _29300_ (
    .A(reg_op1[18]),
    .ZN(_21185_)
  );
  INV_X1 _29301_ (
    .A(reg_op1[19]),
    .ZN(_21186_)
  );
  INV_X1 _29302_ (
    .A(reg_op1[20]),
    .ZN(_21187_)
  );
  INV_X1 _29303_ (
    .A(reg_op1[21]),
    .ZN(_21188_)
  );
  INV_X1 _29304_ (
    .A(reg_op1[22]),
    .ZN(_21189_)
  );
  INV_X1 _29305_ (
    .A(reg_op1[23]),
    .ZN(_21190_)
  );
  INV_X1 _29306_ (
    .A(reg_op1[24]),
    .ZN(_21191_)
  );
  INV_X1 _29307_ (
    .A(reg_op1[25]),
    .ZN(_21192_)
  );
  INV_X1 _29308_ (
    .A(reg_op1[26]),
    .ZN(_21193_)
  );
  INV_X1 _29309_ (
    .A(reg_op1[27]),
    .ZN(_21194_)
  );
  INV_X1 _29310_ (
    .A(reg_op1[28]),
    .ZN(_21195_)
  );
  INV_X1 _29311_ (
    .A(reg_op1[29]),
    .ZN(_21196_)
  );
  INV_X1 _29312_ (
    .A(reg_op1[30]),
    .ZN(_21197_)
  );
  INV_X1 _29313_ (
    .A(instr_sw),
    .ZN(_21198_)
  );
  INV_X1 _29314_ (
    .A(reg_op1[31]),
    .ZN(_21199_)
  );
  INV_X1 _29315_ (
    .A(reg_op2[0]),
    .ZN(_21200_)
  );
  INV_X1 _29316_ (
    .A(reg_op2[1]),
    .ZN(_21201_)
  );
  INV_X1 _29317_ (
    .A(reg_op2[2]),
    .ZN(_21202_)
  );
  INV_X1 _29318_ (
    .A(reg_op2[3]),
    .ZN(_21203_)
  );
  INV_X1 _29319_ (
    .A(reg_op2[4]),
    .ZN(_21204_)
  );
  INV_X1 _29320_ (
    .A(reg_op2[5]),
    .ZN(_21205_)
  );
  INV_X1 _29321_ (
    .A(reg_op2[6]),
    .ZN(_21206_)
  );
  INV_X1 _29322_ (
    .A(reg_op2[7]),
    .ZN(_21207_)
  );
  INV_X1 _29323_ (
    .A(reg_op2[8]),
    .ZN(_21208_)
  );
  INV_X1 _29324_ (
    .A(reg_op2[9]),
    .ZN(_21209_)
  );
  INV_X1 _29325_ (
    .A(reg_op2[10]),
    .ZN(_21210_)
  );
  INV_X1 _29326_ (
    .A(reg_op2[11]),
    .ZN(_21211_)
  );
  INV_X1 _29327_ (
    .A(reg_op2[12]),
    .ZN(_21212_)
  );
  INV_X1 _29328_ (
    .A(reg_op2[13]),
    .ZN(_21213_)
  );
  INV_X1 _29329_ (
    .A(reg_op2[14]),
    .ZN(_21214_)
  );
  INV_X1 _29330_ (
    .A(reg_op2[15]),
    .ZN(_21215_)
  );
  INV_X1 _29331_ (
    .A(reg_op2[16]),
    .ZN(_21216_)
  );
  INV_X1 _29332_ (
    .A(reg_op2[17]),
    .ZN(_21217_)
  );
  INV_X1 _29333_ (
    .A(reg_op2[18]),
    .ZN(_21218_)
  );
  INV_X1 _29334_ (
    .A(reg_op2[19]),
    .ZN(_21219_)
  );
  INV_X1 _29335_ (
    .A(reg_op2[20]),
    .ZN(_21220_)
  );
  INV_X1 _29336_ (
    .A(reg_op2[21]),
    .ZN(_21221_)
  );
  INV_X1 _29337_ (
    .A(reg_op2[22]),
    .ZN(_21222_)
  );
  INV_X1 _29338_ (
    .A(reg_op2[23]),
    .ZN(_21223_)
  );
  INV_X1 _29339_ (
    .A(reg_op2[24]),
    .ZN(_21224_)
  );
  INV_X1 _29340_ (
    .A(reg_op2[25]),
    .ZN(_21225_)
  );
  INV_X1 _29341_ (
    .A(reg_op2[26]),
    .ZN(_21226_)
  );
  INV_X1 _29342_ (
    .A(reg_op2[27]),
    .ZN(_21227_)
  );
  INV_X1 _29343_ (
    .A(reg_op2[28]),
    .ZN(_21228_)
  );
  INV_X1 _29344_ (
    .A(reg_op2[29]),
    .ZN(_21229_)
  );
  INV_X1 _29345_ (
    .A(reg_op2[30]),
    .ZN(_21230_)
  );
  INV_X1 _29346_ (
    .A(reg_op2[31]),
    .ZN(_21231_)
  );
  INV_X1 _29347_ (
    .A(mem_rdata_q[12]),
    .ZN(_21232_)
  );
  INV_X1 _29348_ (
    .A(mem_rdata_q[13]),
    .ZN(_21233_)
  );
  INV_X1 _29349_ (
    .A(mem_rdata_q[14]),
    .ZN(_21234_)
  );
  INV_X1 _29350_ (
    .A(mem_rdata_q[15]),
    .ZN(_21235_)
  );
  INV_X1 _29351_ (
    .A(mem_rdata_q[16]),
    .ZN(_21236_)
  );
  INV_X1 _29352_ (
    .A(mem_rdata_q[17]),
    .ZN(_21237_)
  );
  INV_X1 _29353_ (
    .A(mem_rdata_q[18]),
    .ZN(_21238_)
  );
  INV_X1 _29354_ (
    .A(mem_rdata_q[19]),
    .ZN(_21239_)
  );
  INV_X1 _29355_ (
    .A(mem_rdata_q[20]),
    .ZN(_21240_)
  );
  INV_X1 _29356_ (
    .A(mem_rdata_q[21]),
    .ZN(_21241_)
  );
  INV_X1 _29357_ (
    .A(mem_rdata_q[22]),
    .ZN(_21242_)
  );
  INV_X1 _29358_ (
    .A(mem_rdata_q[23]),
    .ZN(_21243_)
  );
  INV_X1 _29359_ (
    .A(mem_rdata_q[24]),
    .ZN(_21244_)
  );
  INV_X1 _29360_ (
    .A(mem_rdata_q[25]),
    .ZN(_21245_)
  );
  INV_X1 _29361_ (
    .A(mem_rdata_q[26]),
    .ZN(_21246_)
  );
  INV_X1 _29362_ (
    .A(mem_rdata_q[27]),
    .ZN(_21247_)
  );
  INV_X1 _29363_ (
    .A(mem_rdata_q[28]),
    .ZN(_21248_)
  );
  INV_X1 _29364_ (
    .A(mem_rdata_q[29]),
    .ZN(_21249_)
  );
  INV_X1 _29365_ (
    .A(mem_rdata_q[30]),
    .ZN(_21250_)
  );
  INV_X1 _29366_ (
    .A(mem_rdata_q[31]),
    .ZN(_21251_)
  );
  INV_X1 _29367_ (
    .A(mem_wordsize[0]),
    .ZN(_21252_)
  );
  INV_X1 _29368_ (
    .A(mem_wordsize[1]),
    .ZN(_21253_)
  );
  INV_X1 _29369_ (
    .A(latched_rd[0]),
    .ZN(_21254_)
  );
  INV_X1 _29370_ (
    .A(latched_rd[1]),
    .ZN(_21255_)
  );
  INV_X1 _29371_ (
    .A(latched_rd[2]),
    .ZN(_21256_)
  );
  INV_X1 _29372_ (
    .A(latched_rd[3]),
    .ZN(_21257_)
  );
  INV_X1 _29373_ (
    .A(latched_rd[4]),
    .ZN(_21258_)
  );
  INV_X1 _29374_ (
    .A(instr_lui),
    .ZN(_21259_)
  );
  INV_X1 _29375_ (
    .A(instr_auipc),
    .ZN(_21260_)
  );
  INV_X1 _29376_ (
    .A(instr_jal),
    .ZN(_21261_)
  );
  INV_X1 _29377_ (
    .A(instr_jalr),
    .ZN(_21262_)
  );
  INV_X1 _29378_ (
    .A(instr_lb),
    .ZN(_21263_)
  );
  INV_X1 _29379_ (
    .A(instr_lh),
    .ZN(_21264_)
  );
  INV_X1 _29380_ (
    .A(instr_lw),
    .ZN(_21265_)
  );
  INV_X1 _29381_ (
    .A(instr_lbu),
    .ZN(_21266_)
  );
  INV_X1 _29382_ (
    .A(instr_lhu),
    .ZN(_21267_)
  );
  INV_X1 _29383_ (
    .A(instr_sh),
    .ZN(_21268_)
  );
  INV_X1 _29384_ (
    .A(instr_sb),
    .ZN(_21269_)
  );
  INV_X1 _29385_ (
    .A(instr_slli),
    .ZN(_21270_)
  );
  INV_X1 _29386_ (
    .A(instr_srli),
    .ZN(_21271_)
  );
  INV_X1 _29387_ (
    .A(instr_srai),
    .ZN(_21272_)
  );
  INV_X1 _29388_ (
    .A(instr_rdcycle),
    .ZN(_21273_)
  );
  INV_X1 _29389_ (
    .A(instr_rdcycleh),
    .ZN(_21274_)
  );
  INV_X1 _29390_ (
    .A(instr_rdinstr),
    .ZN(_21275_)
  );
  INV_X1 _29391_ (
    .A(instr_rdinstrh),
    .ZN(_21276_)
  );
  INV_X1 _29392_ (
    .A(decoded_rd[0]),
    .ZN(_21277_)
  );
  INV_X1 _29393_ (
    .A(decoded_rd[1]),
    .ZN(_21278_)
  );
  INV_X1 _29394_ (
    .A(decoded_rd[2]),
    .ZN(_21279_)
  );
  INV_X1 _29395_ (
    .A(decoded_rd[3]),
    .ZN(_21280_)
  );
  INV_X1 _29396_ (
    .A(decoded_rd[4]),
    .ZN(_21281_)
  );
  INV_X1 _29397_ (
    .A(decoded_rs2[0]),
    .ZN(_21282_)
  );
  INV_X1 _29398_ (
    .A(decoded_rs2[1]),
    .ZN(_21283_)
  );
  INV_X1 _29399_ (
    .A(decoded_rs2[2]),
    .ZN(_21284_)
  );
  INV_X1 _29400_ (
    .A(decoded_rs2[3]),
    .ZN(_21285_)
  );
  INV_X1 _29401_ (
    .A(decoded_imm[0]),
    .ZN(_21286_)
  );
  INV_X1 _29402_ (
    .A(decoded_imm_j[10]),
    .ZN(_21287_)
  );
  INV_X1 _29403_ (
    .A(is_lb_lh_lw_lbu_lhu),
    .ZN(_21288_)
  );
  INV_X1 _29404_ (
    .A(is_slli_srli_srai),
    .ZN(_21289_)
  );
  INV_X1 _29405_ (
    .A(is_sb_sh_sw),
    .ZN(_21290_)
  );
  INV_X1 _29406_ (
    .A(is_sll_srl_sra),
    .ZN(_21291_)
  );
  INV_X1 _29407_ (
    .A(is_alu_reg_imm),
    .ZN(_21292_)
  );
  INV_X1 _29408_ (
    .A(is_jalr_addi_slti_sltiu_xori_ori_andi),
    .ZN(_21293_)
  );
  INV_X1 _29409_ (
    .A(mem_addr[2]),
    .ZN(_21294_)
  );
  INV_X1 _29410_ (
    .A(mem_addr[3]),
    .ZN(_21295_)
  );
  INV_X1 _29411_ (
    .A(mem_addr[4]),
    .ZN(_21296_)
  );
  INV_X1 _29412_ (
    .A(mem_addr[5]),
    .ZN(_21297_)
  );
  INV_X1 _29413_ (
    .A(mem_addr[6]),
    .ZN(_21298_)
  );
  INV_X1 _29414_ (
    .A(mem_addr[7]),
    .ZN(_21299_)
  );
  INV_X1 _29415_ (
    .A(mem_addr[8]),
    .ZN(_21300_)
  );
  INV_X1 _29416_ (
    .A(mem_addr[9]),
    .ZN(_21301_)
  );
  INV_X1 _29417_ (
    .A(mem_addr[10]),
    .ZN(_21302_)
  );
  INV_X1 _29418_ (
    .A(mem_addr[11]),
    .ZN(_21303_)
  );
  INV_X1 _29419_ (
    .A(mem_addr[12]),
    .ZN(_21304_)
  );
  INV_X1 _29420_ (
    .A(mem_addr[13]),
    .ZN(_21305_)
  );
  INV_X1 _29421_ (
    .A(mem_addr[14]),
    .ZN(_21306_)
  );
  INV_X1 _29422_ (
    .A(mem_addr[15]),
    .ZN(_21307_)
  );
  INV_X1 _29423_ (
    .A(mem_addr[16]),
    .ZN(_21308_)
  );
  INV_X1 _29424_ (
    .A(mem_addr[17]),
    .ZN(_21309_)
  );
  INV_X1 _29425_ (
    .A(mem_addr[18]),
    .ZN(_21310_)
  );
  INV_X1 _29426_ (
    .A(mem_addr[19]),
    .ZN(_21311_)
  );
  INV_X1 _29427_ (
    .A(mem_addr[20]),
    .ZN(_21312_)
  );
  INV_X1 _29428_ (
    .A(mem_addr[21]),
    .ZN(_21313_)
  );
  INV_X1 _29429_ (
    .A(mem_addr[22]),
    .ZN(_21314_)
  );
  INV_X1 _29430_ (
    .A(mem_addr[23]),
    .ZN(_21315_)
  );
  INV_X1 _29431_ (
    .A(mem_addr[24]),
    .ZN(_21316_)
  );
  INV_X1 _29432_ (
    .A(mem_addr[25]),
    .ZN(_21317_)
  );
  INV_X1 _29433_ (
    .A(mem_addr[26]),
    .ZN(_21318_)
  );
  INV_X1 _29434_ (
    .A(mem_addr[27]),
    .ZN(_21319_)
  );
  INV_X1 _29435_ (
    .A(mem_addr[28]),
    .ZN(_21320_)
  );
  INV_X1 _29436_ (
    .A(mem_addr[29]),
    .ZN(_21321_)
  );
  INV_X1 _29437_ (
    .A(mem_addr[30]),
    .ZN(_21322_)
  );
  INV_X1 _29438_ (
    .A(mem_addr[31]),
    .ZN(_21323_)
  );
  INV_X1 _29439_ (
    .A(mem_wdata[8]),
    .ZN(_21324_)
  );
  INV_X1 _29440_ (
    .A(mem_wdata[9]),
    .ZN(_21325_)
  );
  INV_X1 _29441_ (
    .A(mem_wdata[10]),
    .ZN(_21326_)
  );
  INV_X1 _29442_ (
    .A(mem_wdata[11]),
    .ZN(_21327_)
  );
  INV_X1 _29443_ (
    .A(mem_wdata[12]),
    .ZN(_21328_)
  );
  INV_X1 _29444_ (
    .A(mem_wdata[13]),
    .ZN(_21329_)
  );
  INV_X1 _29445_ (
    .A(mem_wdata[14]),
    .ZN(_21330_)
  );
  INV_X1 _29446_ (
    .A(mem_wdata[15]),
    .ZN(_21331_)
  );
  INV_X1 _29447_ (
    .A(mem_wdata[16]),
    .ZN(_21332_)
  );
  INV_X1 _29448_ (
    .A(mem_wdata[17]),
    .ZN(_21333_)
  );
  INV_X1 _29449_ (
    .A(mem_wdata[18]),
    .ZN(_21334_)
  );
  INV_X1 _29450_ (
    .A(mem_wdata[19]),
    .ZN(_21335_)
  );
  INV_X1 _29451_ (
    .A(mem_wdata[20]),
    .ZN(_21336_)
  );
  INV_X1 _29452_ (
    .A(mem_wdata[21]),
    .ZN(_21337_)
  );
  INV_X1 _29453_ (
    .A(mem_wdata[22]),
    .ZN(_21338_)
  );
  INV_X1 _29454_ (
    .A(mem_wdata[23]),
    .ZN(_21339_)
  );
  INV_X1 _29455_ (
    .A(mem_wdata[24]),
    .ZN(_21340_)
  );
  INV_X1 _29456_ (
    .A(mem_wdata[25]),
    .ZN(_21341_)
  );
  INV_X1 _29457_ (
    .A(mem_wdata[26]),
    .ZN(_21342_)
  );
  INV_X1 _29458_ (
    .A(mem_wdata[27]),
    .ZN(_21343_)
  );
  INV_X1 _29459_ (
    .A(mem_wdata[28]),
    .ZN(_21344_)
  );
  INV_X1 _29460_ (
    .A(mem_wdata[29]),
    .ZN(_21345_)
  );
  INV_X1 _29461_ (
    .A(mem_wdata[30]),
    .ZN(_21346_)
  );
  INV_X1 _29462_ (
    .A(mem_wdata[31]),
    .ZN(_21347_)
  );
  INV_X1 _29463_ (
    .A(mem_state[0]),
    .ZN(_21348_)
  );
  INV_X1 _29464_ (
    .A(mem_state[1]),
    .ZN(_21349_)
  );
  INV_X1 _29465_ (
    .A(mem_rdata_q[0]),
    .ZN(_21350_)
  );
  INV_X1 _29466_ (
    .A(mem_rdata[0]),
    .ZN(_21351_)
  );
  INV_X1 _29467_ (
    .A(mem_rdata_q[1]),
    .ZN(_21352_)
  );
  INV_X1 _29468_ (
    .A(mem_rdata[1]),
    .ZN(_21353_)
  );
  INV_X1 _29469_ (
    .A(mem_rdata_q[2]),
    .ZN(_21354_)
  );
  INV_X1 _29470_ (
    .A(mem_rdata[2]),
    .ZN(_21355_)
  );
  INV_X1 _29471_ (
    .A(mem_rdata_q[3]),
    .ZN(_21356_)
  );
  INV_X1 _29472_ (
    .A(mem_rdata_q[4]),
    .ZN(_21357_)
  );
  INV_X1 _29473_ (
    .A(mem_rdata_q[5]),
    .ZN(_21358_)
  );
  INV_X1 _29474_ (
    .A(mem_rdata_q[6]),
    .ZN(_21359_)
  );
  INV_X1 _29475_ (
    .A(\cpuregs[6] [31]),
    .ZN(_21360_)
  );
  INV_X1 _29476_ (
    .A(\cpuregs[2] [31]),
    .ZN(_21361_)
  );
  INV_X1 _29477_ (
    .A(\cpuregs[23] [31]),
    .ZN(_21362_)
  );
  INV_X1 _29478_ (
    .A(\cpuregs[22] [31]),
    .ZN(_21363_)
  );
  INV_X1 _29479_ (
    .A(\cpuregs[21] [31]),
    .ZN(_21364_)
  );
  INV_X1 _29480_ (
    .A(\cpuregs[20] [31]),
    .ZN(_21365_)
  );
  INV_X1 _29481_ (
    .A(\cpuregs[19] [31]),
    .ZN(_21366_)
  );
  INV_X1 _29482_ (
    .A(\cpuregs[18] [31]),
    .ZN(_21367_)
  );
  INV_X1 _29483_ (
    .A(\cpuregs[17] [31]),
    .ZN(_21368_)
  );
  INV_X1 _29484_ (
    .A(\cpuregs[16] [31]),
    .ZN(_21369_)
  );
  INV_X1 _29485_ (
    .A(\cpuregs[23] [0]),
    .ZN(_21370_)
  );
  INV_X1 _29486_ (
    .A(\cpuregs[23] [1]),
    .ZN(_21371_)
  );
  INV_X1 _29487_ (
    .A(\cpuregs[23] [2]),
    .ZN(_21372_)
  );
  INV_X1 _29488_ (
    .A(\cpuregs[23] [3]),
    .ZN(_21373_)
  );
  INV_X1 _29489_ (
    .A(\cpuregs[23] [4]),
    .ZN(_21374_)
  );
  INV_X1 _29490_ (
    .A(\cpuregs[23] [5]),
    .ZN(_21375_)
  );
  INV_X1 _29491_ (
    .A(\cpuregs[23] [7]),
    .ZN(_21376_)
  );
  INV_X1 _29492_ (
    .A(\cpuregs[23] [9]),
    .ZN(_21377_)
  );
  INV_X1 _29493_ (
    .A(\cpuregs[23] [10]),
    .ZN(_21378_)
  );
  INV_X1 _29494_ (
    .A(\cpuregs[23] [12]),
    .ZN(_21379_)
  );
  INV_X1 _29495_ (
    .A(\cpuregs[23] [13]),
    .ZN(_21380_)
  );
  INV_X1 _29496_ (
    .A(\cpuregs[23] [15]),
    .ZN(_21381_)
  );
  INV_X1 _29497_ (
    .A(\cpuregs[23] [16]),
    .ZN(_21382_)
  );
  INV_X1 _29498_ (
    .A(\cpuregs[23] [17]),
    .ZN(_21383_)
  );
  INV_X1 _29499_ (
    .A(\cpuregs[23] [19]),
    .ZN(_21384_)
  );
  INV_X1 _29500_ (
    .A(\cpuregs[23] [20]),
    .ZN(_21385_)
  );
  INV_X1 _29501_ (
    .A(\cpuregs[23] [22]),
    .ZN(_21386_)
  );
  INV_X1 _29502_ (
    .A(\cpuregs[23] [23]),
    .ZN(_21387_)
  );
  INV_X1 _29503_ (
    .A(\cpuregs[23] [24]),
    .ZN(_21388_)
  );
  INV_X1 _29504_ (
    .A(\cpuregs[23] [25]),
    .ZN(_21389_)
  );
  INV_X1 _29505_ (
    .A(\cpuregs[23] [26]),
    .ZN(_21390_)
  );
  INV_X1 _29506_ (
    .A(\cpuregs[23] [28]),
    .ZN(_21391_)
  );
  INV_X1 _29507_ (
    .A(\cpuregs[23] [29]),
    .ZN(_21392_)
  );
  INV_X1 _29508_ (
    .A(\cpuregs[14] [5]),
    .ZN(_21393_)
  );
  INV_X1 _29509_ (
    .A(\cpuregs[14] [6]),
    .ZN(_21394_)
  );
  INV_X1 _29510_ (
    .A(\cpuregs[14] [7]),
    .ZN(_21395_)
  );
  INV_X1 _29511_ (
    .A(\cpuregs[14] [15]),
    .ZN(_21396_)
  );
  INV_X1 _29512_ (
    .A(\cpuregs[14] [17]),
    .ZN(_21397_)
  );
  INV_X1 _29513_ (
    .A(\cpuregs[14] [23]),
    .ZN(_21398_)
  );
  INV_X1 _29514_ (
    .A(\cpuregs[14] [29]),
    .ZN(_21399_)
  );
  INV_X1 _29515_ (
    .A(\cpuregs[14] [30]),
    .ZN(_21400_)
  );
  INV_X1 _29516_ (
    .A(\cpuregs[15] [5]),
    .ZN(_21401_)
  );
  INV_X1 _29517_ (
    .A(\cpuregs[15] [6]),
    .ZN(_21402_)
  );
  INV_X1 _29518_ (
    .A(\cpuregs[15] [7]),
    .ZN(_21403_)
  );
  INV_X1 _29519_ (
    .A(\cpuregs[15] [17]),
    .ZN(_21404_)
  );
  INV_X1 _29520_ (
    .A(\cpuregs[15] [23]),
    .ZN(_21405_)
  );
  INV_X1 _29521_ (
    .A(\cpuregs[15] [29]),
    .ZN(_21406_)
  );
  INV_X1 _29522_ (
    .A(\cpuregs[15] [30]),
    .ZN(_21407_)
  );
  INV_X1 _29523_ (
    .A(\cpuregs[22] [0]),
    .ZN(_21408_)
  );
  INV_X1 _29524_ (
    .A(\cpuregs[22] [1]),
    .ZN(_21409_)
  );
  INV_X1 _29525_ (
    .A(\cpuregs[22] [2]),
    .ZN(_21410_)
  );
  INV_X1 _29526_ (
    .A(\cpuregs[22] [3]),
    .ZN(_21411_)
  );
  INV_X1 _29527_ (
    .A(\cpuregs[22] [4]),
    .ZN(_21412_)
  );
  INV_X1 _29528_ (
    .A(\cpuregs[22] [5]),
    .ZN(_21413_)
  );
  INV_X1 _29529_ (
    .A(\cpuregs[22] [6]),
    .ZN(_21414_)
  );
  INV_X1 _29530_ (
    .A(\cpuregs[22] [7]),
    .ZN(_21415_)
  );
  INV_X1 _29531_ (
    .A(\cpuregs[22] [8]),
    .ZN(_21416_)
  );
  INV_X1 _29532_ (
    .A(\cpuregs[22] [9]),
    .ZN(_21417_)
  );
  INV_X1 _29533_ (
    .A(\cpuregs[22] [10]),
    .ZN(_21418_)
  );
  INV_X1 _29534_ (
    .A(\cpuregs[22] [12]),
    .ZN(_21419_)
  );
  INV_X1 _29535_ (
    .A(\cpuregs[22] [13]),
    .ZN(_21420_)
  );
  INV_X1 _29536_ (
    .A(\cpuregs[22] [14]),
    .ZN(_21421_)
  );
  INV_X1 _29537_ (
    .A(\cpuregs[22] [15]),
    .ZN(_21422_)
  );
  INV_X1 _29538_ (
    .A(\cpuregs[22] [16]),
    .ZN(_21423_)
  );
  INV_X1 _29539_ (
    .A(\cpuregs[22] [17]),
    .ZN(_21424_)
  );
  INV_X1 _29540_ (
    .A(\cpuregs[22] [19]),
    .ZN(_21425_)
  );
  INV_X1 _29541_ (
    .A(\cpuregs[22] [20]),
    .ZN(_21426_)
  );
  INV_X1 _29542_ (
    .A(\cpuregs[22] [22]),
    .ZN(_21427_)
  );
  INV_X1 _29543_ (
    .A(\cpuregs[22] [23]),
    .ZN(_21428_)
  );
  INV_X1 _29544_ (
    .A(\cpuregs[22] [24]),
    .ZN(_21429_)
  );
  INV_X1 _29545_ (
    .A(\cpuregs[22] [25]),
    .ZN(_21430_)
  );
  INV_X1 _29546_ (
    .A(\cpuregs[22] [26]),
    .ZN(_21431_)
  );
  INV_X1 _29547_ (
    .A(\cpuregs[22] [27]),
    .ZN(_21432_)
  );
  INV_X1 _29548_ (
    .A(\cpuregs[22] [28]),
    .ZN(_21433_)
  );
  INV_X1 _29549_ (
    .A(\cpuregs[22] [29]),
    .ZN(_21434_)
  );
  INV_X1 _29550_ (
    .A(\cpuregs[22] [30]),
    .ZN(_21435_)
  );
  INV_X1 _29551_ (
    .A(\cpuregs[16] [0]),
    .ZN(_21436_)
  );
  INV_X1 _29552_ (
    .A(\cpuregs[16] [1]),
    .ZN(_21437_)
  );
  INV_X1 _29553_ (
    .A(\cpuregs[16] [2]),
    .ZN(_21438_)
  );
  INV_X1 _29554_ (
    .A(\cpuregs[16] [3]),
    .ZN(_21439_)
  );
  INV_X1 _29555_ (
    .A(\cpuregs[16] [4]),
    .ZN(_21440_)
  );
  INV_X1 _29556_ (
    .A(\cpuregs[16] [5]),
    .ZN(_21441_)
  );
  INV_X1 _29557_ (
    .A(\cpuregs[16] [7]),
    .ZN(_21442_)
  );
  INV_X1 _29558_ (
    .A(\cpuregs[16] [9]),
    .ZN(_21443_)
  );
  INV_X1 _29559_ (
    .A(\cpuregs[16] [10]),
    .ZN(_21444_)
  );
  INV_X1 _29560_ (
    .A(\cpuregs[16] [12]),
    .ZN(_21445_)
  );
  INV_X1 _29561_ (
    .A(\cpuregs[16] [13]),
    .ZN(_21446_)
  );
  INV_X1 _29562_ (
    .A(\cpuregs[16] [15]),
    .ZN(_21447_)
  );
  INV_X1 _29563_ (
    .A(\cpuregs[16] [16]),
    .ZN(_21448_)
  );
  INV_X1 _29564_ (
    .A(\cpuregs[16] [17]),
    .ZN(_21449_)
  );
  INV_X1 _29565_ (
    .A(\cpuregs[16] [19]),
    .ZN(_21450_)
  );
  INV_X1 _29566_ (
    .A(\cpuregs[16] [20]),
    .ZN(_21451_)
  );
  INV_X1 _29567_ (
    .A(\cpuregs[16] [22]),
    .ZN(_21452_)
  );
  INV_X1 _29568_ (
    .A(\cpuregs[16] [24]),
    .ZN(_21453_)
  );
  INV_X1 _29569_ (
    .A(\cpuregs[16] [25]),
    .ZN(_21454_)
  );
  INV_X1 _29570_ (
    .A(\cpuregs[16] [26]),
    .ZN(_21455_)
  );
  INV_X1 _29571_ (
    .A(\cpuregs[16] [28]),
    .ZN(_21456_)
  );
  INV_X1 _29572_ (
    .A(\cpuregs[16] [29]),
    .ZN(_21457_)
  );
  INV_X1 _29573_ (
    .A(\cpuregs[17] [0]),
    .ZN(_21458_)
  );
  INV_X1 _29574_ (
    .A(\cpuregs[17] [1]),
    .ZN(_21459_)
  );
  INV_X1 _29575_ (
    .A(\cpuregs[17] [2]),
    .ZN(_21460_)
  );
  INV_X1 _29576_ (
    .A(\cpuregs[17] [3]),
    .ZN(_21461_)
  );
  INV_X1 _29577_ (
    .A(\cpuregs[17] [4]),
    .ZN(_21462_)
  );
  INV_X1 _29578_ (
    .A(\cpuregs[17] [5]),
    .ZN(_21463_)
  );
  INV_X1 _29579_ (
    .A(\cpuregs[17] [7]),
    .ZN(_21464_)
  );
  INV_X1 _29580_ (
    .A(\cpuregs[17] [9]),
    .ZN(_21465_)
  );
  INV_X1 _29581_ (
    .A(\cpuregs[17] [10]),
    .ZN(_21466_)
  );
  INV_X1 _29582_ (
    .A(\cpuregs[17] [12]),
    .ZN(_21467_)
  );
  INV_X1 _29583_ (
    .A(\cpuregs[17] [13]),
    .ZN(_21468_)
  );
  INV_X1 _29584_ (
    .A(\cpuregs[17] [15]),
    .ZN(_21469_)
  );
  INV_X1 _29585_ (
    .A(\cpuregs[17] [16]),
    .ZN(_21470_)
  );
  INV_X1 _29586_ (
    .A(\cpuregs[17] [17]),
    .ZN(_21471_)
  );
  INV_X1 _29587_ (
    .A(\cpuregs[17] [19]),
    .ZN(_21472_)
  );
  INV_X1 _29588_ (
    .A(\cpuregs[17] [20]),
    .ZN(_21473_)
  );
  INV_X1 _29589_ (
    .A(\cpuregs[17] [22]),
    .ZN(_21474_)
  );
  INV_X1 _29590_ (
    .A(\cpuregs[17] [24]),
    .ZN(_21475_)
  );
  INV_X1 _29591_ (
    .A(\cpuregs[17] [25]),
    .ZN(_21476_)
  );
  INV_X1 _29592_ (
    .A(\cpuregs[17] [26]),
    .ZN(_21477_)
  );
  INV_X1 _29593_ (
    .A(\cpuregs[17] [28]),
    .ZN(_21478_)
  );
  INV_X1 _29594_ (
    .A(\cpuregs[17] [29]),
    .ZN(_21479_)
  );
  INV_X1 _29595_ (
    .A(\cpuregs[12] [5]),
    .ZN(_21480_)
  );
  INV_X1 _29596_ (
    .A(\cpuregs[12] [6]),
    .ZN(_21481_)
  );
  INV_X1 _29597_ (
    .A(\cpuregs[12] [7]),
    .ZN(_21482_)
  );
  INV_X1 _29598_ (
    .A(\cpuregs[12] [8]),
    .ZN(_21483_)
  );
  INV_X1 _29599_ (
    .A(\cpuregs[12] [23]),
    .ZN(_21484_)
  );
  INV_X1 _29600_ (
    .A(\cpuregs[12] [29]),
    .ZN(_21485_)
  );
  INV_X1 _29601_ (
    .A(\cpuregs[12] [30]),
    .ZN(_21486_)
  );
  INV_X1 _29602_ (
    .A(\cpuregs[3] [0]),
    .ZN(_21487_)
  );
  INV_X1 _29603_ (
    .A(\cpuregs[3] [1]),
    .ZN(_21488_)
  );
  INV_X1 _29604_ (
    .A(\cpuregs[3] [2]),
    .ZN(_21489_)
  );
  INV_X1 _29605_ (
    .A(\cpuregs[3] [3]),
    .ZN(_21490_)
  );
  INV_X1 _29606_ (
    .A(\cpuregs[3] [4]),
    .ZN(_21491_)
  );
  INV_X1 _29607_ (
    .A(\cpuregs[3] [5]),
    .ZN(_21492_)
  );
  INV_X1 _29608_ (
    .A(\cpuregs[3] [6]),
    .ZN(_21493_)
  );
  INV_X1 _29609_ (
    .A(\cpuregs[3] [7]),
    .ZN(_21494_)
  );
  INV_X1 _29610_ (
    .A(\cpuregs[3] [8]),
    .ZN(_21495_)
  );
  INV_X1 _29611_ (
    .A(\cpuregs[3] [11]),
    .ZN(_21496_)
  );
  INV_X1 _29612_ (
    .A(\cpuregs[3] [13]),
    .ZN(_21497_)
  );
  INV_X1 _29613_ (
    .A(\cpuregs[3] [14]),
    .ZN(_21498_)
  );
  INV_X1 _29614_ (
    .A(\cpuregs[3] [15]),
    .ZN(_21499_)
  );
  INV_X1 _29615_ (
    .A(\cpuregs[3] [16]),
    .ZN(_21500_)
  );
  INV_X1 _29616_ (
    .A(\cpuregs[3] [17]),
    .ZN(_21501_)
  );
  INV_X1 _29617_ (
    .A(\cpuregs[3] [18]),
    .ZN(_21502_)
  );
  INV_X1 _29618_ (
    .A(\cpuregs[3] [19]),
    .ZN(_21503_)
  );
  INV_X1 _29619_ (
    .A(\cpuregs[3] [21]),
    .ZN(_21504_)
  );
  INV_X1 _29620_ (
    .A(\cpuregs[3] [23]),
    .ZN(_21505_)
  );
  INV_X1 _29621_ (
    .A(\cpuregs[3] [25]),
    .ZN(_21506_)
  );
  INV_X1 _29622_ (
    .A(\cpuregs[3] [26]),
    .ZN(_21507_)
  );
  INV_X1 _29623_ (
    .A(\cpuregs[3] [27]),
    .ZN(_21508_)
  );
  INV_X1 _29624_ (
    .A(\cpuregs[3] [28]),
    .ZN(_21509_)
  );
  INV_X1 _29625_ (
    .A(\cpuregs[3] [29]),
    .ZN(_21510_)
  );
  INV_X1 _29626_ (
    .A(\cpuregs[3] [30]),
    .ZN(_21511_)
  );
  INV_X1 _29627_ (
    .A(\cpuregs[1] [0]),
    .ZN(_21512_)
  );
  INV_X1 _29628_ (
    .A(\cpuregs[1] [1]),
    .ZN(_21513_)
  );
  INV_X1 _29629_ (
    .A(\cpuregs[1] [2]),
    .ZN(_21514_)
  );
  INV_X1 _29630_ (
    .A(\cpuregs[1] [3]),
    .ZN(_21515_)
  );
  INV_X1 _29631_ (
    .A(\cpuregs[1] [4]),
    .ZN(_21516_)
  );
  INV_X1 _29632_ (
    .A(\cpuregs[1] [5]),
    .ZN(_21517_)
  );
  INV_X1 _29633_ (
    .A(\cpuregs[1] [6]),
    .ZN(_21518_)
  );
  INV_X1 _29634_ (
    .A(\cpuregs[1] [7]),
    .ZN(_21519_)
  );
  INV_X1 _29635_ (
    .A(\cpuregs[1] [8]),
    .ZN(_21520_)
  );
  INV_X1 _29636_ (
    .A(\cpuregs[1] [11]),
    .ZN(_21521_)
  );
  INV_X1 _29637_ (
    .A(\cpuregs[1] [13]),
    .ZN(_21522_)
  );
  INV_X1 _29638_ (
    .A(\cpuregs[1] [14]),
    .ZN(_21523_)
  );
  INV_X1 _29639_ (
    .A(\cpuregs[1] [15]),
    .ZN(_21524_)
  );
  INV_X1 _29640_ (
    .A(\cpuregs[1] [16]),
    .ZN(_21525_)
  );
  INV_X1 _29641_ (
    .A(\cpuregs[1] [17]),
    .ZN(_21526_)
  );
  INV_X1 _29642_ (
    .A(\cpuregs[1] [18]),
    .ZN(_21527_)
  );
  INV_X1 _29643_ (
    .A(\cpuregs[1] [19]),
    .ZN(_21528_)
  );
  INV_X1 _29644_ (
    .A(\cpuregs[1] [21]),
    .ZN(_21529_)
  );
  INV_X1 _29645_ (
    .A(\cpuregs[1] [23]),
    .ZN(_21530_)
  );
  INV_X1 _29646_ (
    .A(\cpuregs[1] [25]),
    .ZN(_21531_)
  );
  INV_X1 _29647_ (
    .A(\cpuregs[1] [26]),
    .ZN(_21532_)
  );
  INV_X1 _29648_ (
    .A(\cpuregs[1] [27]),
    .ZN(_21533_)
  );
  INV_X1 _29649_ (
    .A(\cpuregs[1] [28]),
    .ZN(_21534_)
  );
  INV_X1 _29650_ (
    .A(\cpuregs[1] [29]),
    .ZN(_21535_)
  );
  INV_X1 _29651_ (
    .A(\cpuregs[1] [30]),
    .ZN(_21536_)
  );
  INV_X1 _29652_ (
    .A(\cpuregs[2] [0]),
    .ZN(_21537_)
  );
  INV_X1 _29653_ (
    .A(\cpuregs[2] [1]),
    .ZN(_21538_)
  );
  INV_X1 _29654_ (
    .A(\cpuregs[2] [2]),
    .ZN(_21539_)
  );
  INV_X1 _29655_ (
    .A(\cpuregs[2] [3]),
    .ZN(_21540_)
  );
  INV_X1 _29656_ (
    .A(\cpuregs[2] [4]),
    .ZN(_21541_)
  );
  INV_X1 _29657_ (
    .A(\cpuregs[2] [5]),
    .ZN(_21542_)
  );
  INV_X1 _29658_ (
    .A(\cpuregs[2] [6]),
    .ZN(_21543_)
  );
  INV_X1 _29659_ (
    .A(\cpuregs[2] [7]),
    .ZN(_21544_)
  );
  INV_X1 _29660_ (
    .A(\cpuregs[2] [8]),
    .ZN(_21545_)
  );
  INV_X1 _29661_ (
    .A(\cpuregs[2] [9]),
    .ZN(_21546_)
  );
  INV_X1 _29662_ (
    .A(\cpuregs[2] [10]),
    .ZN(_21547_)
  );
  INV_X1 _29663_ (
    .A(\cpuregs[2] [11]),
    .ZN(_21548_)
  );
  INV_X1 _29664_ (
    .A(\cpuregs[2] [12]),
    .ZN(_21549_)
  );
  INV_X1 _29665_ (
    .A(\cpuregs[2] [13]),
    .ZN(_21550_)
  );
  INV_X1 _29666_ (
    .A(\cpuregs[2] [14]),
    .ZN(_21551_)
  );
  INV_X1 _29667_ (
    .A(\cpuregs[2] [15]),
    .ZN(_21552_)
  );
  INV_X1 _29668_ (
    .A(\cpuregs[2] [16]),
    .ZN(_21553_)
  );
  INV_X1 _29669_ (
    .A(\cpuregs[2] [17]),
    .ZN(_21554_)
  );
  INV_X1 _29670_ (
    .A(\cpuregs[2] [18]),
    .ZN(_21555_)
  );
  INV_X1 _29671_ (
    .A(\cpuregs[2] [19]),
    .ZN(_21556_)
  );
  INV_X1 _29672_ (
    .A(\cpuregs[2] [21]),
    .ZN(_21557_)
  );
  INV_X1 _29673_ (
    .A(\cpuregs[2] [22]),
    .ZN(_21558_)
  );
  INV_X1 _29674_ (
    .A(\cpuregs[2] [23]),
    .ZN(_21559_)
  );
  INV_X1 _29675_ (
    .A(\cpuregs[2] [24]),
    .ZN(_21560_)
  );
  INV_X1 _29676_ (
    .A(\cpuregs[2] [25]),
    .ZN(_21561_)
  );
  INV_X1 _29677_ (
    .A(\cpuregs[2] [26]),
    .ZN(_21562_)
  );
  INV_X1 _29678_ (
    .A(\cpuregs[2] [27]),
    .ZN(_21563_)
  );
  INV_X1 _29679_ (
    .A(\cpuregs[2] [28]),
    .ZN(_21564_)
  );
  INV_X1 _29680_ (
    .A(\cpuregs[2] [29]),
    .ZN(_21565_)
  );
  INV_X1 _29681_ (
    .A(\cpuregs[2] [30]),
    .ZN(_21566_)
  );
  INV_X1 _29682_ (
    .A(\cpuregs[24] [0]),
    .ZN(_21567_)
  );
  INV_X1 _29683_ (
    .A(\cpuregs[24] [1]),
    .ZN(_21568_)
  );
  INV_X1 _29684_ (
    .A(\cpuregs[24] [2]),
    .ZN(_21569_)
  );
  INV_X1 _29685_ (
    .A(\cpuregs[24] [5]),
    .ZN(_21570_)
  );
  INV_X1 _29686_ (
    .A(\cpuregs[24] [6]),
    .ZN(_21571_)
  );
  INV_X1 _29687_ (
    .A(\cpuregs[24] [7]),
    .ZN(_21572_)
  );
  INV_X1 _29688_ (
    .A(\cpuregs[24] [9]),
    .ZN(_21573_)
  );
  INV_X1 _29689_ (
    .A(\cpuregs[24] [13]),
    .ZN(_21574_)
  );
  INV_X1 _29690_ (
    .A(\cpuregs[24] [15]),
    .ZN(_21575_)
  );
  INV_X1 _29691_ (
    .A(\cpuregs[24] [16]),
    .ZN(_21576_)
  );
  INV_X1 _29692_ (
    .A(\cpuregs[24] [19]),
    .ZN(_21577_)
  );
  INV_X1 _29693_ (
    .A(\cpuregs[24] [23]),
    .ZN(_21578_)
  );
  INV_X1 _29694_ (
    .A(\cpuregs[24] [25]),
    .ZN(_21579_)
  );
  INV_X1 _29695_ (
    .A(\cpuregs[24] [26]),
    .ZN(_21580_)
  );
  INV_X1 _29696_ (
    .A(\cpuregs[24] [28]),
    .ZN(_21581_)
  );
  INV_X1 _29697_ (
    .A(\cpuregs[24] [29]),
    .ZN(_21582_)
  );
  INV_X1 _29698_ (
    .A(\cpuregs[11] [5]),
    .ZN(_21583_)
  );
  INV_X1 _29699_ (
    .A(\cpuregs[11] [6]),
    .ZN(_21584_)
  );
  INV_X1 _29700_ (
    .A(\cpuregs[11] [7]),
    .ZN(_21585_)
  );
  INV_X1 _29701_ (
    .A(\cpuregs[11] [17]),
    .ZN(_21586_)
  );
  INV_X1 _29702_ (
    .A(\cpuregs[11] [23]),
    .ZN(_21587_)
  );
  INV_X1 _29703_ (
    .A(\cpuregs[11] [29]),
    .ZN(_21588_)
  );
  INV_X1 _29704_ (
    .A(\cpuregs[11] [30]),
    .ZN(_21589_)
  );
  INV_X1 _29705_ (
    .A(\cpuregs[18] [0]),
    .ZN(_21590_)
  );
  INV_X1 _29706_ (
    .A(\cpuregs[18] [1]),
    .ZN(_21591_)
  );
  INV_X1 _29707_ (
    .A(\cpuregs[18] [2]),
    .ZN(_21592_)
  );
  INV_X1 _29708_ (
    .A(\cpuregs[18] [3]),
    .ZN(_21593_)
  );
  INV_X1 _29709_ (
    .A(\cpuregs[18] [4]),
    .ZN(_21594_)
  );
  INV_X1 _29710_ (
    .A(\cpuregs[18] [5]),
    .ZN(_21595_)
  );
  INV_X1 _29711_ (
    .A(\cpuregs[18] [7]),
    .ZN(_21596_)
  );
  INV_X1 _29712_ (
    .A(\cpuregs[18] [9]),
    .ZN(_21597_)
  );
  INV_X1 _29713_ (
    .A(\cpuregs[18] [10]),
    .ZN(_21598_)
  );
  INV_X1 _29714_ (
    .A(\cpuregs[18] [12]),
    .ZN(_21599_)
  );
  INV_X1 _29715_ (
    .A(\cpuregs[18] [13]),
    .ZN(_21600_)
  );
  INV_X1 _29716_ (
    .A(\cpuregs[18] [14]),
    .ZN(_21601_)
  );
  INV_X1 _29717_ (
    .A(\cpuregs[18] [15]),
    .ZN(_21602_)
  );
  INV_X1 _29718_ (
    .A(\cpuregs[18] [16]),
    .ZN(_21603_)
  );
  INV_X1 _29719_ (
    .A(\cpuregs[18] [17]),
    .ZN(_21604_)
  );
  INV_X1 _29720_ (
    .A(\cpuregs[18] [19]),
    .ZN(_21605_)
  );
  INV_X1 _29721_ (
    .A(\cpuregs[18] [20]),
    .ZN(_21606_)
  );
  INV_X1 _29722_ (
    .A(\cpuregs[18] [22]),
    .ZN(_21607_)
  );
  INV_X1 _29723_ (
    .A(\cpuregs[18] [23]),
    .ZN(_21608_)
  );
  INV_X1 _29724_ (
    .A(\cpuregs[18] [24]),
    .ZN(_21609_)
  );
  INV_X1 _29725_ (
    .A(\cpuregs[18] [25]),
    .ZN(_21610_)
  );
  INV_X1 _29726_ (
    .A(\cpuregs[18] [26]),
    .ZN(_21611_)
  );
  INV_X1 _29727_ (
    .A(\cpuregs[18] [27]),
    .ZN(_21612_)
  );
  INV_X1 _29728_ (
    .A(\cpuregs[18] [28]),
    .ZN(_21613_)
  );
  INV_X1 _29729_ (
    .A(\cpuregs[18] [29]),
    .ZN(_21614_)
  );
  INV_X1 _29730_ (
    .A(\cpuregs[18] [30]),
    .ZN(_21615_)
  );
  INV_X1 _29731_ (
    .A(\cpuregs[19] [0]),
    .ZN(_21616_)
  );
  INV_X1 _29732_ (
    .A(\cpuregs[19] [1]),
    .ZN(_21617_)
  );
  INV_X1 _29733_ (
    .A(\cpuregs[19] [2]),
    .ZN(_21618_)
  );
  INV_X1 _29734_ (
    .A(\cpuregs[19] [3]),
    .ZN(_21619_)
  );
  INV_X1 _29735_ (
    .A(\cpuregs[19] [4]),
    .ZN(_21620_)
  );
  INV_X1 _29736_ (
    .A(\cpuregs[19] [5]),
    .ZN(_21621_)
  );
  INV_X1 _29737_ (
    .A(\cpuregs[19] [7]),
    .ZN(_21622_)
  );
  INV_X1 _29738_ (
    .A(\cpuregs[19] [9]),
    .ZN(_21623_)
  );
  INV_X1 _29739_ (
    .A(\cpuregs[19] [10]),
    .ZN(_21624_)
  );
  INV_X1 _29740_ (
    .A(\cpuregs[19] [12]),
    .ZN(_21625_)
  );
  INV_X1 _29741_ (
    .A(\cpuregs[19] [13]),
    .ZN(_21626_)
  );
  INV_X1 _29742_ (
    .A(\cpuregs[19] [15]),
    .ZN(_21627_)
  );
  INV_X1 _29743_ (
    .A(\cpuregs[19] [16]),
    .ZN(_21628_)
  );
  INV_X1 _29744_ (
    .A(\cpuregs[19] [17]),
    .ZN(_21629_)
  );
  INV_X1 _29745_ (
    .A(\cpuregs[19] [19]),
    .ZN(_21630_)
  );
  INV_X1 _29746_ (
    .A(\cpuregs[19] [20]),
    .ZN(_21631_)
  );
  INV_X1 _29747_ (
    .A(\cpuregs[19] [22]),
    .ZN(_21632_)
  );
  INV_X1 _29748_ (
    .A(\cpuregs[19] [23]),
    .ZN(_21633_)
  );
  INV_X1 _29749_ (
    .A(\cpuregs[19] [24]),
    .ZN(_21634_)
  );
  INV_X1 _29750_ (
    .A(\cpuregs[19] [25]),
    .ZN(_21635_)
  );
  INV_X1 _29751_ (
    .A(\cpuregs[19] [26]),
    .ZN(_21636_)
  );
  INV_X1 _29752_ (
    .A(\cpuregs[19] [28]),
    .ZN(_21637_)
  );
  INV_X1 _29753_ (
    .A(\cpuregs[19] [29]),
    .ZN(_21638_)
  );
  INV_X1 _29754_ (
    .A(\cpuregs[13] [5]),
    .ZN(_21639_)
  );
  INV_X1 _29755_ (
    .A(\cpuregs[13] [6]),
    .ZN(_21640_)
  );
  INV_X1 _29756_ (
    .A(\cpuregs[13] [7]),
    .ZN(_21641_)
  );
  INV_X1 _29757_ (
    .A(\cpuregs[13] [8]),
    .ZN(_21642_)
  );
  INV_X1 _29758_ (
    .A(\cpuregs[13] [17]),
    .ZN(_21643_)
  );
  INV_X1 _29759_ (
    .A(\cpuregs[13] [23]),
    .ZN(_21644_)
  );
  INV_X1 _29760_ (
    .A(\cpuregs[13] [29]),
    .ZN(_21645_)
  );
  INV_X1 _29761_ (
    .A(\cpuregs[13] [30]),
    .ZN(_21646_)
  );
  INV_X1 _29762_ (
    .A(\cpuregs[20] [0]),
    .ZN(_21647_)
  );
  INV_X1 _29763_ (
    .A(\cpuregs[20] [1]),
    .ZN(_21648_)
  );
  INV_X1 _29764_ (
    .A(\cpuregs[20] [2]),
    .ZN(_21649_)
  );
  INV_X1 _29765_ (
    .A(\cpuregs[20] [3]),
    .ZN(_21650_)
  );
  INV_X1 _29766_ (
    .A(\cpuregs[20] [4]),
    .ZN(_21651_)
  );
  INV_X1 _29767_ (
    .A(\cpuregs[20] [5]),
    .ZN(_21652_)
  );
  INV_X1 _29768_ (
    .A(\cpuregs[20] [7]),
    .ZN(_21653_)
  );
  INV_X1 _29769_ (
    .A(\cpuregs[20] [9]),
    .ZN(_21654_)
  );
  INV_X1 _29770_ (
    .A(\cpuregs[20] [10]),
    .ZN(_21655_)
  );
  INV_X1 _29771_ (
    .A(\cpuregs[20] [12]),
    .ZN(_21656_)
  );
  INV_X1 _29772_ (
    .A(\cpuregs[20] [13]),
    .ZN(_21657_)
  );
  INV_X1 _29773_ (
    .A(\cpuregs[20] [15]),
    .ZN(_21658_)
  );
  INV_X1 _29774_ (
    .A(\cpuregs[20] [16]),
    .ZN(_21659_)
  );
  INV_X1 _29775_ (
    .A(\cpuregs[20] [17]),
    .ZN(_21660_)
  );
  INV_X1 _29776_ (
    .A(\cpuregs[20] [19]),
    .ZN(_21661_)
  );
  INV_X1 _29777_ (
    .A(\cpuregs[20] [20]),
    .ZN(_21662_)
  );
  INV_X1 _29778_ (
    .A(\cpuregs[20] [22]),
    .ZN(_21663_)
  );
  INV_X1 _29779_ (
    .A(\cpuregs[20] [24]),
    .ZN(_21664_)
  );
  INV_X1 _29780_ (
    .A(\cpuregs[20] [25]),
    .ZN(_21665_)
  );
  INV_X1 _29781_ (
    .A(\cpuregs[20] [26]),
    .ZN(_21666_)
  );
  INV_X1 _29782_ (
    .A(\cpuregs[20] [28]),
    .ZN(_21667_)
  );
  INV_X1 _29783_ (
    .A(\cpuregs[20] [29]),
    .ZN(_21668_)
  );
  INV_X1 _29784_ (
    .A(\cpuregs[4] [0]),
    .ZN(_21669_)
  );
  INV_X1 _29785_ (
    .A(\cpuregs[4] [1]),
    .ZN(_21670_)
  );
  INV_X1 _29786_ (
    .A(\cpuregs[4] [2]),
    .ZN(_21671_)
  );
  INV_X1 _29787_ (
    .A(\cpuregs[4] [3]),
    .ZN(_21672_)
  );
  INV_X1 _29788_ (
    .A(\cpuregs[4] [4]),
    .ZN(_21673_)
  );
  INV_X1 _29789_ (
    .A(\cpuregs[4] [5]),
    .ZN(_21674_)
  );
  INV_X1 _29790_ (
    .A(\cpuregs[4] [6]),
    .ZN(_21675_)
  );
  INV_X1 _29791_ (
    .A(\cpuregs[4] [7]),
    .ZN(_21676_)
  );
  INV_X1 _29792_ (
    .A(\cpuregs[4] [8]),
    .ZN(_21677_)
  );
  INV_X1 _29793_ (
    .A(\cpuregs[4] [11]),
    .ZN(_21678_)
  );
  INV_X1 _29794_ (
    .A(\cpuregs[4] [13]),
    .ZN(_21679_)
  );
  INV_X1 _29795_ (
    .A(\cpuregs[4] [14]),
    .ZN(_21680_)
  );
  INV_X1 _29796_ (
    .A(\cpuregs[4] [15]),
    .ZN(_21681_)
  );
  INV_X1 _29797_ (
    .A(\cpuregs[4] [16]),
    .ZN(_21682_)
  );
  INV_X1 _29798_ (
    .A(\cpuregs[4] [17]),
    .ZN(_21683_)
  );
  INV_X1 _29799_ (
    .A(\cpuregs[4] [18]),
    .ZN(_21684_)
  );
  INV_X1 _29800_ (
    .A(\cpuregs[4] [19]),
    .ZN(_21685_)
  );
  INV_X1 _29801_ (
    .A(\cpuregs[4] [21]),
    .ZN(_21686_)
  );
  INV_X1 _29802_ (
    .A(\cpuregs[4] [23]),
    .ZN(_21687_)
  );
  INV_X1 _29803_ (
    .A(\cpuregs[4] [25]),
    .ZN(_21688_)
  );
  INV_X1 _29804_ (
    .A(\cpuregs[4] [26]),
    .ZN(_21689_)
  );
  INV_X1 _29805_ (
    .A(\cpuregs[4] [27]),
    .ZN(_21690_)
  );
  INV_X1 _29806_ (
    .A(\cpuregs[4] [28]),
    .ZN(_21691_)
  );
  INV_X1 _29807_ (
    .A(\cpuregs[4] [29]),
    .ZN(_21692_)
  );
  INV_X1 _29808_ (
    .A(\cpuregs[4] [30]),
    .ZN(_21693_)
  );
  INV_X1 _29809_ (
    .A(\cpuregs[10] [0]),
    .ZN(_21694_)
  );
  INV_X1 _29810_ (
    .A(\cpuregs[10] [1]),
    .ZN(_21695_)
  );
  INV_X1 _29811_ (
    .A(\cpuregs[10] [2]),
    .ZN(_21696_)
  );
  INV_X1 _29812_ (
    .A(\cpuregs[10] [3]),
    .ZN(_21697_)
  );
  INV_X1 _29813_ (
    .A(\cpuregs[10] [5]),
    .ZN(_21698_)
  );
  INV_X1 _29814_ (
    .A(\cpuregs[10] [6]),
    .ZN(_21699_)
  );
  INV_X1 _29815_ (
    .A(\cpuregs[10] [7]),
    .ZN(_21700_)
  );
  INV_X1 _29816_ (
    .A(\cpuregs[10] [9]),
    .ZN(_21701_)
  );
  INV_X1 _29817_ (
    .A(\cpuregs[10] [10]),
    .ZN(_21702_)
  );
  INV_X1 _29818_ (
    .A(\cpuregs[10] [11]),
    .ZN(_21703_)
  );
  INV_X1 _29819_ (
    .A(\cpuregs[10] [12]),
    .ZN(_21704_)
  );
  INV_X1 _29820_ (
    .A(\cpuregs[10] [13]),
    .ZN(_21705_)
  );
  INV_X1 _29821_ (
    .A(\cpuregs[10] [15]),
    .ZN(_21706_)
  );
  INV_X1 _29822_ (
    .A(\cpuregs[10] [17]),
    .ZN(_21707_)
  );
  INV_X1 _29823_ (
    .A(\cpuregs[10] [19]),
    .ZN(_21708_)
  );
  INV_X1 _29824_ (
    .A(\cpuregs[10] [22]),
    .ZN(_21709_)
  );
  INV_X1 _29825_ (
    .A(\cpuregs[10] [23]),
    .ZN(_21710_)
  );
  INV_X1 _29826_ (
    .A(\cpuregs[10] [25]),
    .ZN(_21711_)
  );
  INV_X1 _29827_ (
    .A(\cpuregs[10] [26]),
    .ZN(_21712_)
  );
  INV_X1 _29828_ (
    .A(\cpuregs[10] [27]),
    .ZN(_21713_)
  );
  INV_X1 _29829_ (
    .A(\cpuregs[10] [28]),
    .ZN(_21714_)
  );
  INV_X1 _29830_ (
    .A(\cpuregs[10] [29]),
    .ZN(_21715_)
  );
  INV_X1 _29831_ (
    .A(\cpuregs[10] [30]),
    .ZN(_21716_)
  );
  INV_X1 _29832_ (
    .A(\cpuregs[9] [5]),
    .ZN(_21717_)
  );
  INV_X1 _29833_ (
    .A(\cpuregs[9] [6]),
    .ZN(_21718_)
  );
  INV_X1 _29834_ (
    .A(\cpuregs[9] [7]),
    .ZN(_21719_)
  );
  INV_X1 _29835_ (
    .A(\cpuregs[9] [8]),
    .ZN(_21720_)
  );
  INV_X1 _29836_ (
    .A(\cpuregs[9] [17]),
    .ZN(_21721_)
  );
  INV_X1 _29837_ (
    .A(\cpuregs[9] [23]),
    .ZN(_21722_)
  );
  INV_X1 _29838_ (
    .A(\cpuregs[9] [29]),
    .ZN(_21723_)
  );
  INV_X1 _29839_ (
    .A(\cpuregs[9] [30]),
    .ZN(_21724_)
  );
  INV_X1 _29840_ (
    .A(\cpuregs[8] [5]),
    .ZN(_21725_)
  );
  INV_X1 _29841_ (
    .A(\cpuregs[8] [6]),
    .ZN(_21726_)
  );
  INV_X1 _29842_ (
    .A(\cpuregs[8] [7]),
    .ZN(_21727_)
  );
  INV_X1 _29843_ (
    .A(\cpuregs[8] [8]),
    .ZN(_21728_)
  );
  INV_X1 _29844_ (
    .A(\cpuregs[8] [23]),
    .ZN(_21729_)
  );
  INV_X1 _29845_ (
    .A(\cpuregs[8] [29]),
    .ZN(_21730_)
  );
  INV_X1 _29846_ (
    .A(\cpuregs[8] [30]),
    .ZN(_21731_)
  );
  INV_X1 _29847_ (
    .A(\cpuregs[5] [0]),
    .ZN(_21732_)
  );
  INV_X1 _29848_ (
    .A(\cpuregs[5] [1]),
    .ZN(_21733_)
  );
  INV_X1 _29849_ (
    .A(\cpuregs[5] [2]),
    .ZN(_21734_)
  );
  INV_X1 _29850_ (
    .A(\cpuregs[5] [3]),
    .ZN(_21735_)
  );
  INV_X1 _29851_ (
    .A(\cpuregs[5] [4]),
    .ZN(_21736_)
  );
  INV_X1 _29852_ (
    .A(\cpuregs[5] [5]),
    .ZN(_21737_)
  );
  INV_X1 _29853_ (
    .A(\cpuregs[5] [6]),
    .ZN(_21738_)
  );
  INV_X1 _29854_ (
    .A(\cpuregs[5] [7]),
    .ZN(_21739_)
  );
  INV_X1 _29855_ (
    .A(\cpuregs[5] [8]),
    .ZN(_21740_)
  );
  INV_X1 _29856_ (
    .A(\cpuregs[5] [11]),
    .ZN(_21741_)
  );
  INV_X1 _29857_ (
    .A(\cpuregs[5] [13]),
    .ZN(_21742_)
  );
  INV_X1 _29858_ (
    .A(\cpuregs[5] [14]),
    .ZN(_21743_)
  );
  INV_X1 _29859_ (
    .A(\cpuregs[5] [15]),
    .ZN(_21744_)
  );
  INV_X1 _29860_ (
    .A(\cpuregs[5] [16]),
    .ZN(_21745_)
  );
  INV_X1 _29861_ (
    .A(\cpuregs[5] [17]),
    .ZN(_21746_)
  );
  INV_X1 _29862_ (
    .A(\cpuregs[5] [18]),
    .ZN(_21747_)
  );
  INV_X1 _29863_ (
    .A(\cpuregs[5] [19]),
    .ZN(_21748_)
  );
  INV_X1 _29864_ (
    .A(\cpuregs[5] [21]),
    .ZN(_21749_)
  );
  INV_X1 _29865_ (
    .A(\cpuregs[5] [23]),
    .ZN(_21750_)
  );
  INV_X1 _29866_ (
    .A(\cpuregs[5] [25]),
    .ZN(_21751_)
  );
  INV_X1 _29867_ (
    .A(\cpuregs[5] [26]),
    .ZN(_21752_)
  );
  INV_X1 _29868_ (
    .A(\cpuregs[5] [27]),
    .ZN(_21753_)
  );
  INV_X1 _29869_ (
    .A(\cpuregs[5] [28]),
    .ZN(_21754_)
  );
  INV_X1 _29870_ (
    .A(\cpuregs[5] [29]),
    .ZN(_21755_)
  );
  INV_X1 _29871_ (
    .A(\cpuregs[5] [30]),
    .ZN(_21756_)
  );
  INV_X1 _29872_ (
    .A(\cpuregs[21] [0]),
    .ZN(_21757_)
  );
  INV_X1 _29873_ (
    .A(\cpuregs[21] [1]),
    .ZN(_21758_)
  );
  INV_X1 _29874_ (
    .A(\cpuregs[21] [2]),
    .ZN(_21759_)
  );
  INV_X1 _29875_ (
    .A(\cpuregs[21] [3]),
    .ZN(_21760_)
  );
  INV_X1 _29876_ (
    .A(\cpuregs[21] [4]),
    .ZN(_21761_)
  );
  INV_X1 _29877_ (
    .A(\cpuregs[21] [5]),
    .ZN(_21762_)
  );
  INV_X1 _29878_ (
    .A(\cpuregs[21] [7]),
    .ZN(_21763_)
  );
  INV_X1 _29879_ (
    .A(\cpuregs[21] [9]),
    .ZN(_21764_)
  );
  INV_X1 _29880_ (
    .A(\cpuregs[21] [10]),
    .ZN(_21765_)
  );
  INV_X1 _29881_ (
    .A(\cpuregs[21] [12]),
    .ZN(_21766_)
  );
  INV_X1 _29882_ (
    .A(\cpuregs[21] [13]),
    .ZN(_21767_)
  );
  INV_X1 _29883_ (
    .A(\cpuregs[21] [15]),
    .ZN(_21768_)
  );
  INV_X1 _29884_ (
    .A(\cpuregs[21] [16]),
    .ZN(_21769_)
  );
  INV_X1 _29885_ (
    .A(\cpuregs[21] [17]),
    .ZN(_21770_)
  );
  INV_X1 _29886_ (
    .A(\cpuregs[21] [19]),
    .ZN(_21771_)
  );
  INV_X1 _29887_ (
    .A(\cpuregs[21] [20]),
    .ZN(_21772_)
  );
  INV_X1 _29888_ (
    .A(\cpuregs[21] [22]),
    .ZN(_21773_)
  );
  INV_X1 _29889_ (
    .A(\cpuregs[21] [24]),
    .ZN(_21774_)
  );
  INV_X1 _29890_ (
    .A(\cpuregs[21] [25]),
    .ZN(_21775_)
  );
  INV_X1 _29891_ (
    .A(\cpuregs[21] [26]),
    .ZN(_21776_)
  );
  INV_X1 _29892_ (
    .A(\cpuregs[21] [28]),
    .ZN(_21777_)
  );
  INV_X1 _29893_ (
    .A(\cpuregs[21] [29]),
    .ZN(_21778_)
  );
  INV_X1 _29894_ (
    .A(\cpuregs[7] [0]),
    .ZN(_21779_)
  );
  INV_X1 _29895_ (
    .A(\cpuregs[7] [1]),
    .ZN(_21780_)
  );
  INV_X1 _29896_ (
    .A(\cpuregs[7] [2]),
    .ZN(_21781_)
  );
  INV_X1 _29897_ (
    .A(\cpuregs[7] [3]),
    .ZN(_21782_)
  );
  INV_X1 _29898_ (
    .A(\cpuregs[7] [4]),
    .ZN(_21783_)
  );
  INV_X1 _29899_ (
    .A(\cpuregs[7] [5]),
    .ZN(_21784_)
  );
  INV_X1 _29900_ (
    .A(\cpuregs[7] [6]),
    .ZN(_21785_)
  );
  INV_X1 _29901_ (
    .A(\cpuregs[7] [7]),
    .ZN(_21786_)
  );
  INV_X1 _29902_ (
    .A(\cpuregs[7] [8]),
    .ZN(_21787_)
  );
  INV_X1 _29903_ (
    .A(\cpuregs[7] [11]),
    .ZN(_21788_)
  );
  INV_X1 _29904_ (
    .A(\cpuregs[7] [13]),
    .ZN(_21789_)
  );
  INV_X1 _29905_ (
    .A(\cpuregs[7] [14]),
    .ZN(_21790_)
  );
  INV_X1 _29906_ (
    .A(\cpuregs[7] [15]),
    .ZN(_21791_)
  );
  INV_X1 _29907_ (
    .A(\cpuregs[7] [16]),
    .ZN(_21792_)
  );
  INV_X1 _29908_ (
    .A(\cpuregs[7] [17]),
    .ZN(_21793_)
  );
  INV_X1 _29909_ (
    .A(\cpuregs[7] [18]),
    .ZN(_21794_)
  );
  INV_X1 _29910_ (
    .A(\cpuregs[7] [19]),
    .ZN(_21795_)
  );
  INV_X1 _29911_ (
    .A(\cpuregs[7] [21]),
    .ZN(_21796_)
  );
  INV_X1 _29912_ (
    .A(\cpuregs[7] [23]),
    .ZN(_21797_)
  );
  INV_X1 _29913_ (
    .A(\cpuregs[7] [25]),
    .ZN(_21798_)
  );
  INV_X1 _29914_ (
    .A(\cpuregs[7] [26]),
    .ZN(_21799_)
  );
  INV_X1 _29915_ (
    .A(\cpuregs[7] [27]),
    .ZN(_21800_)
  );
  INV_X1 _29916_ (
    .A(\cpuregs[7] [28]),
    .ZN(_21801_)
  );
  INV_X1 _29917_ (
    .A(\cpuregs[7] [29]),
    .ZN(_21802_)
  );
  INV_X1 _29918_ (
    .A(\cpuregs[7] [30]),
    .ZN(_21803_)
  );
  INV_X1 _29919_ (
    .A(\cpuregs[6] [0]),
    .ZN(_21804_)
  );
  INV_X1 _29920_ (
    .A(\cpuregs[6] [1]),
    .ZN(_21805_)
  );
  INV_X1 _29921_ (
    .A(\cpuregs[6] [2]),
    .ZN(_21806_)
  );
  INV_X1 _29922_ (
    .A(\cpuregs[6] [3]),
    .ZN(_21807_)
  );
  INV_X1 _29923_ (
    .A(\cpuregs[6] [4]),
    .ZN(_21808_)
  );
  INV_X1 _29924_ (
    .A(\cpuregs[6] [5]),
    .ZN(_21809_)
  );
  INV_X1 _29925_ (
    .A(\cpuregs[6] [6]),
    .ZN(_21810_)
  );
  INV_X1 _29926_ (
    .A(\cpuregs[6] [7]),
    .ZN(_21811_)
  );
  INV_X1 _29927_ (
    .A(\cpuregs[6] [8]),
    .ZN(_21812_)
  );
  INV_X1 _29928_ (
    .A(\cpuregs[6] [10]),
    .ZN(_21813_)
  );
  INV_X1 _29929_ (
    .A(\cpuregs[6] [11]),
    .ZN(_21814_)
  );
  INV_X1 _29930_ (
    .A(\cpuregs[6] [12]),
    .ZN(_21815_)
  );
  INV_X1 _29931_ (
    .A(\cpuregs[6] [13]),
    .ZN(_21816_)
  );
  INV_X1 _29932_ (
    .A(\cpuregs[6] [14]),
    .ZN(_21817_)
  );
  INV_X1 _29933_ (
    .A(\cpuregs[6] [15]),
    .ZN(_21818_)
  );
  INV_X1 _29934_ (
    .A(\cpuregs[6] [16]),
    .ZN(_21819_)
  );
  INV_X1 _29935_ (
    .A(\cpuregs[6] [17]),
    .ZN(_21820_)
  );
  INV_X1 _29936_ (
    .A(\cpuregs[6] [18]),
    .ZN(_21821_)
  );
  INV_X1 _29937_ (
    .A(\cpuregs[6] [19]),
    .ZN(_21822_)
  );
  INV_X1 _29938_ (
    .A(\cpuregs[6] [21]),
    .ZN(_21823_)
  );
  INV_X1 _29939_ (
    .A(\cpuregs[6] [22]),
    .ZN(_21824_)
  );
  INV_X1 _29940_ (
    .A(\cpuregs[6] [23]),
    .ZN(_21825_)
  );
  INV_X1 _29941_ (
    .A(\cpuregs[6] [24]),
    .ZN(_21826_)
  );
  INV_X1 _29942_ (
    .A(\cpuregs[6] [25]),
    .ZN(_21827_)
  );
  INV_X1 _29943_ (
    .A(\cpuregs[6] [26]),
    .ZN(_21828_)
  );
  INV_X1 _29944_ (
    .A(\cpuregs[6] [27]),
    .ZN(_21829_)
  );
  INV_X1 _29945_ (
    .A(\cpuregs[6] [28]),
    .ZN(_21830_)
  );
  INV_X1 _29946_ (
    .A(\cpuregs[6] [29]),
    .ZN(_21831_)
  );
  INV_X1 _29947_ (
    .A(\cpuregs[6] [30]),
    .ZN(_21832_)
  );
  INV_X1 _29948_ (
    .A(\cpuregs[25] [0]),
    .ZN(_21833_)
  );
  INV_X1 _29949_ (
    .A(\cpuregs[25] [1]),
    .ZN(_21834_)
  );
  INV_X1 _29950_ (
    .A(\cpuregs[25] [2]),
    .ZN(_21835_)
  );
  INV_X1 _29951_ (
    .A(\cpuregs[25] [5]),
    .ZN(_21836_)
  );
  INV_X1 _29952_ (
    .A(\cpuregs[25] [6]),
    .ZN(_21837_)
  );
  INV_X1 _29953_ (
    .A(\cpuregs[25] [7]),
    .ZN(_21838_)
  );
  INV_X1 _29954_ (
    .A(\cpuregs[25] [9]),
    .ZN(_21839_)
  );
  INV_X1 _29955_ (
    .A(\cpuregs[25] [13]),
    .ZN(_21840_)
  );
  INV_X1 _29956_ (
    .A(\cpuregs[25] [15]),
    .ZN(_21841_)
  );
  INV_X1 _29957_ (
    .A(\cpuregs[25] [16]),
    .ZN(_21842_)
  );
  INV_X1 _29958_ (
    .A(\cpuregs[25] [19]),
    .ZN(_21843_)
  );
  INV_X1 _29959_ (
    .A(\cpuregs[25] [23]),
    .ZN(_21844_)
  );
  INV_X1 _29960_ (
    .A(\cpuregs[25] [25]),
    .ZN(_21845_)
  );
  INV_X1 _29961_ (
    .A(\cpuregs[25] [26]),
    .ZN(_21846_)
  );
  INV_X1 _29962_ (
    .A(\cpuregs[25] [28]),
    .ZN(_21847_)
  );
  INV_X1 _29963_ (
    .A(\cpuregs[25] [29]),
    .ZN(_21848_)
  );
  INV_X1 _29964_ (
    .A(\cpuregs[30] [0]),
    .ZN(_21849_)
  );
  INV_X1 _29965_ (
    .A(\cpuregs[30] [1]),
    .ZN(_21850_)
  );
  INV_X1 _29966_ (
    .A(\cpuregs[30] [2]),
    .ZN(_21851_)
  );
  INV_X1 _29967_ (
    .A(\cpuregs[30] [5]),
    .ZN(_21852_)
  );
  INV_X1 _29968_ (
    .A(\cpuregs[30] [6]),
    .ZN(_21853_)
  );
  INV_X1 _29969_ (
    .A(\cpuregs[30] [7]),
    .ZN(_21854_)
  );
  INV_X1 _29970_ (
    .A(\cpuregs[30] [9]),
    .ZN(_21855_)
  );
  INV_X1 _29971_ (
    .A(\cpuregs[30] [13]),
    .ZN(_21856_)
  );
  INV_X1 _29972_ (
    .A(\cpuregs[30] [15]),
    .ZN(_21857_)
  );
  INV_X1 _29973_ (
    .A(\cpuregs[30] [16]),
    .ZN(_21858_)
  );
  INV_X1 _29974_ (
    .A(\cpuregs[30] [19]),
    .ZN(_21859_)
  );
  INV_X1 _29975_ (
    .A(\cpuregs[30] [23]),
    .ZN(_21860_)
  );
  INV_X1 _29976_ (
    .A(\cpuregs[30] [25]),
    .ZN(_21861_)
  );
  INV_X1 _29977_ (
    .A(\cpuregs[30] [26]),
    .ZN(_21862_)
  );
  INV_X1 _29978_ (
    .A(\cpuregs[30] [28]),
    .ZN(_21863_)
  );
  INV_X1 _29979_ (
    .A(\cpuregs[30] [29]),
    .ZN(_21864_)
  );
  INV_X1 _29980_ (
    .A(\cpuregs[26] [0]),
    .ZN(_21865_)
  );
  INV_X1 _29981_ (
    .A(\cpuregs[26] [1]),
    .ZN(_21866_)
  );
  INV_X1 _29982_ (
    .A(\cpuregs[26] [2]),
    .ZN(_21867_)
  );
  INV_X1 _29983_ (
    .A(\cpuregs[26] [5]),
    .ZN(_21868_)
  );
  INV_X1 _29984_ (
    .A(\cpuregs[26] [6]),
    .ZN(_21869_)
  );
  INV_X1 _29985_ (
    .A(\cpuregs[26] [7]),
    .ZN(_21870_)
  );
  INV_X1 _29986_ (
    .A(\cpuregs[26] [8]),
    .ZN(_21871_)
  );
  INV_X1 _29987_ (
    .A(\cpuregs[26] [9]),
    .ZN(_21872_)
  );
  INV_X1 _29988_ (
    .A(\cpuregs[26] [10]),
    .ZN(_21873_)
  );
  INV_X1 _29989_ (
    .A(\cpuregs[26] [11]),
    .ZN(_21874_)
  );
  INV_X1 _29990_ (
    .A(\cpuregs[26] [12]),
    .ZN(_21875_)
  );
  INV_X1 _29991_ (
    .A(\cpuregs[26] [13]),
    .ZN(_21876_)
  );
  INV_X1 _29992_ (
    .A(\cpuregs[26] [15]),
    .ZN(_21877_)
  );
  INV_X1 _29993_ (
    .A(\cpuregs[26] [16]),
    .ZN(_21878_)
  );
  INV_X1 _29994_ (
    .A(\cpuregs[26] [17]),
    .ZN(_21879_)
  );
  INV_X1 _29995_ (
    .A(\cpuregs[26] [19]),
    .ZN(_21880_)
  );
  INV_X1 _29996_ (
    .A(\cpuregs[26] [21]),
    .ZN(_21881_)
  );
  INV_X1 _29997_ (
    .A(\cpuregs[26] [23]),
    .ZN(_21882_)
  );
  INV_X1 _29998_ (
    .A(\cpuregs[26] [25]),
    .ZN(_21883_)
  );
  INV_X1 _29999_ (
    .A(\cpuregs[26] [26]),
    .ZN(_21884_)
  );
  INV_X1 _30000_ (
    .A(\cpuregs[26] [27]),
    .ZN(_21885_)
  );
  INV_X1 _30001_ (
    .A(\cpuregs[26] [28]),
    .ZN(_21886_)
  );
  INV_X1 _30002_ (
    .A(\cpuregs[26] [29]),
    .ZN(_21887_)
  );
  INV_X1 _30003_ (
    .A(\cpuregs[26] [30]),
    .ZN(_21888_)
  );
  INV_X1 _30004_ (
    .A(\cpuregs[29] [0]),
    .ZN(_21889_)
  );
  INV_X1 _30005_ (
    .A(\cpuregs[29] [1]),
    .ZN(_21890_)
  );
  INV_X1 _30006_ (
    .A(\cpuregs[29] [2]),
    .ZN(_21891_)
  );
  INV_X1 _30007_ (
    .A(\cpuregs[29] [5]),
    .ZN(_21892_)
  );
  INV_X1 _30008_ (
    .A(\cpuregs[29] [6]),
    .ZN(_21893_)
  );
  INV_X1 _30009_ (
    .A(\cpuregs[29] [7]),
    .ZN(_21894_)
  );
  INV_X1 _30010_ (
    .A(\cpuregs[29] [9]),
    .ZN(_21895_)
  );
  INV_X1 _30011_ (
    .A(\cpuregs[29] [13]),
    .ZN(_21896_)
  );
  INV_X1 _30012_ (
    .A(\cpuregs[29] [15]),
    .ZN(_21897_)
  );
  INV_X1 _30013_ (
    .A(\cpuregs[29] [16]),
    .ZN(_21898_)
  );
  INV_X1 _30014_ (
    .A(\cpuregs[29] [19]),
    .ZN(_21899_)
  );
  INV_X1 _30015_ (
    .A(\cpuregs[29] [23]),
    .ZN(_21900_)
  );
  INV_X1 _30016_ (
    .A(\cpuregs[29] [25]),
    .ZN(_21901_)
  );
  INV_X1 _30017_ (
    .A(\cpuregs[29] [26]),
    .ZN(_21902_)
  );
  INV_X1 _30018_ (
    .A(\cpuregs[29] [28]),
    .ZN(_21903_)
  );
  INV_X1 _30019_ (
    .A(\cpuregs[29] [29]),
    .ZN(_21904_)
  );
  INV_X1 _30020_ (
    .A(\cpuregs[28] [0]),
    .ZN(_21905_)
  );
  INV_X1 _30021_ (
    .A(\cpuregs[28] [1]),
    .ZN(_21906_)
  );
  INV_X1 _30022_ (
    .A(\cpuregs[28] [2]),
    .ZN(_21907_)
  );
  INV_X1 _30023_ (
    .A(\cpuregs[28] [5]),
    .ZN(_21908_)
  );
  INV_X1 _30024_ (
    .A(\cpuregs[28] [6]),
    .ZN(_21909_)
  );
  INV_X1 _30025_ (
    .A(\cpuregs[28] [7]),
    .ZN(_21910_)
  );
  INV_X1 _30026_ (
    .A(\cpuregs[28] [9]),
    .ZN(_21911_)
  );
  INV_X1 _30027_ (
    .A(\cpuregs[28] [13]),
    .ZN(_21912_)
  );
  INV_X1 _30028_ (
    .A(\cpuregs[28] [15]),
    .ZN(_21913_)
  );
  INV_X1 _30029_ (
    .A(\cpuregs[28] [16]),
    .ZN(_21914_)
  );
  INV_X1 _30030_ (
    .A(\cpuregs[28] [19]),
    .ZN(_21915_)
  );
  INV_X1 _30031_ (
    .A(\cpuregs[28] [23]),
    .ZN(_21916_)
  );
  INV_X1 _30032_ (
    .A(\cpuregs[28] [25]),
    .ZN(_21917_)
  );
  INV_X1 _30033_ (
    .A(\cpuregs[28] [26]),
    .ZN(_21918_)
  );
  INV_X1 _30034_ (
    .A(\cpuregs[28] [28]),
    .ZN(_21919_)
  );
  INV_X1 _30035_ (
    .A(\cpuregs[28] [29]),
    .ZN(_21920_)
  );
  INV_X1 _30036_ (
    .A(\cpuregs[27] [0]),
    .ZN(_21921_)
  );
  INV_X1 _30037_ (
    .A(\cpuregs[27] [1]),
    .ZN(_21922_)
  );
  INV_X1 _30038_ (
    .A(\cpuregs[27] [2]),
    .ZN(_21923_)
  );
  INV_X1 _30039_ (
    .A(\cpuregs[27] [5]),
    .ZN(_21924_)
  );
  INV_X1 _30040_ (
    .A(\cpuregs[27] [6]),
    .ZN(_21925_)
  );
  INV_X1 _30041_ (
    .A(\cpuregs[27] [7]),
    .ZN(_21926_)
  );
  INV_X1 _30042_ (
    .A(\cpuregs[27] [9]),
    .ZN(_21927_)
  );
  INV_X1 _30043_ (
    .A(\cpuregs[27] [13]),
    .ZN(_21928_)
  );
  INV_X1 _30044_ (
    .A(\cpuregs[27] [15]),
    .ZN(_21929_)
  );
  INV_X1 _30045_ (
    .A(\cpuregs[27] [16]),
    .ZN(_21930_)
  );
  INV_X1 _30046_ (
    .A(\cpuregs[27] [19]),
    .ZN(_21931_)
  );
  INV_X1 _30047_ (
    .A(\cpuregs[27] [23]),
    .ZN(_21932_)
  );
  INV_X1 _30048_ (
    .A(\cpuregs[27] [25]),
    .ZN(_21933_)
  );
  INV_X1 _30049_ (
    .A(\cpuregs[27] [26]),
    .ZN(_21934_)
  );
  INV_X1 _30050_ (
    .A(\cpuregs[27] [28]),
    .ZN(_21935_)
  );
  INV_X1 _30051_ (
    .A(\cpuregs[27] [29]),
    .ZN(_21936_)
  );
  INV_X1 _30052_ (
    .A(\cpuregs[31] [0]),
    .ZN(_21937_)
  );
  INV_X1 _30053_ (
    .A(\cpuregs[31] [1]),
    .ZN(_21938_)
  );
  INV_X1 _30054_ (
    .A(\cpuregs[31] [2]),
    .ZN(_21939_)
  );
  INV_X1 _30055_ (
    .A(\cpuregs[31] [5]),
    .ZN(_21940_)
  );
  INV_X1 _30056_ (
    .A(\cpuregs[31] [6]),
    .ZN(_21941_)
  );
  INV_X1 _30057_ (
    .A(\cpuregs[31] [7]),
    .ZN(_21942_)
  );
  INV_X1 _30058_ (
    .A(\cpuregs[31] [9]),
    .ZN(_21943_)
  );
  INV_X1 _30059_ (
    .A(\cpuregs[31] [13]),
    .ZN(_21944_)
  );
  INV_X1 _30060_ (
    .A(\cpuregs[31] [15]),
    .ZN(_21945_)
  );
  INV_X1 _30061_ (
    .A(\cpuregs[31] [16]),
    .ZN(_21946_)
  );
  INV_X1 _30062_ (
    .A(\cpuregs[31] [19]),
    .ZN(_21947_)
  );
  INV_X1 _30063_ (
    .A(\cpuregs[31] [23]),
    .ZN(_21948_)
  );
  INV_X1 _30064_ (
    .A(\cpuregs[31] [25]),
    .ZN(_21949_)
  );
  INV_X1 _30065_ (
    .A(\cpuregs[31] [26]),
    .ZN(_21950_)
  );
  INV_X1 _30066_ (
    .A(\cpuregs[31] [28]),
    .ZN(_21951_)
  );
  INV_X1 _30067_ (
    .A(\cpuregs[31] [29]),
    .ZN(_21952_)
  );
  INV_X1 _30068_ (
    .A(\cpuregs[0] [0]),
    .ZN(_21953_)
  );
  INV_X1 _30069_ (
    .A(\cpuregs[0] [1]),
    .ZN(_21954_)
  );
  INV_X1 _30070_ (
    .A(\cpuregs[0] [2]),
    .ZN(_21955_)
  );
  INV_X1 _30071_ (
    .A(\cpuregs[0] [3]),
    .ZN(_21956_)
  );
  INV_X1 _30072_ (
    .A(\cpuregs[0] [4]),
    .ZN(_21957_)
  );
  INV_X1 _30073_ (
    .A(\cpuregs[0] [5]),
    .ZN(_21958_)
  );
  INV_X1 _30074_ (
    .A(\cpuregs[0] [6]),
    .ZN(_21959_)
  );
  INV_X1 _30075_ (
    .A(\cpuregs[0] [7]),
    .ZN(_21960_)
  );
  INV_X1 _30076_ (
    .A(\cpuregs[0] [8]),
    .ZN(_21961_)
  );
  INV_X1 _30077_ (
    .A(\cpuregs[0] [11]),
    .ZN(_21962_)
  );
  INV_X1 _30078_ (
    .A(\cpuregs[0] [13]),
    .ZN(_21963_)
  );
  INV_X1 _30079_ (
    .A(\cpuregs[0] [14]),
    .ZN(_21964_)
  );
  INV_X1 _30080_ (
    .A(\cpuregs[0] [15]),
    .ZN(_21965_)
  );
  INV_X1 _30081_ (
    .A(\cpuregs[0] [16]),
    .ZN(_21966_)
  );
  INV_X1 _30082_ (
    .A(\cpuregs[0] [17]),
    .ZN(_21967_)
  );
  INV_X1 _30083_ (
    .A(\cpuregs[0] [18]),
    .ZN(_21968_)
  );
  INV_X1 _30084_ (
    .A(\cpuregs[0] [19]),
    .ZN(_21969_)
  );
  INV_X1 _30085_ (
    .A(\cpuregs[0] [21]),
    .ZN(_21970_)
  );
  INV_X1 _30086_ (
    .A(\cpuregs[0] [23]),
    .ZN(_21971_)
  );
  INV_X1 _30087_ (
    .A(\cpuregs[0] [25]),
    .ZN(_21972_)
  );
  INV_X1 _30088_ (
    .A(\cpuregs[0] [26]),
    .ZN(_21973_)
  );
  INV_X1 _30089_ (
    .A(\cpuregs[0] [27]),
    .ZN(_21974_)
  );
  INV_X1 _30090_ (
    .A(\cpuregs[0] [28]),
    .ZN(_21975_)
  );
  INV_X1 _30091_ (
    .A(\cpuregs[0] [29]),
    .ZN(_21976_)
  );
  INV_X1 _30092_ (
    .A(\cpuregs[0] [30]),
    .ZN(_21977_)
  );
  INV_X1 _30093_ (
    .A(decoded_imm[31]),
    .ZN(_21978_)
  );
  INV_X1 _30094_ (
    .A(decoded_imm[30]),
    .ZN(_21979_)
  );
  INV_X1 _30095_ (
    .A(decoded_imm[29]),
    .ZN(_21980_)
  );
  INV_X1 _30096_ (
    .A(decoded_imm[28]),
    .ZN(_21981_)
  );
  INV_X1 _30097_ (
    .A(decoded_imm[27]),
    .ZN(_21982_)
  );
  INV_X1 _30098_ (
    .A(decoded_imm[26]),
    .ZN(_21983_)
  );
  INV_X1 _30099_ (
    .A(decoded_imm[25]),
    .ZN(_21984_)
  );
  INV_X1 _30100_ (
    .A(decoded_imm[24]),
    .ZN(_21985_)
  );
  INV_X1 _30101_ (
    .A(decoded_imm[23]),
    .ZN(_21986_)
  );
  INV_X1 _30102_ (
    .A(decoded_imm[22]),
    .ZN(_21987_)
  );
  INV_X1 _30103_ (
    .A(decoded_imm[21]),
    .ZN(_21988_)
  );
  INV_X1 _30104_ (
    .A(decoded_imm[20]),
    .ZN(_21989_)
  );
  INV_X1 _30105_ (
    .A(decoded_imm[19]),
    .ZN(_21990_)
  );
  INV_X1 _30106_ (
    .A(decoded_imm[18]),
    .ZN(_21991_)
  );
  INV_X1 _30107_ (
    .A(decoded_imm[17]),
    .ZN(_21992_)
  );
  INV_X1 _30108_ (
    .A(decoded_imm[16]),
    .ZN(_21993_)
  );
  INV_X1 _30109_ (
    .A(decoded_imm[15]),
    .ZN(_21994_)
  );
  INV_X1 _30110_ (
    .A(decoded_imm[14]),
    .ZN(_21995_)
  );
  INV_X1 _30111_ (
    .A(decoded_imm[13]),
    .ZN(_21996_)
  );
  INV_X1 _30112_ (
    .A(decoded_imm[12]),
    .ZN(_21997_)
  );
  INV_X1 _30113_ (
    .A(decoded_imm[11]),
    .ZN(_21998_)
  );
  INV_X1 _30114_ (
    .A(decoded_imm[10]),
    .ZN(_21999_)
  );
  INV_X1 _30115_ (
    .A(decoded_imm[9]),
    .ZN(_22000_)
  );
  INV_X1 _30116_ (
    .A(decoded_imm[8]),
    .ZN(_22001_)
  );
  INV_X1 _30117_ (
    .A(decoded_imm[7]),
    .ZN(_22002_)
  );
  INV_X1 _30118_ (
    .A(decoded_imm[6]),
    .ZN(_22003_)
  );
  INV_X1 _30119_ (
    .A(decoded_imm[5]),
    .ZN(_22004_)
  );
  INV_X1 _30120_ (
    .A(decoded_imm[4]),
    .ZN(_22005_)
  );
  INV_X1 _30121_ (
    .A(decoded_imm[3]),
    .ZN(_22006_)
  );
  INV_X1 _30122_ (
    .A(decoded_imm[2]),
    .ZN(_22007_)
  );
  INV_X1 _30123_ (
    .A(decoded_imm[1]),
    .ZN(_22008_)
  );
  INV_X1 _30124_ (
    .A(decoded_imm_j[7]),
    .ZN(_22009_)
  );
  INV_X1 _30125_ (
    .A(decoded_imm_j[6]),
    .ZN(_22010_)
  );
  INV_X1 _30126_ (
    .A(decoded_imm_j[5]),
    .ZN(_22011_)
  );
  INV_X1 _30127_ (
    .A(decoded_imm_j[8]),
    .ZN(_22012_)
  );
  INV_X1 _30128_ (
    .A(decoded_imm_j[9]),
    .ZN(_22013_)
  );
  INV_X1 _30129_ (
    .A(decoded_imm_j[30]),
    .ZN(_22014_)
  );
  INV_X1 _30130_ (
    .A(decoded_imm_j[4]),
    .ZN(_22015_)
  );
  INV_X1 _30131_ (
    .A(decoded_imm_j[12]),
    .ZN(_22016_)
  );
  INV_X1 _30132_ (
    .A(decoded_imm_j[13]),
    .ZN(_22017_)
  );
  INV_X1 _30133_ (
    .A(decoded_imm_j[14]),
    .ZN(_22018_)
  );
  INV_X1 _30134_ (
    .A(decoded_imm_j[18]),
    .ZN(_22019_)
  );
  INV_X1 _30135_ (
    .A(decoded_imm_j[19]),
    .ZN(_22020_)
  );
  INV_X1 _30136_ (
    .A(decoded_rs1[0]),
    .ZN(_22021_)
  );
  INV_X1 _30137_ (
    .A(decoded_rs1[1]),
    .ZN(_22022_)
  );
  INV_X1 _30138_ (
    .A(decoded_rs1[2]),
    .ZN(_22023_)
  );
  INV_X1 _30139_ (
    .A(reg_op1[1]),
    .ZN(_22024_)
  );
  INV_X1 _30140_ (
    .A(cpu_state[6]),
    .ZN(_22025_)
  );
  INV_X1 _30141_ (
    .A(cpu_state[5]),
    .ZN(_22026_)
  );
  INV_X1 _30142_ (
    .A(cpu_state[4]),
    .ZN(_22027_)
  );
  INV_X1 _30143_ (
    .A(reg_sh[4]),
    .ZN(_22028_)
  );
  INV_X1 _30144_ (
    .A(reg_sh[3]),
    .ZN(_22029_)
  );
  INV_X1 _30145_ (
    .A(reg_sh[1]),
    .ZN(_22030_)
  );
  INV_X1 _30146_ (
    .A(cpu_state[2]),
    .ZN(_22031_)
  );
  INV_X1 _30147_ (
    .A(cpu_state[1]),
    .ZN(_22032_)
  );
  INV_X1 _30148_ (
    .A(cpu_state[3]),
    .ZN(_22033_)
  );
  INV_X1 _30149_ (
    .A(cpu_state[0]),
    .ZN(_22034_)
  );
  INV_X1 _30150_ (
    .A(cpu_state[7]),
    .ZN(_22035_)
  );
  INV_X1 _30151_ (
    .A(reg_sh[0]),
    .ZN(_22036_)
  );
  INV_X1 _30152_ (
    .A(reg_sh[2]),
    .ZN(_22037_)
  );
  INV_X1 _30153_ (
    .A(_00039_),
    .ZN(_22038_)
  );
  INV_X1 _30154_ (
    .A(_00038_),
    .ZN(_22039_)
  );
  INV_X1 _30155_ (
    .A(_00037_),
    .ZN(_22040_)
  );
  INV_X1 _30156_ (
    .A(_00036_),
    .ZN(_22041_)
  );
  INV_X1 _30157_ (
    .A(_00020_),
    .ZN(_22042_)
  );
  INV_X1 _30158_ (
    .A(_00019_),
    .ZN(_22043_)
  );
  INV_X1 _30159_ (
    .A(_00018_),
    .ZN(_22044_)
  );
  INV_X1 _30160_ (
    .A(_00024_),
    .ZN(_22045_)
  );
  INV_X1 _30161_ (
    .A(_00023_),
    .ZN(_22046_)
  );
  INV_X1 _30162_ (
    .A(_00022_),
    .ZN(_22047_)
  );
  INV_X1 _30163_ (
    .A(_00021_),
    .ZN(_22048_)
  );
  INV_X1 _30164_ (
    .A(_00045_),
    .ZN(_22049_)
  );
  INV_X1 _30165_ (
    .A(_00041_),
    .ZN(_22050_)
  );
  INV_X1 _30166_ (
    .A(_00043_),
    .ZN(_22051_)
  );
  INV_X1 _30167_ (
    .A(_00042_),
    .ZN(_22052_)
  );
  INV_X1 _30168_ (
    .A(_00009_),
    .ZN(_22053_)
  );
  INV_X1 _30169_ (
    .A(_00013_),
    .ZN(_22054_)
  );
  INV_X1 _30170_ (
    .A(_00016_),
    .ZN(_22055_)
  );
  INV_X1 _30171_ (
    .A(_00015_),
    .ZN(_22056_)
  );
  INV_X1 _30172_ (
    .A(_00014_),
    .ZN(_22057_)
  );
  INV_X1 _30173_ (
    .A(_00011_),
    .ZN(_22058_)
  );
  INV_X1 _30174_ (
    .A(_00010_),
    .ZN(_22059_)
  );
  INV_X1 _30175_ (
    .A(_00012_),
    .ZN(_22060_)
  );
  INV_X1 _30176_ (
    .A(_00026_),
    .ZN(_22061_)
  );
  INV_X1 _30177_ (
    .A(_00025_),
    .ZN(_22062_)
  );
  INV_X1 _30178_ (
    .A(_00044_),
    .ZN(_22063_)
  );
  INV_X1 _30179_ (
    .A(_29146_[1]),
    .ZN(_22064_)
  );
  INV_X1 _30180_ (
    .A(_00032_),
    .ZN(_22065_)
  );
  INV_X1 _30181_ (
    .A(_00031_),
    .ZN(_22066_)
  );
  INV_X1 _30182_ (
    .A(decoder_trigger),
    .ZN(_22067_)
  );
  INV_X1 _30183_ (
    .A(_29149_[1]),
    .ZN(_22068_)
  );
  INV_X1 _30184_ (
    .A(_29149_[4]),
    .ZN(_22069_)
  );
  INV_X1 _30185_ (
    .A(is_lui_auipc_jal),
    .ZN(_22070_)
  );
  INV_X1 _30186_ (
    .A(_00034_),
    .ZN(_22071_)
  );
  INV_X1 _30187_ (
    .A(_00047_),
    .ZN(_22072_)
  );
  INV_X1 _30188_ (
    .A(_00046_),
    .ZN(_22073_)
  );
  INV_X1 _30189_ (
    .A(_00035_),
    .ZN(_22074_)
  );
  INV_X1 _30190_ (
    .A(mem_ready),
    .ZN(_22075_)
  );
  INV_X1 _30191_ (
    .A(trap),
    .ZN(_22076_)
  );
  INV_X1 _30192_ (
    .A(_00007_[2]),
    .ZN(_22077_)
  );
  INV_X1 _30193_ (
    .A(_00007_[1]),
    .ZN(_22078_)
  );
  INV_X1 _30194_ (
    .A(reg_out[2]),
    .ZN(_22079_)
  );
  INV_X1 _30195_ (
    .A(reg_out[3]),
    .ZN(_22080_)
  );
  INV_X1 _30196_ (
    .A(reg_out[4]),
    .ZN(_22081_)
  );
  INV_X1 _30197_ (
    .A(reg_out[5]),
    .ZN(_22082_)
  );
  INV_X1 _30198_ (
    .A(reg_out[6]),
    .ZN(_22083_)
  );
  INV_X1 _30199_ (
    .A(reg_out[7]),
    .ZN(_22084_)
  );
  INV_X1 _30200_ (
    .A(reg_out[8]),
    .ZN(_22085_)
  );
  INV_X1 _30201_ (
    .A(reg_out[9]),
    .ZN(_22086_)
  );
  INV_X1 _30202_ (
    .A(reg_out[10]),
    .ZN(_22087_)
  );
  INV_X1 _30203_ (
    .A(reg_out[11]),
    .ZN(_22088_)
  );
  INV_X1 _30204_ (
    .A(reg_out[12]),
    .ZN(_22089_)
  );
  INV_X1 _30205_ (
    .A(reg_out[13]),
    .ZN(_22090_)
  );
  INV_X1 _30206_ (
    .A(reg_out[14]),
    .ZN(_22091_)
  );
  INV_X1 _30207_ (
    .A(reg_out[15]),
    .ZN(_22092_)
  );
  INV_X1 _30208_ (
    .A(reg_out[16]),
    .ZN(_22093_)
  );
  INV_X1 _30209_ (
    .A(reg_out[17]),
    .ZN(_22094_)
  );
  INV_X1 _30210_ (
    .A(reg_out[18]),
    .ZN(_22095_)
  );
  INV_X1 _30211_ (
    .A(reg_out[19]),
    .ZN(_22096_)
  );
  INV_X1 _30212_ (
    .A(reg_out[20]),
    .ZN(_22097_)
  );
  INV_X1 _30213_ (
    .A(reg_out[21]),
    .ZN(_22098_)
  );
  INV_X1 _30214_ (
    .A(reg_out[22]),
    .ZN(_22099_)
  );
  INV_X1 _30215_ (
    .A(reg_out[23]),
    .ZN(_22100_)
  );
  INV_X1 _30216_ (
    .A(reg_out[24]),
    .ZN(_22101_)
  );
  INV_X1 _30217_ (
    .A(reg_out[25]),
    .ZN(_22102_)
  );
  INV_X1 _30218_ (
    .A(reg_out[26]),
    .ZN(_22103_)
  );
  INV_X1 _30219_ (
    .A(reg_out[27]),
    .ZN(_22104_)
  );
  INV_X1 _30220_ (
    .A(reg_out[28]),
    .ZN(_22105_)
  );
  INV_X1 _30221_ (
    .A(reg_out[29]),
    .ZN(_22106_)
  );
  INV_X1 _30222_ (
    .A(reg_out[30]),
    .ZN(_22107_)
  );
  INV_X1 _30223_ (
    .A(reg_out[31]),
    .ZN(_22108_)
  );
  INV_X1 _30224_ (
    .A(_00007_[3]),
    .ZN(_22109_)
  );
  INV_X1 _30225_ (
    .A(reg_out[0]),
    .ZN(_22110_)
  );
  INV_X1 _30226_ (
    .A(alu_out_q[0]),
    .ZN(_22111_)
  );
  INV_X1 _30227_ (
    .A(reg_out[1]),
    .ZN(_22112_)
  );
  INV_X1 _30228_ (
    .A(alu_out_q[1]),
    .ZN(_22113_)
  );
  INV_X1 _30229_ (
    .A(alu_out_q[2]),
    .ZN(_22114_)
  );
  INV_X1 _30230_ (
    .A(alu_out_q[3]),
    .ZN(_22115_)
  );
  INV_X1 _30231_ (
    .A(alu_out_q[4]),
    .ZN(_22116_)
  );
  INV_X1 _30232_ (
    .A(alu_out_q[5]),
    .ZN(_22117_)
  );
  INV_X1 _30233_ (
    .A(alu_out_q[6]),
    .ZN(_22118_)
  );
  INV_X1 _30234_ (
    .A(alu_out_q[7]),
    .ZN(_22119_)
  );
  INV_X1 _30235_ (
    .A(alu_out_q[8]),
    .ZN(_22120_)
  );
  INV_X1 _30236_ (
    .A(alu_out_q[9]),
    .ZN(_22121_)
  );
  INV_X1 _30237_ (
    .A(alu_out_q[10]),
    .ZN(_22122_)
  );
  INV_X1 _30238_ (
    .A(alu_out_q[11]),
    .ZN(_22123_)
  );
  INV_X1 _30239_ (
    .A(alu_out_q[12]),
    .ZN(_22124_)
  );
  INV_X1 _30240_ (
    .A(alu_out_q[13]),
    .ZN(_22125_)
  );
  INV_X1 _30241_ (
    .A(alu_out_q[14]),
    .ZN(_22126_)
  );
  INV_X1 _30242_ (
    .A(alu_out_q[15]),
    .ZN(_22127_)
  );
  INV_X1 _30243_ (
    .A(alu_out_q[16]),
    .ZN(_22128_)
  );
  INV_X1 _30244_ (
    .A(alu_out_q[17]),
    .ZN(_22129_)
  );
  INV_X1 _30245_ (
    .A(alu_out_q[18]),
    .ZN(_22130_)
  );
  INV_X1 _30246_ (
    .A(alu_out_q[19]),
    .ZN(_22131_)
  );
  INV_X1 _30247_ (
    .A(alu_out_q[20]),
    .ZN(_22132_)
  );
  INV_X1 _30248_ (
    .A(alu_out_q[21]),
    .ZN(_22133_)
  );
  INV_X1 _30249_ (
    .A(alu_out_q[22]),
    .ZN(_22134_)
  );
  INV_X1 _30250_ (
    .A(alu_out_q[23]),
    .ZN(_22135_)
  );
  INV_X1 _30251_ (
    .A(alu_out_q[24]),
    .ZN(_22136_)
  );
  INV_X1 _30252_ (
    .A(alu_out_q[25]),
    .ZN(_22137_)
  );
  INV_X1 _30253_ (
    .A(alu_out_q[26]),
    .ZN(_22138_)
  );
  INV_X1 _30254_ (
    .A(alu_out_q[27]),
    .ZN(_22139_)
  );
  INV_X1 _30255_ (
    .A(alu_out_q[28]),
    .ZN(_22140_)
  );
  INV_X1 _30256_ (
    .A(alu_out_q[29]),
    .ZN(_22141_)
  );
  INV_X1 _30257_ (
    .A(alu_out_q[30]),
    .ZN(_22142_)
  );
  INV_X1 _30258_ (
    .A(alu_out_q[31]),
    .ZN(_22143_)
  );
  INV_X1 _30259_ (
    .A(_00007_[4]),
    .ZN(_22144_)
  );
  INV_X1 _30260_ (
    .A(_29150_[2]),
    .ZN(_22145_)
  );
  INV_X1 _30261_ (
    .A(_00033_),
    .ZN(_22146_)
  );
  INV_X1 _30262_ (
    .A(_00008_[0]),
    .ZN(_22147_)
  );
  INV_X1 _30263_ (
    .A(_00008_[1]),
    .ZN(_22148_)
  );
  INV_X1 _30264_ (
    .A(_00008_[2]),
    .ZN(_22149_)
  );
  INV_X1 _30265_ (
    .A(_00008_[3]),
    .ZN(_22150_)
  );
  INV_X1 _30266_ (
    .A(_00008_[4]),
    .ZN(_22151_)
  );
  INV_X1 _30267_ (
    .A(_00007_[0]),
    .ZN(_22152_)
  );
  INV_X1 _30268_ (
    .A(count_cycle[0]),
    .ZN(_22153_)
  );
  INV_X1 _30269_ (
    .A(count_cycle[1]),
    .ZN(_22154_)
  );
  INV_X1 _30270_ (
    .A(count_cycle[2]),
    .ZN(_22155_)
  );
  INV_X1 _30271_ (
    .A(count_cycle[3]),
    .ZN(_22156_)
  );
  INV_X1 _30272_ (
    .A(count_cycle[4]),
    .ZN(_22157_)
  );
  INV_X1 _30273_ (
    .A(count_cycle[5]),
    .ZN(_22158_)
  );
  INV_X1 _30274_ (
    .A(count_cycle[6]),
    .ZN(_22159_)
  );
  INV_X1 _30275_ (
    .A(count_cycle[7]),
    .ZN(_22160_)
  );
  INV_X1 _30276_ (
    .A(count_cycle[8]),
    .ZN(_22161_)
  );
  INV_X1 _30277_ (
    .A(count_cycle[9]),
    .ZN(_22162_)
  );
  INV_X1 _30278_ (
    .A(count_cycle[10]),
    .ZN(_22163_)
  );
  INV_X1 _30279_ (
    .A(count_cycle[11]),
    .ZN(_22164_)
  );
  INV_X1 _30280_ (
    .A(count_cycle[12]),
    .ZN(_22165_)
  );
  INV_X1 _30281_ (
    .A(count_cycle[13]),
    .ZN(_22166_)
  );
  INV_X1 _30282_ (
    .A(count_cycle[14]),
    .ZN(_22167_)
  );
  INV_X1 _30283_ (
    .A(count_cycle[15]),
    .ZN(_22168_)
  );
  INV_X1 _30284_ (
    .A(count_cycle[16]),
    .ZN(_22169_)
  );
  INV_X1 _30285_ (
    .A(count_cycle[17]),
    .ZN(_22170_)
  );
  INV_X1 _30286_ (
    .A(count_cycle[18]),
    .ZN(_22171_)
  );
  INV_X1 _30287_ (
    .A(count_cycle[19]),
    .ZN(_22172_)
  );
  INV_X1 _30288_ (
    .A(count_cycle[20]),
    .ZN(_22173_)
  );
  INV_X1 _30289_ (
    .A(count_cycle[21]),
    .ZN(_22174_)
  );
  INV_X1 _30290_ (
    .A(count_cycle[22]),
    .ZN(_22175_)
  );
  INV_X1 _30291_ (
    .A(count_cycle[23]),
    .ZN(_22176_)
  );
  INV_X1 _30292_ (
    .A(count_cycle[24]),
    .ZN(_22177_)
  );
  INV_X1 _30293_ (
    .A(count_cycle[25]),
    .ZN(_22178_)
  );
  INV_X1 _30294_ (
    .A(count_cycle[26]),
    .ZN(_22179_)
  );
  INV_X1 _30295_ (
    .A(count_cycle[27]),
    .ZN(_22180_)
  );
  INV_X1 _30296_ (
    .A(count_cycle[28]),
    .ZN(_22181_)
  );
  INV_X1 _30297_ (
    .A(count_cycle[29]),
    .ZN(_22182_)
  );
  INV_X1 _30298_ (
    .A(count_cycle[30]),
    .ZN(_22183_)
  );
  INV_X1 _30299_ (
    .A(count_cycle[31]),
    .ZN(_22184_)
  );
  INV_X1 _30300_ (
    .A(count_cycle[32]),
    .ZN(_22185_)
  );
  INV_X1 _30301_ (
    .A(count_cycle[33]),
    .ZN(_22186_)
  );
  INV_X1 _30302_ (
    .A(count_cycle[34]),
    .ZN(_22187_)
  );
  INV_X1 _30303_ (
    .A(count_cycle[35]),
    .ZN(_22188_)
  );
  INV_X1 _30304_ (
    .A(count_cycle[36]),
    .ZN(_22189_)
  );
  INV_X1 _30305_ (
    .A(count_cycle[37]),
    .ZN(_22190_)
  );
  INV_X1 _30306_ (
    .A(count_cycle[38]),
    .ZN(_22191_)
  );
  INV_X1 _30307_ (
    .A(count_cycle[39]),
    .ZN(_22192_)
  );
  INV_X1 _30308_ (
    .A(count_cycle[40]),
    .ZN(_22193_)
  );
  INV_X1 _30309_ (
    .A(count_cycle[41]),
    .ZN(_22194_)
  );
  INV_X1 _30310_ (
    .A(count_cycle[42]),
    .ZN(_22195_)
  );
  INV_X1 _30311_ (
    .A(count_cycle[43]),
    .ZN(_22196_)
  );
  INV_X1 _30312_ (
    .A(count_cycle[44]),
    .ZN(_22197_)
  );
  INV_X1 _30313_ (
    .A(count_cycle[45]),
    .ZN(_22198_)
  );
  INV_X1 _30314_ (
    .A(count_cycle[46]),
    .ZN(_22199_)
  );
  INV_X1 _30315_ (
    .A(count_cycle[47]),
    .ZN(_22200_)
  );
  INV_X1 _30316_ (
    .A(count_cycle[48]),
    .ZN(_22201_)
  );
  INV_X1 _30317_ (
    .A(count_cycle[49]),
    .ZN(_22202_)
  );
  INV_X1 _30318_ (
    .A(count_cycle[50]),
    .ZN(_22203_)
  );
  INV_X1 _30319_ (
    .A(count_cycle[51]),
    .ZN(_22204_)
  );
  INV_X1 _30320_ (
    .A(count_cycle[52]),
    .ZN(_22205_)
  );
  INV_X1 _30321_ (
    .A(count_cycle[53]),
    .ZN(_22206_)
  );
  INV_X1 _30322_ (
    .A(count_cycle[54]),
    .ZN(_22207_)
  );
  INV_X1 _30323_ (
    .A(count_cycle[55]),
    .ZN(_22208_)
  );
  INV_X1 _30324_ (
    .A(count_cycle[56]),
    .ZN(_22209_)
  );
  INV_X1 _30325_ (
    .A(count_cycle[57]),
    .ZN(_22210_)
  );
  INV_X1 _30326_ (
    .A(count_cycle[58]),
    .ZN(_22211_)
  );
  INV_X1 _30327_ (
    .A(count_cycle[59]),
    .ZN(_22212_)
  );
  INV_X1 _30328_ (
    .A(count_cycle[60]),
    .ZN(_22213_)
  );
  INV_X1 _30329_ (
    .A(count_cycle[61]),
    .ZN(_22214_)
  );
  INV_X1 _30330_ (
    .A(count_cycle[62]),
    .ZN(_22215_)
  );
  INV_X1 _30331_ (
    .A(count_cycle[63]),
    .ZN(_22216_)
  );
  INV_X1 _30332_ (
    .A(_29149_[3]),
    .ZN(_22217_)
  );
  INV_X1 _30333_ (
    .A(_29151_[28]),
    .ZN(_22218_)
  );
  INV_X1 _30334_ (
    .A(_29151_[29]),
    .ZN(_22219_)
  );
  INV_X1 _30335_ (
    .A(_29151_[9]),
    .ZN(_22220_)
  );
  INV_X1 _30336_ (
    .A(_29151_[10]),
    .ZN(_22221_)
  );
  INV_X1 _30337_ (
    .A(_29151_[11]),
    .ZN(_22222_)
  );
  INV_X1 _30338_ (
    .A(_29151_[14]),
    .ZN(_22223_)
  );
  INV_X1 _30339_ (
    .A(_29151_[15]),
    .ZN(_22224_)
  );
  INV_X1 _30340_ (
    .A(_29151_[16]),
    .ZN(_22225_)
  );
  INV_X1 _30341_ (
    .A(_29151_[18]),
    .ZN(_22226_)
  );
  INV_X1 _30342_ (
    .A(_29151_[19]),
    .ZN(_22227_)
  );
  INV_X1 _30343_ (
    .A(_29151_[20]),
    .ZN(_22228_)
  );
  INV_X1 _30344_ (
    .A(_29151_[23]),
    .ZN(_22229_)
  );
  INV_X1 _30345_ (
    .A(_29151_[25]),
    .ZN(_22230_)
  );
  INV_X1 _30346_ (
    .A(_29151_[30]),
    .ZN(_22231_)
  );
  INV_X1 _30347_ (
    .A(_29151_[0]),
    .ZN(_22232_)
  );
  INV_X1 _30348_ (
    .A(_29151_[1]),
    .ZN(_22233_)
  );
  INV_X1 _30349_ (
    .A(_29151_[2]),
    .ZN(_22234_)
  );
  INV_X1 _30350_ (
    .A(_29151_[3]),
    .ZN(_22235_)
  );
  INV_X1 _30351_ (
    .A(_29151_[4]),
    .ZN(_22236_)
  );
  INV_X1 _30352_ (
    .A(_29151_[5]),
    .ZN(_22237_)
  );
  INV_X1 _30353_ (
    .A(_29151_[6]),
    .ZN(_22238_)
  );
  INV_X1 _30354_ (
    .A(_29151_[17]),
    .ZN(_22239_)
  );
  INV_X1 _30355_ (
    .A(_29151_[24]),
    .ZN(_22240_)
  );
  INV_X1 _30356_ (
    .A(_29151_[27]),
    .ZN(_22241_)
  );
  INV_X1 _30357_ (
    .A(_29151_[22]),
    .ZN(_22242_)
  );
  INV_X1 _30358_ (
    .A(_29151_[7]),
    .ZN(_22243_)
  );
  INV_X1 _30359_ (
    .A(_29151_[8]),
    .ZN(_22244_)
  );
  INV_X1 _30360_ (
    .A(_29151_[12]),
    .ZN(_22245_)
  );
  INV_X1 _30361_ (
    .A(_29151_[13]),
    .ZN(_22246_)
  );
  INV_X1 _30362_ (
    .A(_29151_[21]),
    .ZN(_22247_)
  );
  INV_X1 _30363_ (
    .A(_29151_[26]),
    .ZN(_22248_)
  );
  INV_X1 _30364_ (
    .A(_29151_[31]),
    .ZN(_22249_)
  );
  AND2_X1 _30365_ (
    .A1(_22025_),
    .A2(_22035_),
    .ZN(_22250_)
  );
  AND2_X1 _30366_ (
    .A1(_22026_),
    .A2(_22027_),
    .ZN(_22251_)
  );
  AND2_X1 _30367_ (
    .A1(_22250_),
    .A2(_22251_),
    .ZN(_22252_)
  );
  AND2_X1 _30368_ (
    .A1(_22031_),
    .A2(_22033_),
    .ZN(_22253_)
  );
  AND2_X1 _30369_ (
    .A1(_22032_),
    .A2(_22055_),
    .ZN(_22254_)
  );
  AND2_X1 _30370_ (
    .A1(_22253_),
    .A2(_22254_),
    .ZN(_22255_)
  );
  AND2_X1 _30371_ (
    .A1(_22252_),
    .A2(_22255_),
    .ZN(_22256_)
  );
  INV_X1 _30372_ (
    .A(_22256_),
    .ZN(_22257_)
  );
  AND2_X1 _30373_ (
    .A1(_22032_),
    .A2(_22034_),
    .ZN(_22258_)
  );
  AND2_X1 _30374_ (
    .A1(_22033_),
    .A2(_22057_),
    .ZN(_22259_)
  );
  AND2_X1 _30375_ (
    .A1(_22258_),
    .A2(_22259_),
    .ZN(_22260_)
  );
  AND2_X1 _30376_ (
    .A1(_22252_),
    .A2(_22260_),
    .ZN(_22261_)
  );
  INV_X1 _30377_ (
    .A(_22261_),
    .ZN(_22262_)
  );
  AND2_X1 _30378_ (
    .A1(_22257_),
    .A2(_22262_),
    .ZN(_22263_)
  );
  AND2_X1 _30379_ (
    .A1(_22034_),
    .A2(_22056_),
    .ZN(_22264_)
  );
  AND2_X1 _30380_ (
    .A1(_22253_),
    .A2(_22264_),
    .ZN(_22265_)
  );
  AND2_X1 _30381_ (
    .A1(_22252_),
    .A2(_22265_),
    .ZN(_22266_)
  );
  INV_X1 _30382_ (
    .A(_22266_),
    .ZN(_22267_)
  );
  AND2_X1 _30383_ (
    .A1(_22253_),
    .A2(_22258_),
    .ZN(_22268_)
  );
  AND2_X1 _30384_ (
    .A1(_22250_),
    .A2(_22268_),
    .ZN(_22269_)
  );
  AND2_X1 _30385_ (
    .A1(_22027_),
    .A2(_22058_),
    .ZN(_22270_)
  );
  AND2_X1 _30386_ (
    .A1(_22269_),
    .A2(_22270_),
    .ZN(_22271_)
  );
  INV_X1 _30387_ (
    .A(_22271_),
    .ZN(_22272_)
  );
  AND2_X1 _30388_ (
    .A1(_22263_),
    .A2(_22267_),
    .ZN(_22273_)
  );
  AND2_X1 _30389_ (
    .A1(_22272_),
    .A2(_22273_),
    .ZN(_22274_)
  );
  INV_X1 _30390_ (
    .A(_22274_),
    .ZN(_22275_)
  );
  AND2_X1 _30391_ (
    .A1(_22029_),
    .A2(_22037_),
    .ZN(_22276_)
  );
  INV_X1 _30392_ (
    .A(_22276_),
    .ZN(_22277_)
  );
  AND2_X1 _30393_ (
    .A1(_22028_),
    .A2(_22036_),
    .ZN(_22278_)
  );
  AND2_X1 _30394_ (
    .A1(_22030_),
    .A2(_22278_),
    .ZN(_22279_)
  );
  AND2_X1 _30395_ (
    .A1(_22276_),
    .A2(_22279_),
    .ZN(_22280_)
  );
  INV_X1 _30396_ (
    .A(_22280_),
    .ZN(_22281_)
  );
  AND2_X1 _30397_ (
    .A1(_22261_),
    .A2(_22280_),
    .ZN(_22282_)
  );
  INV_X1 _30398_ (
    .A(_22282_),
    .ZN(_22283_)
  );
  AND2_X1 _30399_ (
    .A1(_21048_),
    .A2(_21270_),
    .ZN(_22284_)
  );
  INV_X1 _30400_ (
    .A(_22284_),
    .ZN(_22285_)
  );
  AND2_X1 _30401_ (
    .A1(_21044_),
    .A2(_21271_),
    .ZN(_22286_)
  );
  AND2_X1 _30402_ (
    .A1(_21043_),
    .A2(_21272_),
    .ZN(_22287_)
  );
  INV_X1 _30403_ (
    .A(_22287_),
    .ZN(_22288_)
  );
  AND2_X1 _30404_ (
    .A1(_22286_),
    .A2(_22287_),
    .ZN(_22289_)
  );
  INV_X1 _30405_ (
    .A(_22289_),
    .ZN(_22290_)
  );
  AND2_X1 _30406_ (
    .A1(_22284_),
    .A2(_22289_),
    .ZN(_22291_)
  );
  AND2_X1 _30407_ (
    .A1(_22261_),
    .A2(_22291_),
    .ZN(_22292_)
  );
  INV_X1 _30408_ (
    .A(_22292_),
    .ZN(_22293_)
  );
  AND2_X1 _30409_ (
    .A1(_22283_),
    .A2(_22293_),
    .ZN(_22294_)
  );
  AND2_X1 _30410_ (
    .A1(_22261_),
    .A2(_22281_),
    .ZN(_22295_)
  );
  INV_X1 _30411_ (
    .A(_22295_),
    .ZN(_22296_)
  );
  AND2_X1 _30412_ (
    .A1(_22275_),
    .A2(_22294_),
    .ZN(_22297_)
  );
  AND2_X1 _30413_ (
    .A1(mem_do_rinst),
    .A2(resetn),
    .ZN(_22298_)
  );
  AND2_X1 _30414_ (
    .A1(_21038_),
    .A2(_21069_),
    .ZN(_22299_)
  );
  INV_X1 _30415_ (
    .A(_22299_),
    .ZN(_22300_)
  );
  AND2_X1 _30416_ (
    .A1(resetn),
    .A2(_22300_),
    .ZN(_22301_)
  );
  AND2_X1 _30417_ (
    .A1(mem_state[0]),
    .A2(mem_state[1]),
    .ZN(_22302_)
  );
  AND2_X1 _30418_ (
    .A1(_22298_),
    .A2(_22302_),
    .ZN(_22303_)
  );
  INV_X1 _30419_ (
    .A(_22303_),
    .ZN(_22304_)
  );
  AND2_X1 _30420_ (
    .A1(_21348_),
    .A2(_21349_),
    .ZN(_22305_)
  );
  INV_X1 _30421_ (
    .A(_22305_),
    .ZN(_22306_)
  );
  AND2_X1 _30422_ (
    .A1(mem_valid),
    .A2(mem_ready),
    .ZN(_22307_)
  );
  INV_X1 _30423_ (
    .A(_22307_),
    .ZN(_22308_)
  );
  AND2_X1 _30424_ (
    .A1(resetn),
    .A2(_22307_),
    .ZN(_22309_)
  );
  AND2_X1 _30425_ (
    .A1(_21069_),
    .A2(_21070_),
    .ZN(_22310_)
  );
  AND2_X1 _30426_ (
    .A1(_21038_),
    .A2(_22310_),
    .ZN(_22311_)
  );
  INV_X1 _30427_ (
    .A(_22311_),
    .ZN(_22312_)
  );
  AND2_X1 _30428_ (
    .A1(_22309_),
    .A2(_22312_),
    .ZN(_22313_)
  );
  AND2_X1 _30429_ (
    .A1(_22306_),
    .A2(_22313_),
    .ZN(_22314_)
  );
  INV_X1 _30430_ (
    .A(_22314_),
    .ZN(_22315_)
  );
  AND2_X1 _30431_ (
    .A1(_22304_),
    .A2(_22315_),
    .ZN(_22316_)
  );
  INV_X1 _30432_ (
    .A(_22316_),
    .ZN(_22317_)
  );
  AND2_X1 _30433_ (
    .A1(_22074_),
    .A2(_22316_),
    .ZN(_22318_)
  );
  INV_X1 _30434_ (
    .A(_22318_),
    .ZN(_22319_)
  );
  AND2_X1 _30435_ (
    .A1(_22266_),
    .A2(_22319_),
    .ZN(_22320_)
  );
  AND2_X1 _30436_ (
    .A1(_22049_),
    .A2(_22320_),
    .ZN(_22321_)
  );
  INV_X1 _30437_ (
    .A(_22321_),
    .ZN(_22322_)
  );
  AND2_X1 _30438_ (
    .A1(_22256_),
    .A2(_22319_),
    .ZN(_22323_)
  );
  AND2_X1 _30439_ (
    .A1(_22071_),
    .A2(_22323_),
    .ZN(_22324_)
  );
  INV_X1 _30440_ (
    .A(_22324_),
    .ZN(_22325_)
  );
  AND2_X1 _30441_ (
    .A1(_22257_),
    .A2(_22267_),
    .ZN(_22326_)
  );
  INV_X1 _30442_ (
    .A(_22326_),
    .ZN(_22327_)
  );
  AND2_X1 _30443_ (
    .A1(_22318_),
    .A2(_22327_),
    .ZN(_22328_)
  );
  INV_X1 _30444_ (
    .A(_22328_),
    .ZN(_22329_)
  );
  AND2_X1 _30445_ (
    .A1(resetn),
    .A2(_22329_),
    .ZN(_22330_)
  );
  AND2_X1 _30446_ (
    .A1(_22325_),
    .A2(_22330_),
    .ZN(_22331_)
  );
  AND2_X1 _30447_ (
    .A1(_22322_),
    .A2(_22331_),
    .ZN(_22332_)
  );
  AND2_X1 _30448_ (
    .A1(_22297_),
    .A2(_22332_),
    .ZN(_22333_)
  );
  INV_X1 _30449_ (
    .A(_22333_),
    .ZN(_22334_)
  );
  AND2_X1 _30450_ (
    .A1(_21259_),
    .A2(is_lui_auipc_jal),
    .ZN(_22335_)
  );
  AND2_X1 _30451_ (
    .A1(reg_next_pc[0]),
    .A2(_22335_),
    .ZN(_22336_)
  );
  INV_X1 _30452_ (
    .A(_22336_),
    .ZN(_22337_)
  );
  AND2_X1 _30453_ (
    .A1(_21436_),
    .A2(_22149_),
    .ZN(_22338_)
  );
  INV_X1 _30454_ (
    .A(_22338_),
    .ZN(_22339_)
  );
  AND2_X1 _30455_ (
    .A1(_21647_),
    .A2(_00008_[2]),
    .ZN(_22340_)
  );
  INV_X1 _30456_ (
    .A(_22340_),
    .ZN(_22341_)
  );
  AND2_X1 _30457_ (
    .A1(_22339_),
    .A2(_22341_),
    .ZN(_22342_)
  );
  AND2_X1 _30458_ (
    .A1(_22147_),
    .A2(_22342_),
    .ZN(_22343_)
  );
  INV_X1 _30459_ (
    .A(_22343_),
    .ZN(_22344_)
  );
  AND2_X1 _30460_ (
    .A1(_21757_),
    .A2(_00008_[2]),
    .ZN(_22345_)
  );
  INV_X1 _30461_ (
    .A(_22345_),
    .ZN(_22346_)
  );
  AND2_X1 _30462_ (
    .A1(_21458_),
    .A2(_22149_),
    .ZN(_22347_)
  );
  INV_X1 _30463_ (
    .A(_22347_),
    .ZN(_22348_)
  );
  AND2_X1 _30464_ (
    .A1(_00008_[0]),
    .A2(_22346_),
    .ZN(_22349_)
  );
  AND2_X1 _30465_ (
    .A1(_22348_),
    .A2(_22349_),
    .ZN(_22350_)
  );
  INV_X1 _30466_ (
    .A(_22350_),
    .ZN(_22351_)
  );
  AND2_X1 _30467_ (
    .A1(_22344_),
    .A2(_22351_),
    .ZN(_22352_)
  );
  AND2_X1 _30468_ (
    .A1(_22148_),
    .A2(_22352_),
    .ZN(_22353_)
  );
  INV_X1 _30469_ (
    .A(_22353_),
    .ZN(_22354_)
  );
  AND2_X1 _30470_ (
    .A1(_21590_),
    .A2(_22149_),
    .ZN(_22355_)
  );
  INV_X1 _30471_ (
    .A(_22355_),
    .ZN(_22356_)
  );
  AND2_X1 _30472_ (
    .A1(_21408_),
    .A2(_00008_[2]),
    .ZN(_22357_)
  );
  INV_X1 _30473_ (
    .A(_22357_),
    .ZN(_22358_)
  );
  AND2_X1 _30474_ (
    .A1(_22356_),
    .A2(_22358_),
    .ZN(_22359_)
  );
  AND2_X1 _30475_ (
    .A1(_22147_),
    .A2(_22359_),
    .ZN(_22360_)
  );
  INV_X1 _30476_ (
    .A(_22360_),
    .ZN(_22361_)
  );
  AND2_X1 _30477_ (
    .A1(_21370_),
    .A2(_00008_[2]),
    .ZN(_22362_)
  );
  INV_X1 _30478_ (
    .A(_22362_),
    .ZN(_22363_)
  );
  AND2_X1 _30479_ (
    .A1(_21616_),
    .A2(_22149_),
    .ZN(_22364_)
  );
  INV_X1 _30480_ (
    .A(_22364_),
    .ZN(_22365_)
  );
  AND2_X1 _30481_ (
    .A1(_00008_[0]),
    .A2(_22365_),
    .ZN(_22366_)
  );
  AND2_X1 _30482_ (
    .A1(_22363_),
    .A2(_22366_),
    .ZN(_22367_)
  );
  INV_X1 _30483_ (
    .A(_22367_),
    .ZN(_22368_)
  );
  AND2_X1 _30484_ (
    .A1(_22361_),
    .A2(_22368_),
    .ZN(_22369_)
  );
  AND2_X1 _30485_ (
    .A1(_00008_[1]),
    .A2(_22369_),
    .ZN(_22370_)
  );
  INV_X1 _30486_ (
    .A(_22370_),
    .ZN(_22371_)
  );
  AND2_X1 _30487_ (
    .A1(_22354_),
    .A2(_22371_),
    .ZN(_22372_)
  );
  AND2_X1 _30488_ (
    .A1(_21865_),
    .A2(_22149_),
    .ZN(_22373_)
  );
  INV_X1 _30489_ (
    .A(_22373_),
    .ZN(_22374_)
  );
  AND2_X1 _30490_ (
    .A1(_21849_),
    .A2(_00008_[2]),
    .ZN(_22375_)
  );
  INV_X1 _30491_ (
    .A(_22375_),
    .ZN(_22376_)
  );
  AND2_X1 _30492_ (
    .A1(_22374_),
    .A2(_22376_),
    .ZN(_22377_)
  );
  AND2_X1 _30493_ (
    .A1(_22147_),
    .A2(_22377_),
    .ZN(_22378_)
  );
  INV_X1 _30494_ (
    .A(_22378_),
    .ZN(_22379_)
  );
  AND2_X1 _30495_ (
    .A1(_21937_),
    .A2(_00008_[2]),
    .ZN(_22380_)
  );
  INV_X1 _30496_ (
    .A(_22380_),
    .ZN(_22381_)
  );
  AND2_X1 _30497_ (
    .A1(_21921_),
    .A2(_22149_),
    .ZN(_22382_)
  );
  INV_X1 _30498_ (
    .A(_22382_),
    .ZN(_22383_)
  );
  AND2_X1 _30499_ (
    .A1(_00008_[0]),
    .A2(_22383_),
    .ZN(_22384_)
  );
  AND2_X1 _30500_ (
    .A1(_22381_),
    .A2(_22384_),
    .ZN(_22385_)
  );
  INV_X1 _30501_ (
    .A(_22385_),
    .ZN(_22386_)
  );
  AND2_X1 _30502_ (
    .A1(_22379_),
    .A2(_22386_),
    .ZN(_22387_)
  );
  AND2_X1 _30503_ (
    .A1(_00008_[1]),
    .A2(_22387_),
    .ZN(_22388_)
  );
  INV_X1 _30504_ (
    .A(_22388_),
    .ZN(_22389_)
  );
  AND2_X1 _30505_ (
    .A1(_21889_),
    .A2(_00008_[2]),
    .ZN(_22390_)
  );
  INV_X1 _30506_ (
    .A(_22390_),
    .ZN(_22391_)
  );
  AND2_X1 _30507_ (
    .A1(_21833_),
    .A2(_22149_),
    .ZN(_22392_)
  );
  INV_X1 _30508_ (
    .A(_22392_),
    .ZN(_22393_)
  );
  AND2_X1 _30509_ (
    .A1(_00008_[0]),
    .A2(_22393_),
    .ZN(_22394_)
  );
  AND2_X1 _30510_ (
    .A1(_22391_),
    .A2(_22394_),
    .ZN(_22395_)
  );
  INV_X1 _30511_ (
    .A(_22395_),
    .ZN(_22396_)
  );
  AND2_X1 _30512_ (
    .A1(_21567_),
    .A2(_22149_),
    .ZN(_22397_)
  );
  INV_X1 _30513_ (
    .A(_22397_),
    .ZN(_22398_)
  );
  AND2_X1 _30514_ (
    .A1(_21905_),
    .A2(_00008_[2]),
    .ZN(_22399_)
  );
  INV_X1 _30515_ (
    .A(_22399_),
    .ZN(_22400_)
  );
  AND2_X1 _30516_ (
    .A1(_22398_),
    .A2(_22400_),
    .ZN(_22401_)
  );
  AND2_X1 _30517_ (
    .A1(_22147_),
    .A2(_22401_),
    .ZN(_22402_)
  );
  INV_X1 _30518_ (
    .A(_22402_),
    .ZN(_22403_)
  );
  AND2_X1 _30519_ (
    .A1(_22396_),
    .A2(_22403_),
    .ZN(_22404_)
  );
  AND2_X1 _30520_ (
    .A1(_22148_),
    .A2(_22404_),
    .ZN(_22405_)
  );
  INV_X1 _30521_ (
    .A(_22405_),
    .ZN(_22406_)
  );
  AND2_X1 _30522_ (
    .A1(_00008_[3]),
    .A2(_22389_),
    .ZN(_22407_)
  );
  AND2_X1 _30523_ (
    .A1(_22406_),
    .A2(_22407_),
    .ZN(_22408_)
  );
  INV_X1 _30524_ (
    .A(_22408_),
    .ZN(_22409_)
  );
  AND2_X1 _30525_ (
    .A1(_22150_),
    .A2(_22372_),
    .ZN(_22410_)
  );
  INV_X1 _30526_ (
    .A(_22410_),
    .ZN(_22411_)
  );
  AND2_X1 _30527_ (
    .A1(_00008_[4]),
    .A2(_22411_),
    .ZN(_22412_)
  );
  AND2_X1 _30528_ (
    .A1(_22409_),
    .A2(_22412_),
    .ZN(_22413_)
  );
  INV_X1 _30529_ (
    .A(_22413_),
    .ZN(_22414_)
  );
  AND2_X1 _30530_ (
    .A1(\cpuregs[9] [0]),
    .A2(_22149_),
    .ZN(_22415_)
  );
  INV_X1 _30531_ (
    .A(_22415_),
    .ZN(_22416_)
  );
  AND2_X1 _30532_ (
    .A1(\cpuregs[13] [0]),
    .A2(_00008_[2]),
    .ZN(_22417_)
  );
  INV_X1 _30533_ (
    .A(_22417_),
    .ZN(_22418_)
  );
  AND2_X1 _30534_ (
    .A1(_22148_),
    .A2(_22418_),
    .ZN(_22419_)
  );
  AND2_X1 _30535_ (
    .A1(_22416_),
    .A2(_22419_),
    .ZN(_22420_)
  );
  INV_X1 _30536_ (
    .A(_22420_),
    .ZN(_22421_)
  );
  AND2_X1 _30537_ (
    .A1(\cpuregs[15] [0]),
    .A2(_00008_[2]),
    .ZN(_22422_)
  );
  INV_X1 _30538_ (
    .A(_22422_),
    .ZN(_22423_)
  );
  AND2_X1 _30539_ (
    .A1(\cpuregs[11] [0]),
    .A2(_22149_),
    .ZN(_22424_)
  );
  INV_X1 _30540_ (
    .A(_22424_),
    .ZN(_22425_)
  );
  AND2_X1 _30541_ (
    .A1(_00008_[1]),
    .A2(_22425_),
    .ZN(_22426_)
  );
  AND2_X1 _30542_ (
    .A1(_22423_),
    .A2(_22426_),
    .ZN(_22427_)
  );
  INV_X1 _30543_ (
    .A(_22427_),
    .ZN(_22428_)
  );
  AND2_X1 _30544_ (
    .A1(_22421_),
    .A2(_22428_),
    .ZN(_22429_)
  );
  INV_X1 _30545_ (
    .A(_22429_),
    .ZN(_22430_)
  );
  AND2_X1 _30546_ (
    .A1(_00008_[0]),
    .A2(_22430_),
    .ZN(_22431_)
  );
  INV_X1 _30547_ (
    .A(_22431_),
    .ZN(_22432_)
  );
  AND2_X1 _30548_ (
    .A1(\cpuregs[8] [0]),
    .A2(_22149_),
    .ZN(_22433_)
  );
  INV_X1 _30549_ (
    .A(_22433_),
    .ZN(_22434_)
  );
  AND2_X1 _30550_ (
    .A1(\cpuregs[12] [0]),
    .A2(_00008_[2]),
    .ZN(_22435_)
  );
  INV_X1 _30551_ (
    .A(_22435_),
    .ZN(_22436_)
  );
  AND2_X1 _30552_ (
    .A1(_22148_),
    .A2(_22436_),
    .ZN(_22437_)
  );
  AND2_X1 _30553_ (
    .A1(_22434_),
    .A2(_22437_),
    .ZN(_22438_)
  );
  INV_X1 _30554_ (
    .A(_22438_),
    .ZN(_22439_)
  );
  AND2_X1 _30555_ (
    .A1(\cpuregs[10] [0]),
    .A2(_22149_),
    .ZN(_22440_)
  );
  INV_X1 _30556_ (
    .A(_22440_),
    .ZN(_22441_)
  );
  AND2_X1 _30557_ (
    .A1(\cpuregs[14] [0]),
    .A2(_00008_[2]),
    .ZN(_22442_)
  );
  INV_X1 _30558_ (
    .A(_22442_),
    .ZN(_22443_)
  );
  AND2_X1 _30559_ (
    .A1(_00008_[1]),
    .A2(_22443_),
    .ZN(_22444_)
  );
  AND2_X1 _30560_ (
    .A1(_22441_),
    .A2(_22444_),
    .ZN(_22445_)
  );
  INV_X1 _30561_ (
    .A(_22445_),
    .ZN(_22446_)
  );
  AND2_X1 _30562_ (
    .A1(_22439_),
    .A2(_22446_),
    .ZN(_22447_)
  );
  INV_X1 _30563_ (
    .A(_22447_),
    .ZN(_22448_)
  );
  AND2_X1 _30564_ (
    .A1(_22147_),
    .A2(_22448_),
    .ZN(_22449_)
  );
  INV_X1 _30565_ (
    .A(_22449_),
    .ZN(_22450_)
  );
  AND2_X1 _30566_ (
    .A1(_22432_),
    .A2(_22450_),
    .ZN(_22451_)
  );
  INV_X1 _30567_ (
    .A(_22451_),
    .ZN(_22452_)
  );
  AND2_X1 _30568_ (
    .A1(_00008_[3]),
    .A2(_22452_),
    .ZN(_22453_)
  );
  INV_X1 _30569_ (
    .A(_22453_),
    .ZN(_22454_)
  );
  AND2_X1 _30570_ (
    .A1(_21732_),
    .A2(_00008_[2]),
    .ZN(_22455_)
  );
  INV_X1 _30571_ (
    .A(_22455_),
    .ZN(_22456_)
  );
  AND2_X1 _30572_ (
    .A1(_21512_),
    .A2(_22149_),
    .ZN(_22457_)
  );
  INV_X1 _30573_ (
    .A(_22457_),
    .ZN(_22458_)
  );
  AND2_X1 _30574_ (
    .A1(_00008_[0]),
    .A2(_22458_),
    .ZN(_22459_)
  );
  AND2_X1 _30575_ (
    .A1(_22456_),
    .A2(_22459_),
    .ZN(_22460_)
  );
  INV_X1 _30576_ (
    .A(_22460_),
    .ZN(_22461_)
  );
  AND2_X1 _30577_ (
    .A1(_21953_),
    .A2(_22149_),
    .ZN(_22462_)
  );
  INV_X1 _30578_ (
    .A(_22462_),
    .ZN(_22463_)
  );
  AND2_X1 _30579_ (
    .A1(_21669_),
    .A2(_00008_[2]),
    .ZN(_22464_)
  );
  INV_X1 _30580_ (
    .A(_22464_),
    .ZN(_22465_)
  );
  AND2_X1 _30581_ (
    .A1(_22463_),
    .A2(_22465_),
    .ZN(_22466_)
  );
  AND2_X1 _30582_ (
    .A1(_22147_),
    .A2(_22466_),
    .ZN(_22467_)
  );
  INV_X1 _30583_ (
    .A(_22467_),
    .ZN(_22468_)
  );
  AND2_X1 _30584_ (
    .A1(_22461_),
    .A2(_22468_),
    .ZN(_22469_)
  );
  AND2_X1 _30585_ (
    .A1(_22148_),
    .A2(_22469_),
    .ZN(_22470_)
  );
  INV_X1 _30586_ (
    .A(_22470_),
    .ZN(_22471_)
  );
  AND2_X1 _30587_ (
    .A1(_21779_),
    .A2(_00008_[2]),
    .ZN(_22472_)
  );
  INV_X1 _30588_ (
    .A(_22472_),
    .ZN(_22473_)
  );
  AND2_X1 _30589_ (
    .A1(_21487_),
    .A2(_22149_),
    .ZN(_22474_)
  );
  INV_X1 _30590_ (
    .A(_22474_),
    .ZN(_22475_)
  );
  AND2_X1 _30591_ (
    .A1(_00008_[0]),
    .A2(_22475_),
    .ZN(_22476_)
  );
  AND2_X1 _30592_ (
    .A1(_22473_),
    .A2(_22476_),
    .ZN(_22477_)
  );
  INV_X1 _30593_ (
    .A(_22477_),
    .ZN(_22478_)
  );
  AND2_X1 _30594_ (
    .A1(_21537_),
    .A2(_22149_),
    .ZN(_22479_)
  );
  INV_X1 _30595_ (
    .A(_22479_),
    .ZN(_22480_)
  );
  AND2_X1 _30596_ (
    .A1(_21804_),
    .A2(_00008_[2]),
    .ZN(_22481_)
  );
  INV_X1 _30597_ (
    .A(_22481_),
    .ZN(_22482_)
  );
  AND2_X1 _30598_ (
    .A1(_22480_),
    .A2(_22482_),
    .ZN(_22483_)
  );
  AND2_X1 _30599_ (
    .A1(_22147_),
    .A2(_22483_),
    .ZN(_22484_)
  );
  INV_X1 _30600_ (
    .A(_22484_),
    .ZN(_22485_)
  );
  AND2_X1 _30601_ (
    .A1(_22478_),
    .A2(_22485_),
    .ZN(_22486_)
  );
  AND2_X1 _30602_ (
    .A1(_00008_[1]),
    .A2(_22486_),
    .ZN(_22487_)
  );
  INV_X1 _30603_ (
    .A(_22487_),
    .ZN(_22488_)
  );
  AND2_X1 _30604_ (
    .A1(_22471_),
    .A2(_22488_),
    .ZN(_22489_)
  );
  INV_X1 _30605_ (
    .A(_22489_),
    .ZN(_22490_)
  );
  AND2_X1 _30606_ (
    .A1(_22150_),
    .A2(_22490_),
    .ZN(_22491_)
  );
  INV_X1 _30607_ (
    .A(_22491_),
    .ZN(_22492_)
  );
  AND2_X1 _30608_ (
    .A1(_22454_),
    .A2(_22492_),
    .ZN(_22493_)
  );
  INV_X1 _30609_ (
    .A(_22493_),
    .ZN(_22494_)
  );
  AND2_X1 _30610_ (
    .A1(_22151_),
    .A2(_22494_),
    .ZN(_22495_)
  );
  INV_X1 _30611_ (
    .A(_22495_),
    .ZN(_22496_)
  );
  AND2_X1 _30612_ (
    .A1(_21273_),
    .A2(_21276_),
    .ZN(_22497_)
  );
  AND2_X1 _30613_ (
    .A1(_21274_),
    .A2(_21275_),
    .ZN(_22498_)
  );
  AND2_X1 _30614_ (
    .A1(_22497_),
    .A2(_22498_),
    .ZN(_22499_)
  );
  INV_X1 _30615_ (
    .A(_22499_),
    .ZN(_22500_)
  );
  AND2_X1 _30616_ (
    .A1(_21264_),
    .A2(_21269_),
    .ZN(_22501_)
  );
  AND2_X1 _30617_ (
    .A1(_21051_),
    .A2(_22501_),
    .ZN(_22502_)
  );
  AND2_X1 _30618_ (
    .A1(_22499_),
    .A2(_22502_),
    .ZN(_22503_)
  );
  AND2_X1 _30619_ (
    .A1(_21047_),
    .A2(_21055_),
    .ZN(_22504_)
  );
  AND2_X1 _30620_ (
    .A1(_21046_),
    .A2(_21054_),
    .ZN(_22505_)
  );
  AND2_X1 _30621_ (
    .A1(_22504_),
    .A2(_22505_),
    .ZN(_22506_)
  );
  AND2_X1 _30622_ (
    .A1(_21265_),
    .A2(_21267_),
    .ZN(_22507_)
  );
  AND2_X1 _30623_ (
    .A1(_21266_),
    .A2(_22507_),
    .ZN(_22508_)
  );
  INV_X1 _30624_ (
    .A(_22508_),
    .ZN(_00001_)
  );
  AND2_X1 _30625_ (
    .A1(_22506_),
    .A2(_22508_),
    .ZN(_22509_)
  );
  AND2_X1 _30626_ (
    .A1(_22503_),
    .A2(_22509_),
    .ZN(_22510_)
  );
  AND2_X1 _30627_ (
    .A1(_21040_),
    .A2(_21041_),
    .ZN(_22511_)
  );
  AND2_X1 _30628_ (
    .A1(_22284_),
    .A2(_22511_),
    .ZN(_22512_)
  );
  AND2_X1 _30629_ (
    .A1(_22289_),
    .A2(_22512_),
    .ZN(_22513_)
  );
  AND2_X1 _30630_ (
    .A1(_21060_),
    .A2(_21061_),
    .ZN(_22514_)
  );
  AND2_X1 _30631_ (
    .A1(_21062_),
    .A2(_21263_),
    .ZN(_22515_)
  );
  AND2_X1 _30632_ (
    .A1(_22514_),
    .A2(_22515_),
    .ZN(_22516_)
  );
  AND2_X1 _30633_ (
    .A1(_21056_),
    .A2(_21057_),
    .ZN(_22517_)
  );
  AND2_X1 _30634_ (
    .A1(_21058_),
    .A2(_21059_),
    .ZN(_22518_)
  );
  AND2_X1 _30635_ (
    .A1(_22517_),
    .A2(_22518_),
    .ZN(_22519_)
  );
  AND2_X1 _30636_ (
    .A1(_22516_),
    .A2(_22519_),
    .ZN(_22520_)
  );
  AND2_X1 _30637_ (
    .A1(_22513_),
    .A2(_22520_),
    .ZN(_22521_)
  );
  AND2_X1 _30638_ (
    .A1(_21259_),
    .A2(_21260_),
    .ZN(_22522_)
  );
  INV_X1 _30639_ (
    .A(_22522_),
    .ZN(_22523_)
  );
  AND2_X1 _30640_ (
    .A1(_21261_),
    .A2(_22522_),
    .ZN(_22524_)
  );
  INV_X1 _30641_ (
    .A(_22524_),
    .ZN(_00002_)
  );
  AND2_X1 _30642_ (
    .A1(_21262_),
    .A2(_22524_),
    .ZN(_22525_)
  );
  AND2_X1 _30643_ (
    .A1(_21049_),
    .A2(_21050_),
    .ZN(_22526_)
  );
  AND2_X1 _30644_ (
    .A1(_21045_),
    .A2(_21053_),
    .ZN(_22527_)
  );
  INV_X1 _30645_ (
    .A(_22527_),
    .ZN(_22528_)
  );
  AND2_X1 _30646_ (
    .A1(_22526_),
    .A2(_22527_),
    .ZN(_22529_)
  );
  AND2_X1 _30647_ (
    .A1(_21198_),
    .A2(_21268_),
    .ZN(_22530_)
  );
  AND2_X1 _30648_ (
    .A1(_21042_),
    .A2(_21052_),
    .ZN(_22531_)
  );
  INV_X1 _30649_ (
    .A(_22531_),
    .ZN(_22532_)
  );
  AND2_X1 _30650_ (
    .A1(_22530_),
    .A2(_22531_),
    .ZN(_22533_)
  );
  AND2_X1 _30651_ (
    .A1(_22529_),
    .A2(_22533_),
    .ZN(_22534_)
  );
  AND2_X1 _30652_ (
    .A1(_22525_),
    .A2(_22534_),
    .ZN(_22535_)
  );
  AND2_X1 _30653_ (
    .A1(_22521_),
    .A2(_22535_),
    .ZN(_22536_)
  );
  AND2_X1 _30654_ (
    .A1(_22510_),
    .A2(_22536_),
    .ZN(_22537_)
  );
  INV_X1 _30655_ (
    .A(_22537_),
    .ZN(_22538_)
  );
  AND2_X1 _30656_ (
    .A1(_22070_),
    .A2(_22499_),
    .ZN(_22539_)
  );
  AND2_X1 _30657_ (
    .A1(_22538_),
    .A2(_22539_),
    .ZN(_22540_)
  );
  AND2_X1 _30658_ (
    .A1(_22019_),
    .A2(_22020_),
    .ZN(_22541_)
  );
  AND2_X1 _30659_ (
    .A1(_22021_),
    .A2(_22023_),
    .ZN(_22542_)
  );
  AND2_X1 _30660_ (
    .A1(_22541_),
    .A2(_22542_),
    .ZN(_22543_)
  );
  AND2_X1 _30661_ (
    .A1(_22022_),
    .A2(_22543_),
    .ZN(_22544_)
  );
  INV_X1 _30662_ (
    .A(_22544_),
    .ZN(_22545_)
  );
  AND2_X1 _30663_ (
    .A1(_22540_),
    .A2(_22545_),
    .ZN(_22546_)
  );
  AND2_X1 _30664_ (
    .A1(_22414_),
    .A2(_22546_),
    .ZN(_22547_)
  );
  AND2_X1 _30665_ (
    .A1(_22496_),
    .A2(_22547_),
    .ZN(_22548_)
  );
  INV_X1 _30666_ (
    .A(_22548_),
    .ZN(_22549_)
  );
  AND2_X1 _30667_ (
    .A1(_22337_),
    .A2(_22549_),
    .ZN(_22550_)
  );
  INV_X1 _30668_ (
    .A(_22550_),
    .ZN(_22551_)
  );
  AND2_X1 _30669_ (
    .A1(_22271_),
    .A2(_22551_),
    .ZN(_22552_)
  );
  INV_X1 _30670_ (
    .A(_22552_),
    .ZN(_22553_)
  );
  AND2_X1 _30671_ (
    .A1(_21038_),
    .A2(_22320_),
    .ZN(_22554_)
  );
  INV_X1 _30672_ (
    .A(_22554_),
    .ZN(_22555_)
  );
  AND2_X1 _30673_ (
    .A1(_21069_),
    .A2(_22323_),
    .ZN(_22556_)
  );
  INV_X1 _30674_ (
    .A(_22556_),
    .ZN(_22557_)
  );
  AND2_X1 _30675_ (
    .A1(_22555_),
    .A2(_22557_),
    .ZN(_22558_)
  );
  INV_X1 _30676_ (
    .A(_22558_),
    .ZN(_22559_)
  );
  AND2_X1 _30677_ (
    .A1(reg_op1[0]),
    .A2(decoded_imm[0]),
    .ZN(_22560_)
  );
  INV_X1 _30678_ (
    .A(_22560_),
    .ZN(_22561_)
  );
  AND2_X1 _30679_ (
    .A1(_21168_),
    .A2(_21286_),
    .ZN(_22562_)
  );
  INV_X1 _30680_ (
    .A(_22562_),
    .ZN(_22563_)
  );
  AND2_X1 _30681_ (
    .A1(_22561_),
    .A2(_22563_),
    .ZN(_22564_)
  );
  AND2_X1 _30682_ (
    .A1(_22559_),
    .A2(_22564_),
    .ZN(_22565_)
  );
  INV_X1 _30683_ (
    .A(_22565_),
    .ZN(_22566_)
  );
  AND2_X1 _30684_ (
    .A1(_22029_),
    .A2(_22217_),
    .ZN(_22567_)
  );
  INV_X1 _30685_ (
    .A(_22567_),
    .ZN(_22568_)
  );
  AND2_X1 _30686_ (
    .A1(_29149_[4]),
    .A2(_22277_),
    .ZN(_22569_)
  );
  AND2_X1 _30687_ (
    .A1(_22568_),
    .A2(_22569_),
    .ZN(_22570_)
  );
  INV_X1 _30688_ (
    .A(_22570_),
    .ZN(_22571_)
  );
  AND2_X1 _30689_ (
    .A1(_22028_),
    .A2(_22571_),
    .ZN(_22572_)
  );
  INV_X1 _30690_ (
    .A(_22572_),
    .ZN(_22573_)
  );
  AND2_X1 _30691_ (
    .A1(reg_op1[4]),
    .A2(_22290_),
    .ZN(_22574_)
  );
  INV_X1 _30692_ (
    .A(_22574_),
    .ZN(_22575_)
  );
  AND2_X1 _30693_ (
    .A1(reg_op1[1]),
    .A2(_22290_),
    .ZN(_22576_)
  );
  AND2_X1 _30694_ (
    .A1(_21168_),
    .A2(_22334_),
    .ZN(_22577_)
  );
  INV_X1 _30695_ (
    .A(_22577_),
    .ZN(_22578_)
  );
  AND2_X1 _30696_ (
    .A1(_22572_),
    .A2(_22576_),
    .ZN(_22579_)
  );
  INV_X1 _30697_ (
    .A(_22579_),
    .ZN(_22580_)
  );
  AND2_X1 _30698_ (
    .A1(_22573_),
    .A2(_22574_),
    .ZN(_22581_)
  );
  INV_X1 _30699_ (
    .A(_22581_),
    .ZN(_22582_)
  );
  AND2_X1 _30700_ (
    .A1(_22580_),
    .A2(_22582_),
    .ZN(_22583_)
  );
  INV_X1 _30701_ (
    .A(_22583_),
    .ZN(_22584_)
  );
  AND2_X1 _30702_ (
    .A1(_22295_),
    .A2(_22584_),
    .ZN(_22585_)
  );
  INV_X1 _30703_ (
    .A(_22585_),
    .ZN(_22586_)
  );
  AND2_X1 _30704_ (
    .A1(_22566_),
    .A2(_22586_),
    .ZN(_22587_)
  );
  AND2_X1 _30705_ (
    .A1(_22553_),
    .A2(_22587_),
    .ZN(_22588_)
  );
  AND2_X1 _30706_ (
    .A1(_22333_),
    .A2(_22588_),
    .ZN(_22589_)
  );
  INV_X1 _30707_ (
    .A(_22589_),
    .ZN(_22590_)
  );
  AND2_X1 _30708_ (
    .A1(_22578_),
    .A2(_22590_),
    .ZN(_00058_)
  );
  AND2_X1 _30709_ (
    .A1(reg_pc[2]),
    .A2(_22335_),
    .ZN(_22591_)
  );
  INV_X1 _30710_ (
    .A(_22591_),
    .ZN(_22592_)
  );
  AND2_X1 _30711_ (
    .A1(_21867_),
    .A2(_22149_),
    .ZN(_22593_)
  );
  INV_X1 _30712_ (
    .A(_22593_),
    .ZN(_22594_)
  );
  AND2_X1 _30713_ (
    .A1(_21851_),
    .A2(_00008_[2]),
    .ZN(_22595_)
  );
  INV_X1 _30714_ (
    .A(_22595_),
    .ZN(_22596_)
  );
  AND2_X1 _30715_ (
    .A1(_22594_),
    .A2(_22596_),
    .ZN(_22597_)
  );
  AND2_X1 _30716_ (
    .A1(_22147_),
    .A2(_22597_),
    .ZN(_22598_)
  );
  INV_X1 _30717_ (
    .A(_22598_),
    .ZN(_22599_)
  );
  AND2_X1 _30718_ (
    .A1(_21939_),
    .A2(_00008_[2]),
    .ZN(_22600_)
  );
  INV_X1 _30719_ (
    .A(_22600_),
    .ZN(_22601_)
  );
  AND2_X1 _30720_ (
    .A1(_21923_),
    .A2(_22149_),
    .ZN(_22602_)
  );
  INV_X1 _30721_ (
    .A(_22602_),
    .ZN(_22603_)
  );
  AND2_X1 _30722_ (
    .A1(_00008_[0]),
    .A2(_22603_),
    .ZN(_22604_)
  );
  AND2_X1 _30723_ (
    .A1(_22601_),
    .A2(_22604_),
    .ZN(_22605_)
  );
  INV_X1 _30724_ (
    .A(_22605_),
    .ZN(_22606_)
  );
  AND2_X1 _30725_ (
    .A1(_22599_),
    .A2(_22606_),
    .ZN(_22607_)
  );
  AND2_X1 _30726_ (
    .A1(_00008_[3]),
    .A2(_22607_),
    .ZN(_22608_)
  );
  INV_X1 _30727_ (
    .A(_22608_),
    .ZN(_22609_)
  );
  AND2_X1 _30728_ (
    .A1(\cpuregs[18] [2]),
    .A2(_22149_),
    .ZN(_22610_)
  );
  INV_X1 _30729_ (
    .A(_22610_),
    .ZN(_22611_)
  );
  AND2_X1 _30730_ (
    .A1(\cpuregs[22] [2]),
    .A2(_00008_[2]),
    .ZN(_22612_)
  );
  INV_X1 _30731_ (
    .A(_22612_),
    .ZN(_22613_)
  );
  AND2_X1 _30732_ (
    .A1(_22147_),
    .A2(_22613_),
    .ZN(_22614_)
  );
  AND2_X1 _30733_ (
    .A1(_22611_),
    .A2(_22614_),
    .ZN(_22615_)
  );
  INV_X1 _30734_ (
    .A(_22615_),
    .ZN(_22616_)
  );
  AND2_X1 _30735_ (
    .A1(\cpuregs[19] [2]),
    .A2(_22149_),
    .ZN(_22617_)
  );
  INV_X1 _30736_ (
    .A(_22617_),
    .ZN(_22618_)
  );
  AND2_X1 _30737_ (
    .A1(\cpuregs[23] [2]),
    .A2(_00008_[2]),
    .ZN(_22619_)
  );
  INV_X1 _30738_ (
    .A(_22619_),
    .ZN(_22620_)
  );
  AND2_X1 _30739_ (
    .A1(_00008_[0]),
    .A2(_22620_),
    .ZN(_22621_)
  );
  AND2_X1 _30740_ (
    .A1(_22618_),
    .A2(_22621_),
    .ZN(_22622_)
  );
  INV_X1 _30741_ (
    .A(_22622_),
    .ZN(_22623_)
  );
  AND2_X1 _30742_ (
    .A1(_22616_),
    .A2(_22623_),
    .ZN(_22624_)
  );
  INV_X1 _30743_ (
    .A(_22624_),
    .ZN(_22625_)
  );
  AND2_X1 _30744_ (
    .A1(_22150_),
    .A2(_22625_),
    .ZN(_22626_)
  );
  INV_X1 _30745_ (
    .A(_22626_),
    .ZN(_22627_)
  );
  AND2_X1 _30746_ (
    .A1(_22609_),
    .A2(_22627_),
    .ZN(_22628_)
  );
  AND2_X1 _30747_ (
    .A1(\cpuregs[17] [2]),
    .A2(_22149_),
    .ZN(_22629_)
  );
  INV_X1 _30748_ (
    .A(_22629_),
    .ZN(_22630_)
  );
  AND2_X1 _30749_ (
    .A1(\cpuregs[21] [2]),
    .A2(_00008_[2]),
    .ZN(_22631_)
  );
  INV_X1 _30750_ (
    .A(_22631_),
    .ZN(_22632_)
  );
  AND2_X1 _30751_ (
    .A1(_00008_[0]),
    .A2(_22632_),
    .ZN(_22633_)
  );
  AND2_X1 _30752_ (
    .A1(_22630_),
    .A2(_22633_),
    .ZN(_22634_)
  );
  INV_X1 _30753_ (
    .A(_22634_),
    .ZN(_22635_)
  );
  AND2_X1 _30754_ (
    .A1(\cpuregs[20] [2]),
    .A2(_00008_[2]),
    .ZN(_22636_)
  );
  INV_X1 _30755_ (
    .A(_22636_),
    .ZN(_22637_)
  );
  AND2_X1 _30756_ (
    .A1(\cpuregs[16] [2]),
    .A2(_22149_),
    .ZN(_22638_)
  );
  INV_X1 _30757_ (
    .A(_22638_),
    .ZN(_22639_)
  );
  AND2_X1 _30758_ (
    .A1(_22147_),
    .A2(_22639_),
    .ZN(_22640_)
  );
  AND2_X1 _30759_ (
    .A1(_22637_),
    .A2(_22640_),
    .ZN(_22641_)
  );
  INV_X1 _30760_ (
    .A(_22641_),
    .ZN(_22642_)
  );
  AND2_X1 _30761_ (
    .A1(_22635_),
    .A2(_22642_),
    .ZN(_22643_)
  );
  INV_X1 _30762_ (
    .A(_22643_),
    .ZN(_22644_)
  );
  AND2_X1 _30763_ (
    .A1(_22150_),
    .A2(_22644_),
    .ZN(_22645_)
  );
  INV_X1 _30764_ (
    .A(_22645_),
    .ZN(_22646_)
  );
  AND2_X1 _30765_ (
    .A1(_21835_),
    .A2(_22149_),
    .ZN(_22647_)
  );
  INV_X1 _30766_ (
    .A(_22647_),
    .ZN(_22648_)
  );
  AND2_X1 _30767_ (
    .A1(_21891_),
    .A2(_00008_[2]),
    .ZN(_22649_)
  );
  INV_X1 _30768_ (
    .A(_22649_),
    .ZN(_22650_)
  );
  AND2_X1 _30769_ (
    .A1(_21569_),
    .A2(_22149_),
    .ZN(_22651_)
  );
  INV_X1 _30770_ (
    .A(_22651_),
    .ZN(_22652_)
  );
  AND2_X1 _30771_ (
    .A1(_21907_),
    .A2(_00008_[2]),
    .ZN(_22653_)
  );
  INV_X1 _30772_ (
    .A(_22653_),
    .ZN(_22654_)
  );
  AND2_X1 _30773_ (
    .A1(_22652_),
    .A2(_22654_),
    .ZN(_22655_)
  );
  AND2_X1 _30774_ (
    .A1(_00008_[0]),
    .A2(_22648_),
    .ZN(_22656_)
  );
  AND2_X1 _30775_ (
    .A1(_22650_),
    .A2(_22656_),
    .ZN(_22657_)
  );
  INV_X1 _30776_ (
    .A(_22657_),
    .ZN(_22658_)
  );
  AND2_X1 _30777_ (
    .A1(_22147_),
    .A2(_22655_),
    .ZN(_22659_)
  );
  INV_X1 _30778_ (
    .A(_22659_),
    .ZN(_22660_)
  );
  AND2_X1 _30779_ (
    .A1(_22658_),
    .A2(_22660_),
    .ZN(_22661_)
  );
  AND2_X1 _30780_ (
    .A1(_00008_[3]),
    .A2(_22661_),
    .ZN(_22662_)
  );
  INV_X1 _30781_ (
    .A(_22662_),
    .ZN(_22663_)
  );
  AND2_X1 _30782_ (
    .A1(_22148_),
    .A2(_22663_),
    .ZN(_22664_)
  );
  AND2_X1 _30783_ (
    .A1(_22646_),
    .A2(_22664_),
    .ZN(_22665_)
  );
  INV_X1 _30784_ (
    .A(_22665_),
    .ZN(_22666_)
  );
  AND2_X1 _30785_ (
    .A1(_00008_[1]),
    .A2(_22628_),
    .ZN(_22667_)
  );
  INV_X1 _30786_ (
    .A(_22667_),
    .ZN(_22668_)
  );
  AND2_X1 _30787_ (
    .A1(_00008_[4]),
    .A2(_22668_),
    .ZN(_22669_)
  );
  AND2_X1 _30788_ (
    .A1(_22666_),
    .A2(_22669_),
    .ZN(_22670_)
  );
  INV_X1 _30789_ (
    .A(_22670_),
    .ZN(_22671_)
  );
  AND2_X1 _30790_ (
    .A1(_21781_),
    .A2(_00008_[2]),
    .ZN(_22672_)
  );
  INV_X1 _30791_ (
    .A(_22672_),
    .ZN(_22673_)
  );
  AND2_X1 _30792_ (
    .A1(_21489_),
    .A2(_22149_),
    .ZN(_22674_)
  );
  INV_X1 _30793_ (
    .A(_22674_),
    .ZN(_22675_)
  );
  AND2_X1 _30794_ (
    .A1(_21539_),
    .A2(_22149_),
    .ZN(_22676_)
  );
  INV_X1 _30795_ (
    .A(_22676_),
    .ZN(_22677_)
  );
  AND2_X1 _30796_ (
    .A1(_21806_),
    .A2(_00008_[2]),
    .ZN(_22678_)
  );
  INV_X1 _30797_ (
    .A(_22678_),
    .ZN(_22679_)
  );
  AND2_X1 _30798_ (
    .A1(_22677_),
    .A2(_22679_),
    .ZN(_22680_)
  );
  AND2_X1 _30799_ (
    .A1(_00008_[0]),
    .A2(_22675_),
    .ZN(_22681_)
  );
  AND2_X1 _30800_ (
    .A1(_22673_),
    .A2(_22681_),
    .ZN(_22682_)
  );
  INV_X1 _30801_ (
    .A(_22682_),
    .ZN(_22683_)
  );
  AND2_X1 _30802_ (
    .A1(_22147_),
    .A2(_22680_),
    .ZN(_22684_)
  );
  INV_X1 _30803_ (
    .A(_22684_),
    .ZN(_22685_)
  );
  AND2_X1 _30804_ (
    .A1(_22683_),
    .A2(_22685_),
    .ZN(_22686_)
  );
  AND2_X1 _30805_ (
    .A1(_00008_[1]),
    .A2(_22686_),
    .ZN(_22687_)
  );
  INV_X1 _30806_ (
    .A(_22687_),
    .ZN(_22688_)
  );
  AND2_X1 _30807_ (
    .A1(_21514_),
    .A2(_22149_),
    .ZN(_22689_)
  );
  INV_X1 _30808_ (
    .A(_22689_),
    .ZN(_22690_)
  );
  AND2_X1 _30809_ (
    .A1(_21734_),
    .A2(_00008_[2]),
    .ZN(_22691_)
  );
  INV_X1 _30810_ (
    .A(_22691_),
    .ZN(_22692_)
  );
  AND2_X1 _30811_ (
    .A1(_21955_),
    .A2(_22149_),
    .ZN(_22693_)
  );
  INV_X1 _30812_ (
    .A(_22693_),
    .ZN(_22694_)
  );
  AND2_X1 _30813_ (
    .A1(_21671_),
    .A2(_00008_[2]),
    .ZN(_22695_)
  );
  INV_X1 _30814_ (
    .A(_22695_),
    .ZN(_22696_)
  );
  AND2_X1 _30815_ (
    .A1(_22694_),
    .A2(_22696_),
    .ZN(_22697_)
  );
  AND2_X1 _30816_ (
    .A1(_00008_[0]),
    .A2(_22690_),
    .ZN(_22698_)
  );
  AND2_X1 _30817_ (
    .A1(_22692_),
    .A2(_22698_),
    .ZN(_22699_)
  );
  INV_X1 _30818_ (
    .A(_22699_),
    .ZN(_22700_)
  );
  AND2_X1 _30819_ (
    .A1(_22147_),
    .A2(_22697_),
    .ZN(_22701_)
  );
  INV_X1 _30820_ (
    .A(_22701_),
    .ZN(_22702_)
  );
  AND2_X1 _30821_ (
    .A1(_22700_),
    .A2(_22702_),
    .ZN(_22703_)
  );
  AND2_X1 _30822_ (
    .A1(_22148_),
    .A2(_22703_),
    .ZN(_22704_)
  );
  INV_X1 _30823_ (
    .A(_22704_),
    .ZN(_22705_)
  );
  AND2_X1 _30824_ (
    .A1(_22688_),
    .A2(_22705_),
    .ZN(_22706_)
  );
  INV_X1 _30825_ (
    .A(_22706_),
    .ZN(_22707_)
  );
  AND2_X1 _30826_ (
    .A1(_22150_),
    .A2(_22707_),
    .ZN(_22708_)
  );
  INV_X1 _30827_ (
    .A(_22708_),
    .ZN(_22709_)
  );
  AND2_X1 _30828_ (
    .A1(\cpuregs[9] [2]),
    .A2(_22148_),
    .ZN(_22710_)
  );
  INV_X1 _30829_ (
    .A(_22710_),
    .ZN(_22711_)
  );
  AND2_X1 _30830_ (
    .A1(\cpuregs[11] [2]),
    .A2(_00008_[1]),
    .ZN(_22712_)
  );
  INV_X1 _30831_ (
    .A(_22712_),
    .ZN(_22713_)
  );
  AND2_X1 _30832_ (
    .A1(_22149_),
    .A2(_22713_),
    .ZN(_22714_)
  );
  AND2_X1 _30833_ (
    .A1(_22711_),
    .A2(_22714_),
    .ZN(_22715_)
  );
  INV_X1 _30834_ (
    .A(_22715_),
    .ZN(_22716_)
  );
  AND2_X1 _30835_ (
    .A1(\cpuregs[13] [2]),
    .A2(_22148_),
    .ZN(_22717_)
  );
  INV_X1 _30836_ (
    .A(_22717_),
    .ZN(_22718_)
  );
  AND2_X1 _30837_ (
    .A1(\cpuregs[15] [2]),
    .A2(_00008_[1]),
    .ZN(_22719_)
  );
  INV_X1 _30838_ (
    .A(_22719_),
    .ZN(_22720_)
  );
  AND2_X1 _30839_ (
    .A1(_00008_[2]),
    .A2(_22720_),
    .ZN(_22721_)
  );
  AND2_X1 _30840_ (
    .A1(_22718_),
    .A2(_22721_),
    .ZN(_22722_)
  );
  INV_X1 _30841_ (
    .A(_22722_),
    .ZN(_22723_)
  );
  AND2_X1 _30842_ (
    .A1(_22716_),
    .A2(_22723_),
    .ZN(_22724_)
  );
  INV_X1 _30843_ (
    .A(_22724_),
    .ZN(_22725_)
  );
  AND2_X1 _30844_ (
    .A1(_00008_[0]),
    .A2(_22725_),
    .ZN(_22726_)
  );
  INV_X1 _30845_ (
    .A(_22726_),
    .ZN(_22727_)
  );
  AND2_X1 _30846_ (
    .A1(\cpuregs[8] [2]),
    .A2(_22148_),
    .ZN(_22728_)
  );
  INV_X1 _30847_ (
    .A(_22728_),
    .ZN(_22729_)
  );
  AND2_X1 _30848_ (
    .A1(\cpuregs[10] [2]),
    .A2(_00008_[1]),
    .ZN(_22730_)
  );
  INV_X1 _30849_ (
    .A(_22730_),
    .ZN(_22731_)
  );
  AND2_X1 _30850_ (
    .A1(_22149_),
    .A2(_22731_),
    .ZN(_22732_)
  );
  AND2_X1 _30851_ (
    .A1(_22729_),
    .A2(_22732_),
    .ZN(_22733_)
  );
  INV_X1 _30852_ (
    .A(_22733_),
    .ZN(_22734_)
  );
  AND2_X1 _30853_ (
    .A1(\cpuregs[12] [2]),
    .A2(_22148_),
    .ZN(_22735_)
  );
  INV_X1 _30854_ (
    .A(_22735_),
    .ZN(_22736_)
  );
  AND2_X1 _30855_ (
    .A1(\cpuregs[14] [2]),
    .A2(_00008_[1]),
    .ZN(_22737_)
  );
  INV_X1 _30856_ (
    .A(_22737_),
    .ZN(_22738_)
  );
  AND2_X1 _30857_ (
    .A1(_00008_[2]),
    .A2(_22738_),
    .ZN(_22739_)
  );
  AND2_X1 _30858_ (
    .A1(_22736_),
    .A2(_22739_),
    .ZN(_22740_)
  );
  INV_X1 _30859_ (
    .A(_22740_),
    .ZN(_22741_)
  );
  AND2_X1 _30860_ (
    .A1(_22734_),
    .A2(_22741_),
    .ZN(_22742_)
  );
  INV_X1 _30861_ (
    .A(_22742_),
    .ZN(_22743_)
  );
  AND2_X1 _30862_ (
    .A1(_22147_),
    .A2(_22743_),
    .ZN(_22744_)
  );
  INV_X1 _30863_ (
    .A(_22744_),
    .ZN(_22745_)
  );
  AND2_X1 _30864_ (
    .A1(_22727_),
    .A2(_22745_),
    .ZN(_22746_)
  );
  INV_X1 _30865_ (
    .A(_22746_),
    .ZN(_22747_)
  );
  AND2_X1 _30866_ (
    .A1(_00008_[3]),
    .A2(_22747_),
    .ZN(_22748_)
  );
  INV_X1 _30867_ (
    .A(_22748_),
    .ZN(_22749_)
  );
  AND2_X1 _30868_ (
    .A1(_22709_),
    .A2(_22749_),
    .ZN(_22750_)
  );
  INV_X1 _30869_ (
    .A(_22750_),
    .ZN(_22751_)
  );
  AND2_X1 _30870_ (
    .A1(_22151_),
    .A2(_22751_),
    .ZN(_22752_)
  );
  INV_X1 _30871_ (
    .A(_22752_),
    .ZN(_22753_)
  );
  AND2_X1 _30872_ (
    .A1(_22546_),
    .A2(_22671_),
    .ZN(_22754_)
  );
  AND2_X1 _30873_ (
    .A1(_22753_),
    .A2(_22754_),
    .ZN(_22755_)
  );
  INV_X1 _30874_ (
    .A(_22755_),
    .ZN(_22756_)
  );
  AND2_X1 _30875_ (
    .A1(_22592_),
    .A2(_22756_),
    .ZN(_22757_)
  );
  INV_X1 _30876_ (
    .A(_22757_),
    .ZN(_22758_)
  );
  AND2_X1 _30877_ (
    .A1(_22271_),
    .A2(_22758_),
    .ZN(_22759_)
  );
  INV_X1 _30878_ (
    .A(_22759_),
    .ZN(_22760_)
  );
  AND2_X1 _30879_ (
    .A1(decoded_imm[1]),
    .A2(reg_op1[1]),
    .ZN(_22761_)
  );
  INV_X1 _30880_ (
    .A(_22761_),
    .ZN(_22762_)
  );
  AND2_X1 _30881_ (
    .A1(_22008_),
    .A2(_22024_),
    .ZN(_22763_)
  );
  INV_X1 _30882_ (
    .A(_22763_),
    .ZN(_22764_)
  );
  AND2_X1 _30883_ (
    .A1(_22762_),
    .A2(_22764_),
    .ZN(_22765_)
  );
  INV_X1 _30884_ (
    .A(_22765_),
    .ZN(_22766_)
  );
  AND2_X1 _30885_ (
    .A1(_22560_),
    .A2(_22765_),
    .ZN(_22767_)
  );
  INV_X1 _30886_ (
    .A(_22767_),
    .ZN(_22768_)
  );
  AND2_X1 _30887_ (
    .A1(_22762_),
    .A2(_22768_),
    .ZN(_22769_)
  );
  INV_X1 _30888_ (
    .A(_22769_),
    .ZN(_22770_)
  );
  AND2_X1 _30889_ (
    .A1(reg_op1[2]),
    .A2(decoded_imm[2]),
    .ZN(_22771_)
  );
  INV_X1 _30890_ (
    .A(_22771_),
    .ZN(_22772_)
  );
  AND2_X1 _30891_ (
    .A1(_21169_),
    .A2(_22007_),
    .ZN(_22773_)
  );
  INV_X1 _30892_ (
    .A(_22773_),
    .ZN(_22774_)
  );
  AND2_X1 _30893_ (
    .A1(_22772_),
    .A2(_22774_),
    .ZN(_22775_)
  );
  INV_X1 _30894_ (
    .A(_22775_),
    .ZN(_22776_)
  );
  AND2_X1 _30895_ (
    .A1(_22769_),
    .A2(_22776_),
    .ZN(_22777_)
  );
  INV_X1 _30896_ (
    .A(_22777_),
    .ZN(_22778_)
  );
  AND2_X1 _30897_ (
    .A1(_22770_),
    .A2(_22775_),
    .ZN(_22779_)
  );
  INV_X1 _30898_ (
    .A(_22779_),
    .ZN(_22780_)
  );
  AND2_X1 _30899_ (
    .A1(reg_op1[6]),
    .A2(_22290_),
    .ZN(_22781_)
  );
  INV_X1 _30900_ (
    .A(_22781_),
    .ZN(_22782_)
  );
  AND2_X1 _30901_ (
    .A1(_22573_),
    .A2(_22782_),
    .ZN(_22783_)
  );
  INV_X1 _30902_ (
    .A(_22783_),
    .ZN(_22784_)
  );
  AND2_X1 _30903_ (
    .A1(reg_op1[1]),
    .A2(_22285_),
    .ZN(_22785_)
  );
  INV_X1 _30904_ (
    .A(_22785_),
    .ZN(_22786_)
  );
  AND2_X1 _30905_ (
    .A1(reg_op1[3]),
    .A2(_22290_),
    .ZN(_22787_)
  );
  INV_X1 _30906_ (
    .A(_22787_),
    .ZN(_22788_)
  );
  AND2_X1 _30907_ (
    .A1(_22786_),
    .A2(_22788_),
    .ZN(_22789_)
  );
  AND2_X1 _30908_ (
    .A1(_22572_),
    .A2(_22789_),
    .ZN(_22790_)
  );
  INV_X1 _30909_ (
    .A(_22790_),
    .ZN(_22791_)
  );
  AND2_X1 _30910_ (
    .A1(_21169_),
    .A2(_22334_),
    .ZN(_22792_)
  );
  INV_X1 _30911_ (
    .A(_22792_),
    .ZN(_22793_)
  );
  AND2_X1 _30912_ (
    .A1(_22295_),
    .A2(_22784_),
    .ZN(_22794_)
  );
  AND2_X1 _30913_ (
    .A1(_22791_),
    .A2(_22794_),
    .ZN(_22795_)
  );
  INV_X1 _30914_ (
    .A(_22795_),
    .ZN(_22796_)
  );
  AND2_X1 _30915_ (
    .A1(_22559_),
    .A2(_22780_),
    .ZN(_22797_)
  );
  AND2_X1 _30916_ (
    .A1(_22778_),
    .A2(_22797_),
    .ZN(_22798_)
  );
  INV_X1 _30917_ (
    .A(_22798_),
    .ZN(_22799_)
  );
  AND2_X1 _30918_ (
    .A1(_22796_),
    .A2(_22799_),
    .ZN(_22800_)
  );
  AND2_X1 _30919_ (
    .A1(_22333_),
    .A2(_22800_),
    .ZN(_22801_)
  );
  AND2_X1 _30920_ (
    .A1(_22760_),
    .A2(_22801_),
    .ZN(_22802_)
  );
  INV_X1 _30921_ (
    .A(_22802_),
    .ZN(_22803_)
  );
  AND2_X1 _30922_ (
    .A1(_22793_),
    .A2(_22803_),
    .ZN(_00059_)
  );
  AND2_X1 _30923_ (
    .A1(reg_pc[3]),
    .A2(_22335_),
    .ZN(_22804_)
  );
  INV_X1 _30924_ (
    .A(_22804_),
    .ZN(_22805_)
  );
  AND2_X1 _30925_ (
    .A1(\cpuregs[26] [3]),
    .A2(_22149_),
    .ZN(_22806_)
  );
  INV_X1 _30926_ (
    .A(_22806_),
    .ZN(_22807_)
  );
  AND2_X1 _30927_ (
    .A1(\cpuregs[30] [3]),
    .A2(_00008_[2]),
    .ZN(_22808_)
  );
  INV_X1 _30928_ (
    .A(_22808_),
    .ZN(_22809_)
  );
  AND2_X1 _30929_ (
    .A1(_22147_),
    .A2(_22809_),
    .ZN(_22810_)
  );
  AND2_X1 _30930_ (
    .A1(_22807_),
    .A2(_22810_),
    .ZN(_22811_)
  );
  INV_X1 _30931_ (
    .A(_22811_),
    .ZN(_22812_)
  );
  AND2_X1 _30932_ (
    .A1(\cpuregs[31] [3]),
    .A2(_00008_[2]),
    .ZN(_22813_)
  );
  INV_X1 _30933_ (
    .A(_22813_),
    .ZN(_22814_)
  );
  AND2_X1 _30934_ (
    .A1(\cpuregs[27] [3]),
    .A2(_22149_),
    .ZN(_22815_)
  );
  INV_X1 _30935_ (
    .A(_22815_),
    .ZN(_22816_)
  );
  AND2_X1 _30936_ (
    .A1(_00008_[0]),
    .A2(_22816_),
    .ZN(_22817_)
  );
  AND2_X1 _30937_ (
    .A1(_22814_),
    .A2(_22817_),
    .ZN(_22818_)
  );
  INV_X1 _30938_ (
    .A(_22818_),
    .ZN(_22819_)
  );
  AND2_X1 _30939_ (
    .A1(_22812_),
    .A2(_22819_),
    .ZN(_22820_)
  );
  INV_X1 _30940_ (
    .A(_22820_),
    .ZN(_22821_)
  );
  AND2_X1 _30941_ (
    .A1(_00008_[1]),
    .A2(_22821_),
    .ZN(_22822_)
  );
  INV_X1 _30942_ (
    .A(_22822_),
    .ZN(_22823_)
  );
  AND2_X1 _30943_ (
    .A1(\cpuregs[24] [3]),
    .A2(_22149_),
    .ZN(_22824_)
  );
  INV_X1 _30944_ (
    .A(_22824_),
    .ZN(_22825_)
  );
  AND2_X1 _30945_ (
    .A1(\cpuregs[28] [3]),
    .A2(_00008_[2]),
    .ZN(_22826_)
  );
  INV_X1 _30946_ (
    .A(_22826_),
    .ZN(_22827_)
  );
  AND2_X1 _30947_ (
    .A1(_22147_),
    .A2(_22827_),
    .ZN(_22828_)
  );
  AND2_X1 _30948_ (
    .A1(_22825_),
    .A2(_22828_),
    .ZN(_22829_)
  );
  INV_X1 _30949_ (
    .A(_22829_),
    .ZN(_22830_)
  );
  AND2_X1 _30950_ (
    .A1(\cpuregs[25] [3]),
    .A2(_22149_),
    .ZN(_22831_)
  );
  INV_X1 _30951_ (
    .A(_22831_),
    .ZN(_22832_)
  );
  AND2_X1 _30952_ (
    .A1(\cpuregs[29] [3]),
    .A2(_00008_[2]),
    .ZN(_22833_)
  );
  INV_X1 _30953_ (
    .A(_22833_),
    .ZN(_22834_)
  );
  AND2_X1 _30954_ (
    .A1(_00008_[0]),
    .A2(_22834_),
    .ZN(_22835_)
  );
  AND2_X1 _30955_ (
    .A1(_22832_),
    .A2(_22835_),
    .ZN(_22836_)
  );
  INV_X1 _30956_ (
    .A(_22836_),
    .ZN(_22837_)
  );
  AND2_X1 _30957_ (
    .A1(_22830_),
    .A2(_22837_),
    .ZN(_22838_)
  );
  INV_X1 _30958_ (
    .A(_22838_),
    .ZN(_22839_)
  );
  AND2_X1 _30959_ (
    .A1(_22148_),
    .A2(_22839_),
    .ZN(_22840_)
  );
  INV_X1 _30960_ (
    .A(_22840_),
    .ZN(_22841_)
  );
  AND2_X1 _30961_ (
    .A1(_21373_),
    .A2(_00008_[2]),
    .ZN(_22842_)
  );
  INV_X1 _30962_ (
    .A(_22842_),
    .ZN(_22843_)
  );
  AND2_X1 _30963_ (
    .A1(_21619_),
    .A2(_22149_),
    .ZN(_22844_)
  );
  INV_X1 _30964_ (
    .A(_22844_),
    .ZN(_22845_)
  );
  AND2_X1 _30965_ (
    .A1(_21593_),
    .A2(_22149_),
    .ZN(_22846_)
  );
  INV_X1 _30966_ (
    .A(_22846_),
    .ZN(_22847_)
  );
  AND2_X1 _30967_ (
    .A1(_21411_),
    .A2(_00008_[2]),
    .ZN(_22848_)
  );
  INV_X1 _30968_ (
    .A(_22848_),
    .ZN(_22849_)
  );
  AND2_X1 _30969_ (
    .A1(_22847_),
    .A2(_22849_),
    .ZN(_22850_)
  );
  AND2_X1 _30970_ (
    .A1(_00008_[0]),
    .A2(_22845_),
    .ZN(_22851_)
  );
  AND2_X1 _30971_ (
    .A1(_22843_),
    .A2(_22851_),
    .ZN(_22852_)
  );
  INV_X1 _30972_ (
    .A(_22852_),
    .ZN(_22853_)
  );
  AND2_X1 _30973_ (
    .A1(_22147_),
    .A2(_22850_),
    .ZN(_22854_)
  );
  INV_X1 _30974_ (
    .A(_22854_),
    .ZN(_22855_)
  );
  AND2_X1 _30975_ (
    .A1(_22853_),
    .A2(_22855_),
    .ZN(_22856_)
  );
  AND2_X1 _30976_ (
    .A1(_00008_[1]),
    .A2(_22856_),
    .ZN(_22857_)
  );
  INV_X1 _30977_ (
    .A(_22857_),
    .ZN(_22858_)
  );
  AND2_X1 _30978_ (
    .A1(_21461_),
    .A2(_22149_),
    .ZN(_22859_)
  );
  INV_X1 _30979_ (
    .A(_22859_),
    .ZN(_22860_)
  );
  AND2_X1 _30980_ (
    .A1(_21760_),
    .A2(_00008_[2]),
    .ZN(_22861_)
  );
  INV_X1 _30981_ (
    .A(_22861_),
    .ZN(_22862_)
  );
  AND2_X1 _30982_ (
    .A1(_21439_),
    .A2(_22149_),
    .ZN(_22863_)
  );
  INV_X1 _30983_ (
    .A(_22863_),
    .ZN(_22864_)
  );
  AND2_X1 _30984_ (
    .A1(_21650_),
    .A2(_00008_[2]),
    .ZN(_22865_)
  );
  INV_X1 _30985_ (
    .A(_22865_),
    .ZN(_22866_)
  );
  AND2_X1 _30986_ (
    .A1(_22864_),
    .A2(_22866_),
    .ZN(_22867_)
  );
  AND2_X1 _30987_ (
    .A1(_00008_[0]),
    .A2(_22860_),
    .ZN(_22868_)
  );
  AND2_X1 _30988_ (
    .A1(_22862_),
    .A2(_22868_),
    .ZN(_22869_)
  );
  INV_X1 _30989_ (
    .A(_22869_),
    .ZN(_22870_)
  );
  AND2_X1 _30990_ (
    .A1(_22147_),
    .A2(_22867_),
    .ZN(_22871_)
  );
  INV_X1 _30991_ (
    .A(_22871_),
    .ZN(_22872_)
  );
  AND2_X1 _30992_ (
    .A1(_22870_),
    .A2(_22872_),
    .ZN(_22873_)
  );
  AND2_X1 _30993_ (
    .A1(_22148_),
    .A2(_22873_),
    .ZN(_22874_)
  );
  INV_X1 _30994_ (
    .A(_22874_),
    .ZN(_22875_)
  );
  AND2_X1 _30995_ (
    .A1(_22858_),
    .A2(_22875_),
    .ZN(_22876_)
  );
  AND2_X1 _30996_ (
    .A1(_22150_),
    .A2(_22876_),
    .ZN(_22877_)
  );
  INV_X1 _30997_ (
    .A(_22877_),
    .ZN(_22878_)
  );
  AND2_X1 _30998_ (
    .A1(_00008_[3]),
    .A2(_22841_),
    .ZN(_22879_)
  );
  AND2_X1 _30999_ (
    .A1(_22823_),
    .A2(_22879_),
    .ZN(_22880_)
  );
  INV_X1 _31000_ (
    .A(_22880_),
    .ZN(_22881_)
  );
  AND2_X1 _31001_ (
    .A1(_00008_[4]),
    .A2(_22881_),
    .ZN(_22882_)
  );
  AND2_X1 _31002_ (
    .A1(_22878_),
    .A2(_22882_),
    .ZN(_22883_)
  );
  INV_X1 _31003_ (
    .A(_22883_),
    .ZN(_22884_)
  );
  AND2_X1 _31004_ (
    .A1(_21782_),
    .A2(_00008_[2]),
    .ZN(_22885_)
  );
  INV_X1 _31005_ (
    .A(_22885_),
    .ZN(_22886_)
  );
  AND2_X1 _31006_ (
    .A1(_21490_),
    .A2(_22149_),
    .ZN(_22887_)
  );
  INV_X1 _31007_ (
    .A(_22887_),
    .ZN(_22888_)
  );
  AND2_X1 _31008_ (
    .A1(_21540_),
    .A2(_22149_),
    .ZN(_22889_)
  );
  INV_X1 _31009_ (
    .A(_22889_),
    .ZN(_22890_)
  );
  AND2_X1 _31010_ (
    .A1(_21807_),
    .A2(_00008_[2]),
    .ZN(_22891_)
  );
  INV_X1 _31011_ (
    .A(_22891_),
    .ZN(_22892_)
  );
  AND2_X1 _31012_ (
    .A1(_22890_),
    .A2(_22892_),
    .ZN(_22893_)
  );
  AND2_X1 _31013_ (
    .A1(_00008_[0]),
    .A2(_22888_),
    .ZN(_22894_)
  );
  AND2_X1 _31014_ (
    .A1(_22886_),
    .A2(_22894_),
    .ZN(_22895_)
  );
  INV_X1 _31015_ (
    .A(_22895_),
    .ZN(_22896_)
  );
  AND2_X1 _31016_ (
    .A1(_22147_),
    .A2(_22893_),
    .ZN(_22897_)
  );
  INV_X1 _31017_ (
    .A(_22897_),
    .ZN(_22898_)
  );
  AND2_X1 _31018_ (
    .A1(_22896_),
    .A2(_22898_),
    .ZN(_22899_)
  );
  AND2_X1 _31019_ (
    .A1(_00008_[1]),
    .A2(_22899_),
    .ZN(_22900_)
  );
  INV_X1 _31020_ (
    .A(_22900_),
    .ZN(_22901_)
  );
  AND2_X1 _31021_ (
    .A1(_21515_),
    .A2(_22149_),
    .ZN(_22902_)
  );
  INV_X1 _31022_ (
    .A(_22902_),
    .ZN(_22903_)
  );
  AND2_X1 _31023_ (
    .A1(_21735_),
    .A2(_00008_[2]),
    .ZN(_22904_)
  );
  INV_X1 _31024_ (
    .A(_22904_),
    .ZN(_22905_)
  );
  AND2_X1 _31025_ (
    .A1(_21956_),
    .A2(_22149_),
    .ZN(_22906_)
  );
  INV_X1 _31026_ (
    .A(_22906_),
    .ZN(_22907_)
  );
  AND2_X1 _31027_ (
    .A1(_21672_),
    .A2(_00008_[2]),
    .ZN(_22908_)
  );
  INV_X1 _31028_ (
    .A(_22908_),
    .ZN(_22909_)
  );
  AND2_X1 _31029_ (
    .A1(_22907_),
    .A2(_22909_),
    .ZN(_22910_)
  );
  AND2_X1 _31030_ (
    .A1(_00008_[0]),
    .A2(_22903_),
    .ZN(_22911_)
  );
  AND2_X1 _31031_ (
    .A1(_22905_),
    .A2(_22911_),
    .ZN(_22912_)
  );
  INV_X1 _31032_ (
    .A(_22912_),
    .ZN(_22913_)
  );
  AND2_X1 _31033_ (
    .A1(_22147_),
    .A2(_22910_),
    .ZN(_22914_)
  );
  INV_X1 _31034_ (
    .A(_22914_),
    .ZN(_22915_)
  );
  AND2_X1 _31035_ (
    .A1(_22913_),
    .A2(_22915_),
    .ZN(_22916_)
  );
  AND2_X1 _31036_ (
    .A1(_22148_),
    .A2(_22916_),
    .ZN(_22917_)
  );
  INV_X1 _31037_ (
    .A(_22917_),
    .ZN(_22918_)
  );
  AND2_X1 _31038_ (
    .A1(_22901_),
    .A2(_22918_),
    .ZN(_22919_)
  );
  INV_X1 _31039_ (
    .A(_22919_),
    .ZN(_22920_)
  );
  AND2_X1 _31040_ (
    .A1(_22150_),
    .A2(_22920_),
    .ZN(_22921_)
  );
  INV_X1 _31041_ (
    .A(_22921_),
    .ZN(_22922_)
  );
  AND2_X1 _31042_ (
    .A1(\cpuregs[9] [3]),
    .A2(_22148_),
    .ZN(_22923_)
  );
  INV_X1 _31043_ (
    .A(_22923_),
    .ZN(_22924_)
  );
  AND2_X1 _31044_ (
    .A1(\cpuregs[11] [3]),
    .A2(_00008_[1]),
    .ZN(_22925_)
  );
  INV_X1 _31045_ (
    .A(_22925_),
    .ZN(_22926_)
  );
  AND2_X1 _31046_ (
    .A1(_22149_),
    .A2(_22926_),
    .ZN(_22927_)
  );
  AND2_X1 _31047_ (
    .A1(_22924_),
    .A2(_22927_),
    .ZN(_22928_)
  );
  INV_X1 _31048_ (
    .A(_22928_),
    .ZN(_22929_)
  );
  AND2_X1 _31049_ (
    .A1(\cpuregs[13] [3]),
    .A2(_22148_),
    .ZN(_22930_)
  );
  INV_X1 _31050_ (
    .A(_22930_),
    .ZN(_22931_)
  );
  AND2_X1 _31051_ (
    .A1(\cpuregs[15] [3]),
    .A2(_00008_[1]),
    .ZN(_22932_)
  );
  INV_X1 _31052_ (
    .A(_22932_),
    .ZN(_22933_)
  );
  AND2_X1 _31053_ (
    .A1(_00008_[2]),
    .A2(_22933_),
    .ZN(_22934_)
  );
  AND2_X1 _31054_ (
    .A1(_22931_),
    .A2(_22934_),
    .ZN(_22935_)
  );
  INV_X1 _31055_ (
    .A(_22935_),
    .ZN(_22936_)
  );
  AND2_X1 _31056_ (
    .A1(_22929_),
    .A2(_22936_),
    .ZN(_22937_)
  );
  INV_X1 _31057_ (
    .A(_22937_),
    .ZN(_22938_)
  );
  AND2_X1 _31058_ (
    .A1(_00008_[0]),
    .A2(_22938_),
    .ZN(_22939_)
  );
  INV_X1 _31059_ (
    .A(_22939_),
    .ZN(_22940_)
  );
  AND2_X1 _31060_ (
    .A1(\cpuregs[8] [3]),
    .A2(_22148_),
    .ZN(_22941_)
  );
  INV_X1 _31061_ (
    .A(_22941_),
    .ZN(_22942_)
  );
  AND2_X1 _31062_ (
    .A1(\cpuregs[10] [3]),
    .A2(_00008_[1]),
    .ZN(_22943_)
  );
  INV_X1 _31063_ (
    .A(_22943_),
    .ZN(_22944_)
  );
  AND2_X1 _31064_ (
    .A1(_22149_),
    .A2(_22944_),
    .ZN(_22945_)
  );
  AND2_X1 _31065_ (
    .A1(_22942_),
    .A2(_22945_),
    .ZN(_22946_)
  );
  INV_X1 _31066_ (
    .A(_22946_),
    .ZN(_22947_)
  );
  AND2_X1 _31067_ (
    .A1(\cpuregs[12] [3]),
    .A2(_22148_),
    .ZN(_22948_)
  );
  INV_X1 _31068_ (
    .A(_22948_),
    .ZN(_22949_)
  );
  AND2_X1 _31069_ (
    .A1(\cpuregs[14] [3]),
    .A2(_00008_[1]),
    .ZN(_22950_)
  );
  INV_X1 _31070_ (
    .A(_22950_),
    .ZN(_22951_)
  );
  AND2_X1 _31071_ (
    .A1(_00008_[2]),
    .A2(_22951_),
    .ZN(_22952_)
  );
  AND2_X1 _31072_ (
    .A1(_22949_),
    .A2(_22952_),
    .ZN(_22953_)
  );
  INV_X1 _31073_ (
    .A(_22953_),
    .ZN(_22954_)
  );
  AND2_X1 _31074_ (
    .A1(_22947_),
    .A2(_22954_),
    .ZN(_22955_)
  );
  INV_X1 _31075_ (
    .A(_22955_),
    .ZN(_22956_)
  );
  AND2_X1 _31076_ (
    .A1(_22147_),
    .A2(_22956_),
    .ZN(_22957_)
  );
  INV_X1 _31077_ (
    .A(_22957_),
    .ZN(_22958_)
  );
  AND2_X1 _31078_ (
    .A1(_22940_),
    .A2(_22958_),
    .ZN(_22959_)
  );
  INV_X1 _31079_ (
    .A(_22959_),
    .ZN(_22960_)
  );
  AND2_X1 _31080_ (
    .A1(_00008_[3]),
    .A2(_22960_),
    .ZN(_22961_)
  );
  INV_X1 _31081_ (
    .A(_22961_),
    .ZN(_22962_)
  );
  AND2_X1 _31082_ (
    .A1(_22922_),
    .A2(_22962_),
    .ZN(_22963_)
  );
  INV_X1 _31083_ (
    .A(_22963_),
    .ZN(_22964_)
  );
  AND2_X1 _31084_ (
    .A1(_22151_),
    .A2(_22964_),
    .ZN(_22965_)
  );
  INV_X1 _31085_ (
    .A(_22965_),
    .ZN(_22966_)
  );
  AND2_X1 _31086_ (
    .A1(_22546_),
    .A2(_22884_),
    .ZN(_22967_)
  );
  AND2_X1 _31087_ (
    .A1(_22966_),
    .A2(_22967_),
    .ZN(_22968_)
  );
  INV_X1 _31088_ (
    .A(_22968_),
    .ZN(_22969_)
  );
  AND2_X1 _31089_ (
    .A1(_22805_),
    .A2(_22969_),
    .ZN(_22970_)
  );
  INV_X1 _31090_ (
    .A(_22970_),
    .ZN(_22971_)
  );
  AND2_X1 _31091_ (
    .A1(_22271_),
    .A2(_22971_),
    .ZN(_22972_)
  );
  INV_X1 _31092_ (
    .A(_22972_),
    .ZN(_22973_)
  );
  AND2_X1 _31093_ (
    .A1(reg_op1[2]),
    .A2(_22285_),
    .ZN(_22974_)
  );
  INV_X1 _31094_ (
    .A(_22974_),
    .ZN(_22975_)
  );
  AND2_X1 _31095_ (
    .A1(_22575_),
    .A2(_22975_),
    .ZN(_22976_)
  );
  AND2_X1 _31096_ (
    .A1(_22572_),
    .A2(_22976_),
    .ZN(_22977_)
  );
  INV_X1 _31097_ (
    .A(_22977_),
    .ZN(_22978_)
  );
  AND2_X1 _31098_ (
    .A1(reg_op1[7]),
    .A2(_22290_),
    .ZN(_22979_)
  );
  INV_X1 _31099_ (
    .A(_22979_),
    .ZN(_22980_)
  );
  AND2_X1 _31100_ (
    .A1(_22573_),
    .A2(_22980_),
    .ZN(_22981_)
  );
  INV_X1 _31101_ (
    .A(_22981_),
    .ZN(_22982_)
  );
  AND2_X1 _31102_ (
    .A1(_22295_),
    .A2(_22982_),
    .ZN(_22983_)
  );
  AND2_X1 _31103_ (
    .A1(_22978_),
    .A2(_22983_),
    .ZN(_22984_)
  );
  INV_X1 _31104_ (
    .A(_22984_),
    .ZN(_22985_)
  );
  AND2_X1 _31105_ (
    .A1(_22772_),
    .A2(_22780_),
    .ZN(_22986_)
  );
  INV_X1 _31106_ (
    .A(_22986_),
    .ZN(_22987_)
  );
  AND2_X1 _31107_ (
    .A1(reg_op1[3]),
    .A2(decoded_imm[3]),
    .ZN(_22988_)
  );
  INV_X1 _31108_ (
    .A(_22988_),
    .ZN(_22989_)
  );
  AND2_X1 _31109_ (
    .A1(_21170_),
    .A2(_22006_),
    .ZN(_22990_)
  );
  INV_X1 _31110_ (
    .A(_22990_),
    .ZN(_22991_)
  );
  AND2_X1 _31111_ (
    .A1(_22989_),
    .A2(_22991_),
    .ZN(_22992_)
  );
  INV_X1 _31112_ (
    .A(_22992_),
    .ZN(_22993_)
  );
  AND2_X1 _31113_ (
    .A1(_22986_),
    .A2(_22993_),
    .ZN(_22994_)
  );
  INV_X1 _31114_ (
    .A(_22994_),
    .ZN(_22995_)
  );
  AND2_X1 _31115_ (
    .A1(_22987_),
    .A2(_22992_),
    .ZN(_22996_)
  );
  INV_X1 _31116_ (
    .A(_22996_),
    .ZN(_22997_)
  );
  AND2_X1 _31117_ (
    .A1(_21170_),
    .A2(_22334_),
    .ZN(_22998_)
  );
  INV_X1 _31118_ (
    .A(_22998_),
    .ZN(_22999_)
  );
  AND2_X1 _31119_ (
    .A1(_22559_),
    .A2(_22997_),
    .ZN(_23000_)
  );
  AND2_X1 _31120_ (
    .A1(_22995_),
    .A2(_23000_),
    .ZN(_23001_)
  );
  INV_X1 _31121_ (
    .A(_23001_),
    .ZN(_23002_)
  );
  AND2_X1 _31122_ (
    .A1(_22985_),
    .A2(_23002_),
    .ZN(_23003_)
  );
  AND2_X1 _31123_ (
    .A1(_22333_),
    .A2(_23003_),
    .ZN(_23004_)
  );
  AND2_X1 _31124_ (
    .A1(_22973_),
    .A2(_23004_),
    .ZN(_23005_)
  );
  INV_X1 _31125_ (
    .A(_23005_),
    .ZN(_23006_)
  );
  AND2_X1 _31126_ (
    .A1(_22999_),
    .A2(_23006_),
    .ZN(_00060_)
  );
  AND2_X1 _31127_ (
    .A1(_21171_),
    .A2(_22334_),
    .ZN(_23007_)
  );
  INV_X1 _31128_ (
    .A(_23007_),
    .ZN(_23008_)
  );
  AND2_X1 _31129_ (
    .A1(reg_pc[4]),
    .A2(_22335_),
    .ZN(_23009_)
  );
  INV_X1 _31130_ (
    .A(_23009_),
    .ZN(_23010_)
  );
  AND2_X1 _31131_ (
    .A1(\cpuregs[26] [4]),
    .A2(_22149_),
    .ZN(_23011_)
  );
  INV_X1 _31132_ (
    .A(_23011_),
    .ZN(_23012_)
  );
  AND2_X1 _31133_ (
    .A1(\cpuregs[30] [4]),
    .A2(_00008_[2]),
    .ZN(_23013_)
  );
  INV_X1 _31134_ (
    .A(_23013_),
    .ZN(_23014_)
  );
  AND2_X1 _31135_ (
    .A1(_22147_),
    .A2(_23014_),
    .ZN(_23015_)
  );
  AND2_X1 _31136_ (
    .A1(_23012_),
    .A2(_23015_),
    .ZN(_23016_)
  );
  INV_X1 _31137_ (
    .A(_23016_),
    .ZN(_23017_)
  );
  AND2_X1 _31138_ (
    .A1(\cpuregs[31] [4]),
    .A2(_00008_[2]),
    .ZN(_23018_)
  );
  INV_X1 _31139_ (
    .A(_23018_),
    .ZN(_23019_)
  );
  AND2_X1 _31140_ (
    .A1(\cpuregs[27] [4]),
    .A2(_22149_),
    .ZN(_23020_)
  );
  INV_X1 _31141_ (
    .A(_23020_),
    .ZN(_23021_)
  );
  AND2_X1 _31142_ (
    .A1(_00008_[0]),
    .A2(_23021_),
    .ZN(_23022_)
  );
  AND2_X1 _31143_ (
    .A1(_23019_),
    .A2(_23022_),
    .ZN(_23023_)
  );
  INV_X1 _31144_ (
    .A(_23023_),
    .ZN(_23024_)
  );
  AND2_X1 _31145_ (
    .A1(_23017_),
    .A2(_23024_),
    .ZN(_23025_)
  );
  INV_X1 _31146_ (
    .A(_23025_),
    .ZN(_23026_)
  );
  AND2_X1 _31147_ (
    .A1(_00008_[1]),
    .A2(_23026_),
    .ZN(_23027_)
  );
  INV_X1 _31148_ (
    .A(_23027_),
    .ZN(_23028_)
  );
  AND2_X1 _31149_ (
    .A1(\cpuregs[24] [4]),
    .A2(_22149_),
    .ZN(_23029_)
  );
  INV_X1 _31150_ (
    .A(_23029_),
    .ZN(_23030_)
  );
  AND2_X1 _31151_ (
    .A1(\cpuregs[28] [4]),
    .A2(_00008_[2]),
    .ZN(_23031_)
  );
  INV_X1 _31152_ (
    .A(_23031_),
    .ZN(_23032_)
  );
  AND2_X1 _31153_ (
    .A1(_22147_),
    .A2(_23032_),
    .ZN(_23033_)
  );
  AND2_X1 _31154_ (
    .A1(_23030_),
    .A2(_23033_),
    .ZN(_23034_)
  );
  INV_X1 _31155_ (
    .A(_23034_),
    .ZN(_23035_)
  );
  AND2_X1 _31156_ (
    .A1(\cpuregs[25] [4]),
    .A2(_22149_),
    .ZN(_23036_)
  );
  INV_X1 _31157_ (
    .A(_23036_),
    .ZN(_23037_)
  );
  AND2_X1 _31158_ (
    .A1(\cpuregs[29] [4]),
    .A2(_00008_[2]),
    .ZN(_23038_)
  );
  INV_X1 _31159_ (
    .A(_23038_),
    .ZN(_23039_)
  );
  AND2_X1 _31160_ (
    .A1(_00008_[0]),
    .A2(_23039_),
    .ZN(_23040_)
  );
  AND2_X1 _31161_ (
    .A1(_23037_),
    .A2(_23040_),
    .ZN(_23041_)
  );
  INV_X1 _31162_ (
    .A(_23041_),
    .ZN(_23042_)
  );
  AND2_X1 _31163_ (
    .A1(_23035_),
    .A2(_23042_),
    .ZN(_23043_)
  );
  INV_X1 _31164_ (
    .A(_23043_),
    .ZN(_23044_)
  );
  AND2_X1 _31165_ (
    .A1(_22148_),
    .A2(_23044_),
    .ZN(_23045_)
  );
  INV_X1 _31166_ (
    .A(_23045_),
    .ZN(_23046_)
  );
  AND2_X1 _31167_ (
    .A1(_21374_),
    .A2(_00008_[2]),
    .ZN(_23047_)
  );
  INV_X1 _31168_ (
    .A(_23047_),
    .ZN(_23048_)
  );
  AND2_X1 _31169_ (
    .A1(_21620_),
    .A2(_22149_),
    .ZN(_23049_)
  );
  INV_X1 _31170_ (
    .A(_23049_),
    .ZN(_23050_)
  );
  AND2_X1 _31171_ (
    .A1(_21594_),
    .A2(_22149_),
    .ZN(_23051_)
  );
  INV_X1 _31172_ (
    .A(_23051_),
    .ZN(_23052_)
  );
  AND2_X1 _31173_ (
    .A1(_21412_),
    .A2(_00008_[2]),
    .ZN(_23053_)
  );
  INV_X1 _31174_ (
    .A(_23053_),
    .ZN(_23054_)
  );
  AND2_X1 _31175_ (
    .A1(_23052_),
    .A2(_23054_),
    .ZN(_23055_)
  );
  AND2_X1 _31176_ (
    .A1(_00008_[0]),
    .A2(_23050_),
    .ZN(_23056_)
  );
  AND2_X1 _31177_ (
    .A1(_23048_),
    .A2(_23056_),
    .ZN(_23057_)
  );
  INV_X1 _31178_ (
    .A(_23057_),
    .ZN(_23058_)
  );
  AND2_X1 _31179_ (
    .A1(_22147_),
    .A2(_23055_),
    .ZN(_23059_)
  );
  INV_X1 _31180_ (
    .A(_23059_),
    .ZN(_23060_)
  );
  AND2_X1 _31181_ (
    .A1(_23058_),
    .A2(_23060_),
    .ZN(_23061_)
  );
  AND2_X1 _31182_ (
    .A1(_00008_[1]),
    .A2(_23061_),
    .ZN(_23062_)
  );
  INV_X1 _31183_ (
    .A(_23062_),
    .ZN(_23063_)
  );
  AND2_X1 _31184_ (
    .A1(_21462_),
    .A2(_22149_),
    .ZN(_23064_)
  );
  INV_X1 _31185_ (
    .A(_23064_),
    .ZN(_23065_)
  );
  AND2_X1 _31186_ (
    .A1(_21761_),
    .A2(_00008_[2]),
    .ZN(_23066_)
  );
  INV_X1 _31187_ (
    .A(_23066_),
    .ZN(_23067_)
  );
  AND2_X1 _31188_ (
    .A1(_21440_),
    .A2(_22149_),
    .ZN(_23068_)
  );
  INV_X1 _31189_ (
    .A(_23068_),
    .ZN(_23069_)
  );
  AND2_X1 _31190_ (
    .A1(_21651_),
    .A2(_00008_[2]),
    .ZN(_23070_)
  );
  INV_X1 _31191_ (
    .A(_23070_),
    .ZN(_23071_)
  );
  AND2_X1 _31192_ (
    .A1(_23069_),
    .A2(_23071_),
    .ZN(_23072_)
  );
  AND2_X1 _31193_ (
    .A1(_00008_[0]),
    .A2(_23065_),
    .ZN(_23073_)
  );
  AND2_X1 _31194_ (
    .A1(_23067_),
    .A2(_23073_),
    .ZN(_23074_)
  );
  INV_X1 _31195_ (
    .A(_23074_),
    .ZN(_23075_)
  );
  AND2_X1 _31196_ (
    .A1(_22147_),
    .A2(_23072_),
    .ZN(_23076_)
  );
  INV_X1 _31197_ (
    .A(_23076_),
    .ZN(_23077_)
  );
  AND2_X1 _31198_ (
    .A1(_23075_),
    .A2(_23077_),
    .ZN(_23078_)
  );
  AND2_X1 _31199_ (
    .A1(_22148_),
    .A2(_23078_),
    .ZN(_23079_)
  );
  INV_X1 _31200_ (
    .A(_23079_),
    .ZN(_23080_)
  );
  AND2_X1 _31201_ (
    .A1(_23063_),
    .A2(_23080_),
    .ZN(_23081_)
  );
  AND2_X1 _31202_ (
    .A1(_22150_),
    .A2(_23081_),
    .ZN(_23082_)
  );
  INV_X1 _31203_ (
    .A(_23082_),
    .ZN(_23083_)
  );
  AND2_X1 _31204_ (
    .A1(_00008_[3]),
    .A2(_23046_),
    .ZN(_23084_)
  );
  AND2_X1 _31205_ (
    .A1(_23028_),
    .A2(_23084_),
    .ZN(_23085_)
  );
  INV_X1 _31206_ (
    .A(_23085_),
    .ZN(_23086_)
  );
  AND2_X1 _31207_ (
    .A1(_00008_[4]),
    .A2(_23086_),
    .ZN(_23087_)
  );
  AND2_X1 _31208_ (
    .A1(_23083_),
    .A2(_23087_),
    .ZN(_23088_)
  );
  INV_X1 _31209_ (
    .A(_23088_),
    .ZN(_23089_)
  );
  AND2_X1 _31210_ (
    .A1(_21783_),
    .A2(_00008_[2]),
    .ZN(_23090_)
  );
  INV_X1 _31211_ (
    .A(_23090_),
    .ZN(_23091_)
  );
  AND2_X1 _31212_ (
    .A1(_21491_),
    .A2(_22149_),
    .ZN(_23092_)
  );
  INV_X1 _31213_ (
    .A(_23092_),
    .ZN(_23093_)
  );
  AND2_X1 _31214_ (
    .A1(_21541_),
    .A2(_22149_),
    .ZN(_23094_)
  );
  INV_X1 _31215_ (
    .A(_23094_),
    .ZN(_23095_)
  );
  AND2_X1 _31216_ (
    .A1(_21808_),
    .A2(_00008_[2]),
    .ZN(_23096_)
  );
  INV_X1 _31217_ (
    .A(_23096_),
    .ZN(_23097_)
  );
  AND2_X1 _31218_ (
    .A1(_23095_),
    .A2(_23097_),
    .ZN(_23098_)
  );
  AND2_X1 _31219_ (
    .A1(_00008_[0]),
    .A2(_23093_),
    .ZN(_23099_)
  );
  AND2_X1 _31220_ (
    .A1(_23091_),
    .A2(_23099_),
    .ZN(_23100_)
  );
  INV_X1 _31221_ (
    .A(_23100_),
    .ZN(_23101_)
  );
  AND2_X1 _31222_ (
    .A1(_22147_),
    .A2(_23098_),
    .ZN(_23102_)
  );
  INV_X1 _31223_ (
    .A(_23102_),
    .ZN(_23103_)
  );
  AND2_X1 _31224_ (
    .A1(_23101_),
    .A2(_23103_),
    .ZN(_23104_)
  );
  AND2_X1 _31225_ (
    .A1(_00008_[1]),
    .A2(_23104_),
    .ZN(_23105_)
  );
  INV_X1 _31226_ (
    .A(_23105_),
    .ZN(_23106_)
  );
  AND2_X1 _31227_ (
    .A1(_21516_),
    .A2(_22149_),
    .ZN(_23107_)
  );
  INV_X1 _31228_ (
    .A(_23107_),
    .ZN(_23108_)
  );
  AND2_X1 _31229_ (
    .A1(_21736_),
    .A2(_00008_[2]),
    .ZN(_23109_)
  );
  INV_X1 _31230_ (
    .A(_23109_),
    .ZN(_23110_)
  );
  AND2_X1 _31231_ (
    .A1(_21957_),
    .A2(_22149_),
    .ZN(_23111_)
  );
  INV_X1 _31232_ (
    .A(_23111_),
    .ZN(_23112_)
  );
  AND2_X1 _31233_ (
    .A1(_21673_),
    .A2(_00008_[2]),
    .ZN(_23113_)
  );
  INV_X1 _31234_ (
    .A(_23113_),
    .ZN(_23114_)
  );
  AND2_X1 _31235_ (
    .A1(_23112_),
    .A2(_23114_),
    .ZN(_23115_)
  );
  AND2_X1 _31236_ (
    .A1(_00008_[0]),
    .A2(_23108_),
    .ZN(_23116_)
  );
  AND2_X1 _31237_ (
    .A1(_23110_),
    .A2(_23116_),
    .ZN(_23117_)
  );
  INV_X1 _31238_ (
    .A(_23117_),
    .ZN(_23118_)
  );
  AND2_X1 _31239_ (
    .A1(_22147_),
    .A2(_23115_),
    .ZN(_23119_)
  );
  INV_X1 _31240_ (
    .A(_23119_),
    .ZN(_23120_)
  );
  AND2_X1 _31241_ (
    .A1(_23118_),
    .A2(_23120_),
    .ZN(_23121_)
  );
  AND2_X1 _31242_ (
    .A1(_22148_),
    .A2(_23121_),
    .ZN(_23122_)
  );
  INV_X1 _31243_ (
    .A(_23122_),
    .ZN(_23123_)
  );
  AND2_X1 _31244_ (
    .A1(_23106_),
    .A2(_23123_),
    .ZN(_23124_)
  );
  INV_X1 _31245_ (
    .A(_23124_),
    .ZN(_23125_)
  );
  AND2_X1 _31246_ (
    .A1(_22150_),
    .A2(_23125_),
    .ZN(_23126_)
  );
  INV_X1 _31247_ (
    .A(_23126_),
    .ZN(_23127_)
  );
  AND2_X1 _31248_ (
    .A1(\cpuregs[9] [4]),
    .A2(_22148_),
    .ZN(_23128_)
  );
  INV_X1 _31249_ (
    .A(_23128_),
    .ZN(_23129_)
  );
  AND2_X1 _31250_ (
    .A1(\cpuregs[11] [4]),
    .A2(_00008_[1]),
    .ZN(_23130_)
  );
  INV_X1 _31251_ (
    .A(_23130_),
    .ZN(_23131_)
  );
  AND2_X1 _31252_ (
    .A1(_22149_),
    .A2(_23131_),
    .ZN(_23132_)
  );
  AND2_X1 _31253_ (
    .A1(_23129_),
    .A2(_23132_),
    .ZN(_23133_)
  );
  INV_X1 _31254_ (
    .A(_23133_),
    .ZN(_23134_)
  );
  AND2_X1 _31255_ (
    .A1(\cpuregs[13] [4]),
    .A2(_22148_),
    .ZN(_23135_)
  );
  INV_X1 _31256_ (
    .A(_23135_),
    .ZN(_23136_)
  );
  AND2_X1 _31257_ (
    .A1(\cpuregs[15] [4]),
    .A2(_00008_[1]),
    .ZN(_23137_)
  );
  INV_X1 _31258_ (
    .A(_23137_),
    .ZN(_23138_)
  );
  AND2_X1 _31259_ (
    .A1(_00008_[2]),
    .A2(_23138_),
    .ZN(_23139_)
  );
  AND2_X1 _31260_ (
    .A1(_23136_),
    .A2(_23139_),
    .ZN(_23140_)
  );
  INV_X1 _31261_ (
    .A(_23140_),
    .ZN(_23141_)
  );
  AND2_X1 _31262_ (
    .A1(_23134_),
    .A2(_23141_),
    .ZN(_23142_)
  );
  INV_X1 _31263_ (
    .A(_23142_),
    .ZN(_23143_)
  );
  AND2_X1 _31264_ (
    .A1(_00008_[0]),
    .A2(_23143_),
    .ZN(_23144_)
  );
  INV_X1 _31265_ (
    .A(_23144_),
    .ZN(_23145_)
  );
  AND2_X1 _31266_ (
    .A1(\cpuregs[8] [4]),
    .A2(_22148_),
    .ZN(_23146_)
  );
  INV_X1 _31267_ (
    .A(_23146_),
    .ZN(_23147_)
  );
  AND2_X1 _31268_ (
    .A1(\cpuregs[10] [4]),
    .A2(_00008_[1]),
    .ZN(_23148_)
  );
  INV_X1 _31269_ (
    .A(_23148_),
    .ZN(_23149_)
  );
  AND2_X1 _31270_ (
    .A1(_22149_),
    .A2(_23149_),
    .ZN(_23150_)
  );
  AND2_X1 _31271_ (
    .A1(_23147_),
    .A2(_23150_),
    .ZN(_23151_)
  );
  INV_X1 _31272_ (
    .A(_23151_),
    .ZN(_23152_)
  );
  AND2_X1 _31273_ (
    .A1(\cpuregs[12] [4]),
    .A2(_22148_),
    .ZN(_23153_)
  );
  INV_X1 _31274_ (
    .A(_23153_),
    .ZN(_23154_)
  );
  AND2_X1 _31275_ (
    .A1(\cpuregs[14] [4]),
    .A2(_00008_[1]),
    .ZN(_23155_)
  );
  INV_X1 _31276_ (
    .A(_23155_),
    .ZN(_23156_)
  );
  AND2_X1 _31277_ (
    .A1(_00008_[2]),
    .A2(_23156_),
    .ZN(_23157_)
  );
  AND2_X1 _31278_ (
    .A1(_23154_),
    .A2(_23157_),
    .ZN(_23158_)
  );
  INV_X1 _31279_ (
    .A(_23158_),
    .ZN(_23159_)
  );
  AND2_X1 _31280_ (
    .A1(_23152_),
    .A2(_23159_),
    .ZN(_23160_)
  );
  INV_X1 _31281_ (
    .A(_23160_),
    .ZN(_23161_)
  );
  AND2_X1 _31282_ (
    .A1(_22147_),
    .A2(_23161_),
    .ZN(_23162_)
  );
  INV_X1 _31283_ (
    .A(_23162_),
    .ZN(_23163_)
  );
  AND2_X1 _31284_ (
    .A1(_23145_),
    .A2(_23163_),
    .ZN(_23164_)
  );
  INV_X1 _31285_ (
    .A(_23164_),
    .ZN(_23165_)
  );
  AND2_X1 _31286_ (
    .A1(_00008_[3]),
    .A2(_23165_),
    .ZN(_23166_)
  );
  INV_X1 _31287_ (
    .A(_23166_),
    .ZN(_23167_)
  );
  AND2_X1 _31288_ (
    .A1(_23127_),
    .A2(_23167_),
    .ZN(_23168_)
  );
  INV_X1 _31289_ (
    .A(_23168_),
    .ZN(_23169_)
  );
  AND2_X1 _31290_ (
    .A1(_22151_),
    .A2(_23169_),
    .ZN(_23170_)
  );
  INV_X1 _31291_ (
    .A(_23170_),
    .ZN(_23171_)
  );
  AND2_X1 _31292_ (
    .A1(_22546_),
    .A2(_23089_),
    .ZN(_23172_)
  );
  AND2_X1 _31293_ (
    .A1(_23171_),
    .A2(_23172_),
    .ZN(_23173_)
  );
  INV_X1 _31294_ (
    .A(_23173_),
    .ZN(_23174_)
  );
  AND2_X1 _31295_ (
    .A1(_23010_),
    .A2(_23174_),
    .ZN(_23175_)
  );
  INV_X1 _31296_ (
    .A(_23175_),
    .ZN(_23176_)
  );
  AND2_X1 _31297_ (
    .A1(_22271_),
    .A2(_23176_),
    .ZN(_23177_)
  );
  INV_X1 _31298_ (
    .A(_23177_),
    .ZN(_23178_)
  );
  AND2_X1 _31299_ (
    .A1(_22989_),
    .A2(_22997_),
    .ZN(_23179_)
  );
  INV_X1 _31300_ (
    .A(_23179_),
    .ZN(_23180_)
  );
  AND2_X1 _31301_ (
    .A1(reg_op1[4]),
    .A2(decoded_imm[4]),
    .ZN(_23181_)
  );
  INV_X1 _31302_ (
    .A(_23181_),
    .ZN(_23182_)
  );
  AND2_X1 _31303_ (
    .A1(_21171_),
    .A2(_22005_),
    .ZN(_23183_)
  );
  INV_X1 _31304_ (
    .A(_23183_),
    .ZN(_23184_)
  );
  AND2_X1 _31305_ (
    .A1(_23182_),
    .A2(_23184_),
    .ZN(_23185_)
  );
  INV_X1 _31306_ (
    .A(_23185_),
    .ZN(_23186_)
  );
  AND2_X1 _31307_ (
    .A1(_23180_),
    .A2(_23185_),
    .ZN(_23187_)
  );
  INV_X1 _31308_ (
    .A(_23187_),
    .ZN(_23188_)
  );
  AND2_X1 _31309_ (
    .A1(_23179_),
    .A2(_23186_),
    .ZN(_23189_)
  );
  INV_X1 _31310_ (
    .A(_23189_),
    .ZN(_23190_)
  );
  AND2_X1 _31311_ (
    .A1(_22559_),
    .A2(_23190_),
    .ZN(_23191_)
  );
  AND2_X1 _31312_ (
    .A1(_23188_),
    .A2(_23191_),
    .ZN(_23192_)
  );
  INV_X1 _31313_ (
    .A(_23192_),
    .ZN(_23193_)
  );
  AND2_X1 _31314_ (
    .A1(reg_op1[3]),
    .A2(_22285_),
    .ZN(_23194_)
  );
  INV_X1 _31315_ (
    .A(_23194_),
    .ZN(_23195_)
  );
  AND2_X1 _31316_ (
    .A1(reg_op1[5]),
    .A2(_22290_),
    .ZN(_23196_)
  );
  INV_X1 _31317_ (
    .A(_23196_),
    .ZN(_23197_)
  );
  AND2_X1 _31318_ (
    .A1(_23195_),
    .A2(_23197_),
    .ZN(_23198_)
  );
  AND2_X1 _31319_ (
    .A1(_22572_),
    .A2(_23198_),
    .ZN(_23199_)
  );
  INV_X1 _31320_ (
    .A(_23199_),
    .ZN(_23200_)
  );
  AND2_X1 _31321_ (
    .A1(reg_op1[0]),
    .A2(_22285_),
    .ZN(_23201_)
  );
  INV_X1 _31322_ (
    .A(_23201_),
    .ZN(_23202_)
  );
  AND2_X1 _31323_ (
    .A1(reg_op1[8]),
    .A2(_22290_),
    .ZN(_23203_)
  );
  INV_X1 _31324_ (
    .A(_23203_),
    .ZN(_23204_)
  );
  AND2_X1 _31325_ (
    .A1(_23202_),
    .A2(_23204_),
    .ZN(_23205_)
  );
  AND2_X1 _31326_ (
    .A1(_22573_),
    .A2(_23205_),
    .ZN(_23206_)
  );
  INV_X1 _31327_ (
    .A(_23206_),
    .ZN(_23207_)
  );
  AND2_X1 _31328_ (
    .A1(_22295_),
    .A2(_23207_),
    .ZN(_23208_)
  );
  AND2_X1 _31329_ (
    .A1(_23200_),
    .A2(_23208_),
    .ZN(_23209_)
  );
  INV_X1 _31330_ (
    .A(_23209_),
    .ZN(_23210_)
  );
  AND2_X1 _31331_ (
    .A1(_22333_),
    .A2(_23210_),
    .ZN(_23211_)
  );
  AND2_X1 _31332_ (
    .A1(_23193_),
    .A2(_23211_),
    .ZN(_23212_)
  );
  AND2_X1 _31333_ (
    .A1(_23178_),
    .A2(_23212_),
    .ZN(_23213_)
  );
  INV_X1 _31334_ (
    .A(_23213_),
    .ZN(_23214_)
  );
  AND2_X1 _31335_ (
    .A1(_23008_),
    .A2(_23214_),
    .ZN(_00061_)
  );
  AND2_X1 _31336_ (
    .A1(_21172_),
    .A2(_22334_),
    .ZN(_23215_)
  );
  INV_X1 _31337_ (
    .A(_23215_),
    .ZN(_23216_)
  );
  AND2_X1 _31338_ (
    .A1(reg_pc[5]),
    .A2(_22335_),
    .ZN(_23217_)
  );
  INV_X1 _31339_ (
    .A(_23217_),
    .ZN(_23218_)
  );
  AND2_X1 _31340_ (
    .A1(_21639_),
    .A2(_00008_[2]),
    .ZN(_23219_)
  );
  INV_X1 _31341_ (
    .A(_23219_),
    .ZN(_23220_)
  );
  AND2_X1 _31342_ (
    .A1(_21717_),
    .A2(_22149_),
    .ZN(_23221_)
  );
  INV_X1 _31343_ (
    .A(_23221_),
    .ZN(_23222_)
  );
  AND2_X1 _31344_ (
    .A1(_00008_[0]),
    .A2(_23220_),
    .ZN(_23223_)
  );
  AND2_X1 _31345_ (
    .A1(_23222_),
    .A2(_23223_),
    .ZN(_23224_)
  );
  INV_X1 _31346_ (
    .A(_23224_),
    .ZN(_23225_)
  );
  AND2_X1 _31347_ (
    .A1(_21725_),
    .A2(_22149_),
    .ZN(_23226_)
  );
  INV_X1 _31348_ (
    .A(_23226_),
    .ZN(_23227_)
  );
  AND2_X1 _31349_ (
    .A1(_21480_),
    .A2(_00008_[2]),
    .ZN(_23228_)
  );
  INV_X1 _31350_ (
    .A(_23228_),
    .ZN(_23229_)
  );
  AND2_X1 _31351_ (
    .A1(_23227_),
    .A2(_23229_),
    .ZN(_23230_)
  );
  AND2_X1 _31352_ (
    .A1(_22147_),
    .A2(_23230_),
    .ZN(_23231_)
  );
  INV_X1 _31353_ (
    .A(_23231_),
    .ZN(_23232_)
  );
  AND2_X1 _31354_ (
    .A1(_23225_),
    .A2(_23232_),
    .ZN(_23233_)
  );
  AND2_X1 _31355_ (
    .A1(_21674_),
    .A2(_00008_[2]),
    .ZN(_23234_)
  );
  INV_X1 _31356_ (
    .A(_23234_),
    .ZN(_23235_)
  );
  AND2_X1 _31357_ (
    .A1(_21958_),
    .A2(_22149_),
    .ZN(_23236_)
  );
  INV_X1 _31358_ (
    .A(_23236_),
    .ZN(_23237_)
  );
  AND2_X1 _31359_ (
    .A1(_23235_),
    .A2(_23237_),
    .ZN(_23238_)
  );
  AND2_X1 _31360_ (
    .A1(_22147_),
    .A2(_23238_),
    .ZN(_23239_)
  );
  INV_X1 _31361_ (
    .A(_23239_),
    .ZN(_23240_)
  );
  AND2_X1 _31362_ (
    .A1(_21737_),
    .A2(_00008_[2]),
    .ZN(_23241_)
  );
  INV_X1 _31363_ (
    .A(_23241_),
    .ZN(_23242_)
  );
  AND2_X1 _31364_ (
    .A1(_21517_),
    .A2(_22149_),
    .ZN(_23243_)
  );
  INV_X1 _31365_ (
    .A(_23243_),
    .ZN(_23244_)
  );
  AND2_X1 _31366_ (
    .A1(_00008_[0]),
    .A2(_23244_),
    .ZN(_23245_)
  );
  AND2_X1 _31367_ (
    .A1(_23242_),
    .A2(_23245_),
    .ZN(_23246_)
  );
  INV_X1 _31368_ (
    .A(_23246_),
    .ZN(_23247_)
  );
  AND2_X1 _31369_ (
    .A1(_23240_),
    .A2(_23247_),
    .ZN(_23248_)
  );
  AND2_X1 _31370_ (
    .A1(_21401_),
    .A2(_00008_[2]),
    .ZN(_23249_)
  );
  INV_X1 _31371_ (
    .A(_23249_),
    .ZN(_23250_)
  );
  AND2_X1 _31372_ (
    .A1(_21583_),
    .A2(_22149_),
    .ZN(_23251_)
  );
  INV_X1 _31373_ (
    .A(_23251_),
    .ZN(_23252_)
  );
  AND2_X1 _31374_ (
    .A1(_00008_[0]),
    .A2(_23250_),
    .ZN(_23253_)
  );
  AND2_X1 _31375_ (
    .A1(_23252_),
    .A2(_23253_),
    .ZN(_23254_)
  );
  INV_X1 _31376_ (
    .A(_23254_),
    .ZN(_23255_)
  );
  AND2_X1 _31377_ (
    .A1(_21698_),
    .A2(_22149_),
    .ZN(_23256_)
  );
  INV_X1 _31378_ (
    .A(_23256_),
    .ZN(_23257_)
  );
  AND2_X1 _31379_ (
    .A1(_21393_),
    .A2(_00008_[2]),
    .ZN(_23258_)
  );
  INV_X1 _31380_ (
    .A(_23258_),
    .ZN(_23259_)
  );
  AND2_X1 _31381_ (
    .A1(_23257_),
    .A2(_23259_),
    .ZN(_23260_)
  );
  AND2_X1 _31382_ (
    .A1(_22147_),
    .A2(_23260_),
    .ZN(_23261_)
  );
  INV_X1 _31383_ (
    .A(_23261_),
    .ZN(_23262_)
  );
  AND2_X1 _31384_ (
    .A1(_23255_),
    .A2(_23262_),
    .ZN(_23263_)
  );
  AND2_X1 _31385_ (
    .A1(_21809_),
    .A2(_00008_[2]),
    .ZN(_23264_)
  );
  INV_X1 _31386_ (
    .A(_23264_),
    .ZN(_23265_)
  );
  AND2_X1 _31387_ (
    .A1(_21542_),
    .A2(_22149_),
    .ZN(_23266_)
  );
  INV_X1 _31388_ (
    .A(_23266_),
    .ZN(_23267_)
  );
  AND2_X1 _31389_ (
    .A1(_23265_),
    .A2(_23267_),
    .ZN(_23268_)
  );
  AND2_X1 _31390_ (
    .A1(_22147_),
    .A2(_23268_),
    .ZN(_23269_)
  );
  INV_X1 _31391_ (
    .A(_23269_),
    .ZN(_23270_)
  );
  AND2_X1 _31392_ (
    .A1(_21784_),
    .A2(_00008_[2]),
    .ZN(_23271_)
  );
  INV_X1 _31393_ (
    .A(_23271_),
    .ZN(_23272_)
  );
  AND2_X1 _31394_ (
    .A1(_21492_),
    .A2(_22149_),
    .ZN(_23273_)
  );
  INV_X1 _31395_ (
    .A(_23273_),
    .ZN(_23274_)
  );
  AND2_X1 _31396_ (
    .A1(_00008_[0]),
    .A2(_23274_),
    .ZN(_23275_)
  );
  AND2_X1 _31397_ (
    .A1(_23272_),
    .A2(_23275_),
    .ZN(_23276_)
  );
  INV_X1 _31398_ (
    .A(_23276_),
    .ZN(_23277_)
  );
  AND2_X1 _31399_ (
    .A1(_23270_),
    .A2(_23277_),
    .ZN(_23278_)
  );
  AND2_X1 _31400_ (
    .A1(_22148_),
    .A2(_23248_),
    .ZN(_23279_)
  );
  INV_X1 _31401_ (
    .A(_23279_),
    .ZN(_23280_)
  );
  AND2_X1 _31402_ (
    .A1(_00008_[1]),
    .A2(_23278_),
    .ZN(_23281_)
  );
  INV_X1 _31403_ (
    .A(_23281_),
    .ZN(_23282_)
  );
  AND2_X1 _31404_ (
    .A1(_23280_),
    .A2(_23282_),
    .ZN(_23283_)
  );
  AND2_X1 _31405_ (
    .A1(_22150_),
    .A2(_23283_),
    .ZN(_23284_)
  );
  INV_X1 _31406_ (
    .A(_23284_),
    .ZN(_23285_)
  );
  AND2_X1 _31407_ (
    .A1(_00008_[1]),
    .A2(_23263_),
    .ZN(_23286_)
  );
  INV_X1 _31408_ (
    .A(_23286_),
    .ZN(_23287_)
  );
  AND2_X1 _31409_ (
    .A1(_22148_),
    .A2(_23233_),
    .ZN(_23288_)
  );
  INV_X1 _31410_ (
    .A(_23288_),
    .ZN(_23289_)
  );
  AND2_X1 _31411_ (
    .A1(_00008_[3]),
    .A2(_23289_),
    .ZN(_23290_)
  );
  AND2_X1 _31412_ (
    .A1(_23287_),
    .A2(_23290_),
    .ZN(_23291_)
  );
  INV_X1 _31413_ (
    .A(_23291_),
    .ZN(_23292_)
  );
  AND2_X1 _31414_ (
    .A1(_22151_),
    .A2(_23292_),
    .ZN(_23293_)
  );
  AND2_X1 _31415_ (
    .A1(_23285_),
    .A2(_23293_),
    .ZN(_23294_)
  );
  INV_X1 _31416_ (
    .A(_23294_),
    .ZN(_23295_)
  );
  AND2_X1 _31417_ (
    .A1(_21375_),
    .A2(_00008_[2]),
    .ZN(_23296_)
  );
  INV_X1 _31418_ (
    .A(_23296_),
    .ZN(_23297_)
  );
  AND2_X1 _31419_ (
    .A1(_21621_),
    .A2(_22149_),
    .ZN(_23298_)
  );
  INV_X1 _31420_ (
    .A(_23298_),
    .ZN(_23299_)
  );
  AND2_X1 _31421_ (
    .A1(_21595_),
    .A2(_22149_),
    .ZN(_23300_)
  );
  INV_X1 _31422_ (
    .A(_23300_),
    .ZN(_23301_)
  );
  AND2_X1 _31423_ (
    .A1(_21413_),
    .A2(_00008_[2]),
    .ZN(_23302_)
  );
  INV_X1 _31424_ (
    .A(_23302_),
    .ZN(_23303_)
  );
  AND2_X1 _31425_ (
    .A1(_23301_),
    .A2(_23303_),
    .ZN(_23304_)
  );
  AND2_X1 _31426_ (
    .A1(_00008_[0]),
    .A2(_23299_),
    .ZN(_23305_)
  );
  AND2_X1 _31427_ (
    .A1(_23297_),
    .A2(_23305_),
    .ZN(_23306_)
  );
  INV_X1 _31428_ (
    .A(_23306_),
    .ZN(_23307_)
  );
  AND2_X1 _31429_ (
    .A1(_22147_),
    .A2(_23304_),
    .ZN(_23308_)
  );
  INV_X1 _31430_ (
    .A(_23308_),
    .ZN(_23309_)
  );
  AND2_X1 _31431_ (
    .A1(_23307_),
    .A2(_23309_),
    .ZN(_23310_)
  );
  AND2_X1 _31432_ (
    .A1(_00008_[1]),
    .A2(_23310_),
    .ZN(_23311_)
  );
  INV_X1 _31433_ (
    .A(_23311_),
    .ZN(_23312_)
  );
  AND2_X1 _31434_ (
    .A1(_21463_),
    .A2(_22149_),
    .ZN(_23313_)
  );
  INV_X1 _31435_ (
    .A(_23313_),
    .ZN(_23314_)
  );
  AND2_X1 _31436_ (
    .A1(_21762_),
    .A2(_00008_[2]),
    .ZN(_23315_)
  );
  INV_X1 _31437_ (
    .A(_23315_),
    .ZN(_23316_)
  );
  AND2_X1 _31438_ (
    .A1(_21441_),
    .A2(_22149_),
    .ZN(_23317_)
  );
  INV_X1 _31439_ (
    .A(_23317_),
    .ZN(_23318_)
  );
  AND2_X1 _31440_ (
    .A1(_21652_),
    .A2(_00008_[2]),
    .ZN(_23319_)
  );
  INV_X1 _31441_ (
    .A(_23319_),
    .ZN(_23320_)
  );
  AND2_X1 _31442_ (
    .A1(_23318_),
    .A2(_23320_),
    .ZN(_23321_)
  );
  AND2_X1 _31443_ (
    .A1(_00008_[0]),
    .A2(_23314_),
    .ZN(_23322_)
  );
  AND2_X1 _31444_ (
    .A1(_23316_),
    .A2(_23322_),
    .ZN(_23323_)
  );
  INV_X1 _31445_ (
    .A(_23323_),
    .ZN(_23324_)
  );
  AND2_X1 _31446_ (
    .A1(_22147_),
    .A2(_23321_),
    .ZN(_23325_)
  );
  INV_X1 _31447_ (
    .A(_23325_),
    .ZN(_23326_)
  );
  AND2_X1 _31448_ (
    .A1(_23324_),
    .A2(_23326_),
    .ZN(_23327_)
  );
  AND2_X1 _31449_ (
    .A1(_22148_),
    .A2(_23327_),
    .ZN(_23328_)
  );
  INV_X1 _31450_ (
    .A(_23328_),
    .ZN(_23329_)
  );
  AND2_X1 _31451_ (
    .A1(_23312_),
    .A2(_23329_),
    .ZN(_23330_)
  );
  AND2_X1 _31452_ (
    .A1(_22150_),
    .A2(_23330_),
    .ZN(_23331_)
  );
  INV_X1 _31453_ (
    .A(_23331_),
    .ZN(_23332_)
  );
  AND2_X1 _31454_ (
    .A1(_21892_),
    .A2(_00008_[2]),
    .ZN(_23333_)
  );
  INV_X1 _31455_ (
    .A(_23333_),
    .ZN(_23334_)
  );
  AND2_X1 _31456_ (
    .A1(_21836_),
    .A2(_22149_),
    .ZN(_23335_)
  );
  INV_X1 _31457_ (
    .A(_23335_),
    .ZN(_23336_)
  );
  AND2_X1 _31458_ (
    .A1(_00008_[0]),
    .A2(_23336_),
    .ZN(_23337_)
  );
  AND2_X1 _31459_ (
    .A1(_23334_),
    .A2(_23337_),
    .ZN(_23338_)
  );
  INV_X1 _31460_ (
    .A(_23338_),
    .ZN(_23339_)
  );
  AND2_X1 _31461_ (
    .A1(_21570_),
    .A2(_22149_),
    .ZN(_23340_)
  );
  INV_X1 _31462_ (
    .A(_23340_),
    .ZN(_23341_)
  );
  AND2_X1 _31463_ (
    .A1(_21908_),
    .A2(_00008_[2]),
    .ZN(_23342_)
  );
  INV_X1 _31464_ (
    .A(_23342_),
    .ZN(_23343_)
  );
  AND2_X1 _31465_ (
    .A1(_23341_),
    .A2(_23343_),
    .ZN(_23344_)
  );
  AND2_X1 _31466_ (
    .A1(_22147_),
    .A2(_23344_),
    .ZN(_23345_)
  );
  INV_X1 _31467_ (
    .A(_23345_),
    .ZN(_23346_)
  );
  AND2_X1 _31468_ (
    .A1(_23339_),
    .A2(_23346_),
    .ZN(_23347_)
  );
  AND2_X1 _31469_ (
    .A1(_22148_),
    .A2(_23347_),
    .ZN(_23348_)
  );
  INV_X1 _31470_ (
    .A(_23348_),
    .ZN(_23349_)
  );
  AND2_X1 _31471_ (
    .A1(_21868_),
    .A2(_22149_),
    .ZN(_23350_)
  );
  INV_X1 _31472_ (
    .A(_23350_),
    .ZN(_23351_)
  );
  AND2_X1 _31473_ (
    .A1(_21852_),
    .A2(_00008_[2]),
    .ZN(_23352_)
  );
  INV_X1 _31474_ (
    .A(_23352_),
    .ZN(_23353_)
  );
  AND2_X1 _31475_ (
    .A1(_23351_),
    .A2(_23353_),
    .ZN(_23354_)
  );
  AND2_X1 _31476_ (
    .A1(_22147_),
    .A2(_23354_),
    .ZN(_23355_)
  );
  INV_X1 _31477_ (
    .A(_23355_),
    .ZN(_23356_)
  );
  AND2_X1 _31478_ (
    .A1(_21940_),
    .A2(_00008_[2]),
    .ZN(_23357_)
  );
  INV_X1 _31479_ (
    .A(_23357_),
    .ZN(_23358_)
  );
  AND2_X1 _31480_ (
    .A1(_21924_),
    .A2(_22149_),
    .ZN(_23359_)
  );
  INV_X1 _31481_ (
    .A(_23359_),
    .ZN(_23360_)
  );
  AND2_X1 _31482_ (
    .A1(_00008_[0]),
    .A2(_23360_),
    .ZN(_23361_)
  );
  AND2_X1 _31483_ (
    .A1(_23358_),
    .A2(_23361_),
    .ZN(_23362_)
  );
  INV_X1 _31484_ (
    .A(_23362_),
    .ZN(_23363_)
  );
  AND2_X1 _31485_ (
    .A1(_23356_),
    .A2(_23363_),
    .ZN(_23364_)
  );
  AND2_X1 _31486_ (
    .A1(_00008_[1]),
    .A2(_23364_),
    .ZN(_23365_)
  );
  INV_X1 _31487_ (
    .A(_23365_),
    .ZN(_23366_)
  );
  AND2_X1 _31488_ (
    .A1(_00008_[3]),
    .A2(_23366_),
    .ZN(_23367_)
  );
  AND2_X1 _31489_ (
    .A1(_23349_),
    .A2(_23367_),
    .ZN(_23368_)
  );
  INV_X1 _31490_ (
    .A(_23368_),
    .ZN(_23369_)
  );
  AND2_X1 _31491_ (
    .A1(_00008_[4]),
    .A2(_23369_),
    .ZN(_23370_)
  );
  AND2_X1 _31492_ (
    .A1(_23332_),
    .A2(_23370_),
    .ZN(_23371_)
  );
  INV_X1 _31493_ (
    .A(_23371_),
    .ZN(_23372_)
  );
  AND2_X1 _31494_ (
    .A1(_22546_),
    .A2(_23295_),
    .ZN(_23373_)
  );
  AND2_X1 _31495_ (
    .A1(_23372_),
    .A2(_23373_),
    .ZN(_23374_)
  );
  INV_X1 _31496_ (
    .A(_23374_),
    .ZN(_23375_)
  );
  AND2_X1 _31497_ (
    .A1(_23218_),
    .A2(_23375_),
    .ZN(_23376_)
  );
  INV_X1 _31498_ (
    .A(_23376_),
    .ZN(_23377_)
  );
  AND2_X1 _31499_ (
    .A1(_22271_),
    .A2(_23377_),
    .ZN(_23378_)
  );
  INV_X1 _31500_ (
    .A(_23378_),
    .ZN(_23379_)
  );
  AND2_X1 _31501_ (
    .A1(_23182_),
    .A2(_23188_),
    .ZN(_23380_)
  );
  INV_X1 _31502_ (
    .A(_23380_),
    .ZN(_23381_)
  );
  AND2_X1 _31503_ (
    .A1(reg_op1[5]),
    .A2(decoded_imm[5]),
    .ZN(_23382_)
  );
  INV_X1 _31504_ (
    .A(_23382_),
    .ZN(_23383_)
  );
  AND2_X1 _31505_ (
    .A1(_21172_),
    .A2(_22004_),
    .ZN(_23384_)
  );
  INV_X1 _31506_ (
    .A(_23384_),
    .ZN(_23385_)
  );
  AND2_X1 _31507_ (
    .A1(_23383_),
    .A2(_23385_),
    .ZN(_23386_)
  );
  INV_X1 _31508_ (
    .A(_23386_),
    .ZN(_23387_)
  );
  AND2_X1 _31509_ (
    .A1(_23380_),
    .A2(_23387_),
    .ZN(_23388_)
  );
  INV_X1 _31510_ (
    .A(_23388_),
    .ZN(_23389_)
  );
  AND2_X1 _31511_ (
    .A1(_23381_),
    .A2(_23386_),
    .ZN(_23390_)
  );
  INV_X1 _31512_ (
    .A(_23390_),
    .ZN(_23391_)
  );
  AND2_X1 _31513_ (
    .A1(reg_op1[9]),
    .A2(_22290_),
    .ZN(_23392_)
  );
  INV_X1 _31514_ (
    .A(_23392_),
    .ZN(_23393_)
  );
  AND2_X1 _31515_ (
    .A1(_22786_),
    .A2(_23393_),
    .ZN(_23394_)
  );
  AND2_X1 _31516_ (
    .A1(_22573_),
    .A2(_23394_),
    .ZN(_23395_)
  );
  INV_X1 _31517_ (
    .A(_23395_),
    .ZN(_23396_)
  );
  AND2_X1 _31518_ (
    .A1(reg_op1[4]),
    .A2(_22285_),
    .ZN(_23397_)
  );
  INV_X1 _31519_ (
    .A(_23397_),
    .ZN(_23398_)
  );
  AND2_X1 _31520_ (
    .A1(_22782_),
    .A2(_23398_),
    .ZN(_23399_)
  );
  AND2_X1 _31521_ (
    .A1(_22572_),
    .A2(_23399_),
    .ZN(_23400_)
  );
  INV_X1 _31522_ (
    .A(_23400_),
    .ZN(_23401_)
  );
  AND2_X1 _31523_ (
    .A1(_22295_),
    .A2(_23401_),
    .ZN(_23402_)
  );
  AND2_X1 _31524_ (
    .A1(_23396_),
    .A2(_23402_),
    .ZN(_23403_)
  );
  INV_X1 _31525_ (
    .A(_23403_),
    .ZN(_23404_)
  );
  AND2_X1 _31526_ (
    .A1(_22559_),
    .A2(_23389_),
    .ZN(_23405_)
  );
  AND2_X1 _31527_ (
    .A1(_23391_),
    .A2(_23405_),
    .ZN(_23406_)
  );
  INV_X1 _31528_ (
    .A(_23406_),
    .ZN(_23407_)
  );
  AND2_X1 _31529_ (
    .A1(_23404_),
    .A2(_23407_),
    .ZN(_23408_)
  );
  AND2_X1 _31530_ (
    .A1(_22333_),
    .A2(_23408_),
    .ZN(_23409_)
  );
  AND2_X1 _31531_ (
    .A1(_23379_),
    .A2(_23409_),
    .ZN(_23410_)
  );
  INV_X1 _31532_ (
    .A(_23410_),
    .ZN(_23411_)
  );
  AND2_X1 _31533_ (
    .A1(_23216_),
    .A2(_23411_),
    .ZN(_00062_)
  );
  AND2_X1 _31534_ (
    .A1(_21173_),
    .A2(_22334_),
    .ZN(_23412_)
  );
  INV_X1 _31535_ (
    .A(_23412_),
    .ZN(_23413_)
  );
  AND2_X1 _31536_ (
    .A1(_23383_),
    .A2(_23391_),
    .ZN(_23414_)
  );
  INV_X1 _31537_ (
    .A(_23414_),
    .ZN(_23415_)
  );
  AND2_X1 _31538_ (
    .A1(reg_op1[6]),
    .A2(decoded_imm[6]),
    .ZN(_23416_)
  );
  INV_X1 _31539_ (
    .A(_23416_),
    .ZN(_23417_)
  );
  AND2_X1 _31540_ (
    .A1(_21173_),
    .A2(_22003_),
    .ZN(_23418_)
  );
  INV_X1 _31541_ (
    .A(_23418_),
    .ZN(_23419_)
  );
  AND2_X1 _31542_ (
    .A1(_23417_),
    .A2(_23419_),
    .ZN(_23420_)
  );
  INV_X1 _31543_ (
    .A(_23420_),
    .ZN(_23421_)
  );
  AND2_X1 _31544_ (
    .A1(_23415_),
    .A2(_23420_),
    .ZN(_23422_)
  );
  INV_X1 _31545_ (
    .A(_23422_),
    .ZN(_23423_)
  );
  AND2_X1 _31546_ (
    .A1(_23414_),
    .A2(_23421_),
    .ZN(_23424_)
  );
  INV_X1 _31547_ (
    .A(_23424_),
    .ZN(_23425_)
  );
  AND2_X1 _31548_ (
    .A1(reg_pc[6]),
    .A2(_22335_),
    .ZN(_23426_)
  );
  INV_X1 _31549_ (
    .A(_23426_),
    .ZN(_23427_)
  );
  AND2_X1 _31550_ (
    .A1(_21699_),
    .A2(_22149_),
    .ZN(_23428_)
  );
  INV_X1 _31551_ (
    .A(_23428_),
    .ZN(_23429_)
  );
  AND2_X1 _31552_ (
    .A1(_21394_),
    .A2(_00008_[2]),
    .ZN(_23430_)
  );
  INV_X1 _31553_ (
    .A(_23430_),
    .ZN(_23431_)
  );
  AND2_X1 _31554_ (
    .A1(_23429_),
    .A2(_23431_),
    .ZN(_23432_)
  );
  AND2_X1 _31555_ (
    .A1(_22147_),
    .A2(_23432_),
    .ZN(_23433_)
  );
  INV_X1 _31556_ (
    .A(_23433_),
    .ZN(_23434_)
  );
  AND2_X1 _31557_ (
    .A1(_21402_),
    .A2(_00008_[2]),
    .ZN(_23435_)
  );
  INV_X1 _31558_ (
    .A(_23435_),
    .ZN(_23436_)
  );
  AND2_X1 _31559_ (
    .A1(_21584_),
    .A2(_22149_),
    .ZN(_23437_)
  );
  INV_X1 _31560_ (
    .A(_23437_),
    .ZN(_23438_)
  );
  AND2_X1 _31561_ (
    .A1(_00008_[0]),
    .A2(_23438_),
    .ZN(_23439_)
  );
  AND2_X1 _31562_ (
    .A1(_23436_),
    .A2(_23439_),
    .ZN(_23440_)
  );
  INV_X1 _31563_ (
    .A(_23440_),
    .ZN(_23441_)
  );
  AND2_X1 _31564_ (
    .A1(_23434_),
    .A2(_23441_),
    .ZN(_23442_)
  );
  AND2_X1 _31565_ (
    .A1(_00008_[1]),
    .A2(_23442_),
    .ZN(_23443_)
  );
  INV_X1 _31566_ (
    .A(_23443_),
    .ZN(_23444_)
  );
  AND2_X1 _31567_ (
    .A1(_21640_),
    .A2(_00008_[2]),
    .ZN(_23445_)
  );
  INV_X1 _31568_ (
    .A(_23445_),
    .ZN(_23446_)
  );
  AND2_X1 _31569_ (
    .A1(_21718_),
    .A2(_22149_),
    .ZN(_23447_)
  );
  INV_X1 _31570_ (
    .A(_23447_),
    .ZN(_23448_)
  );
  AND2_X1 _31571_ (
    .A1(_00008_[0]),
    .A2(_23448_),
    .ZN(_23449_)
  );
  AND2_X1 _31572_ (
    .A1(_23446_),
    .A2(_23449_),
    .ZN(_23450_)
  );
  INV_X1 _31573_ (
    .A(_23450_),
    .ZN(_23451_)
  );
  AND2_X1 _31574_ (
    .A1(_21726_),
    .A2(_22149_),
    .ZN(_23452_)
  );
  INV_X1 _31575_ (
    .A(_23452_),
    .ZN(_23453_)
  );
  AND2_X1 _31576_ (
    .A1(_21481_),
    .A2(_00008_[2]),
    .ZN(_23454_)
  );
  INV_X1 _31577_ (
    .A(_23454_),
    .ZN(_23455_)
  );
  AND2_X1 _31578_ (
    .A1(_23453_),
    .A2(_23455_),
    .ZN(_23456_)
  );
  AND2_X1 _31579_ (
    .A1(_22147_),
    .A2(_23456_),
    .ZN(_23457_)
  );
  INV_X1 _31580_ (
    .A(_23457_),
    .ZN(_23458_)
  );
  AND2_X1 _31581_ (
    .A1(_23451_),
    .A2(_23458_),
    .ZN(_23459_)
  );
  AND2_X1 _31582_ (
    .A1(_22148_),
    .A2(_23459_),
    .ZN(_23460_)
  );
  INV_X1 _31583_ (
    .A(_23460_),
    .ZN(_23461_)
  );
  AND2_X1 _31584_ (
    .A1(_23444_),
    .A2(_23461_),
    .ZN(_23462_)
  );
  AND2_X1 _31585_ (
    .A1(_22151_),
    .A2(_23462_),
    .ZN(_23463_)
  );
  INV_X1 _31586_ (
    .A(_23463_),
    .ZN(_23464_)
  );
  AND2_X1 _31587_ (
    .A1(_21571_),
    .A2(_22149_),
    .ZN(_23465_)
  );
  INV_X1 _31588_ (
    .A(_23465_),
    .ZN(_23466_)
  );
  AND2_X1 _31589_ (
    .A1(_21909_),
    .A2(_00008_[2]),
    .ZN(_23467_)
  );
  INV_X1 _31590_ (
    .A(_23467_),
    .ZN(_23468_)
  );
  AND2_X1 _31591_ (
    .A1(_23466_),
    .A2(_23468_),
    .ZN(_23469_)
  );
  AND2_X1 _31592_ (
    .A1(_22147_),
    .A2(_23469_),
    .ZN(_23470_)
  );
  INV_X1 _31593_ (
    .A(_23470_),
    .ZN(_23471_)
  );
  AND2_X1 _31594_ (
    .A1(_21893_),
    .A2(_00008_[2]),
    .ZN(_23472_)
  );
  INV_X1 _31595_ (
    .A(_23472_),
    .ZN(_23473_)
  );
  AND2_X1 _31596_ (
    .A1(_21837_),
    .A2(_22149_),
    .ZN(_23474_)
  );
  INV_X1 _31597_ (
    .A(_23474_),
    .ZN(_23475_)
  );
  AND2_X1 _31598_ (
    .A1(_00008_[0]),
    .A2(_23475_),
    .ZN(_23476_)
  );
  AND2_X1 _31599_ (
    .A1(_23473_),
    .A2(_23476_),
    .ZN(_23477_)
  );
  INV_X1 _31600_ (
    .A(_23477_),
    .ZN(_23478_)
  );
  AND2_X1 _31601_ (
    .A1(_23471_),
    .A2(_23478_),
    .ZN(_23479_)
  );
  AND2_X1 _31602_ (
    .A1(_22148_),
    .A2(_23479_),
    .ZN(_23480_)
  );
  INV_X1 _31603_ (
    .A(_23480_),
    .ZN(_23481_)
  );
  AND2_X1 _31604_ (
    .A1(_21941_),
    .A2(_00008_[2]),
    .ZN(_23482_)
  );
  INV_X1 _31605_ (
    .A(_23482_),
    .ZN(_23483_)
  );
  AND2_X1 _31606_ (
    .A1(_21925_),
    .A2(_22149_),
    .ZN(_23484_)
  );
  INV_X1 _31607_ (
    .A(_23484_),
    .ZN(_23485_)
  );
  AND2_X1 _31608_ (
    .A1(_00008_[0]),
    .A2(_23485_),
    .ZN(_23486_)
  );
  AND2_X1 _31609_ (
    .A1(_23483_),
    .A2(_23486_),
    .ZN(_23487_)
  );
  INV_X1 _31610_ (
    .A(_23487_),
    .ZN(_23488_)
  );
  AND2_X1 _31611_ (
    .A1(_21869_),
    .A2(_22149_),
    .ZN(_23489_)
  );
  INV_X1 _31612_ (
    .A(_23489_),
    .ZN(_23490_)
  );
  AND2_X1 _31613_ (
    .A1(_21853_),
    .A2(_00008_[2]),
    .ZN(_23491_)
  );
  INV_X1 _31614_ (
    .A(_23491_),
    .ZN(_23492_)
  );
  AND2_X1 _31615_ (
    .A1(_23490_),
    .A2(_23492_),
    .ZN(_23493_)
  );
  AND2_X1 _31616_ (
    .A1(_22147_),
    .A2(_23493_),
    .ZN(_23494_)
  );
  INV_X1 _31617_ (
    .A(_23494_),
    .ZN(_23495_)
  );
  AND2_X1 _31618_ (
    .A1(_23488_),
    .A2(_23495_),
    .ZN(_23496_)
  );
  AND2_X1 _31619_ (
    .A1(_00008_[1]),
    .A2(_23496_),
    .ZN(_23497_)
  );
  INV_X1 _31620_ (
    .A(_23497_),
    .ZN(_23498_)
  );
  AND2_X1 _31621_ (
    .A1(_00008_[4]),
    .A2(_23498_),
    .ZN(_23499_)
  );
  AND2_X1 _31622_ (
    .A1(_23481_),
    .A2(_23499_),
    .ZN(_23500_)
  );
  INV_X1 _31623_ (
    .A(_23500_),
    .ZN(_23501_)
  );
  AND2_X1 _31624_ (
    .A1(_23464_),
    .A2(_23501_),
    .ZN(_23502_)
  );
  AND2_X1 _31625_ (
    .A1(_00008_[3]),
    .A2(_23502_),
    .ZN(_23503_)
  );
  INV_X1 _31626_ (
    .A(_23503_),
    .ZN(_23504_)
  );
  AND2_X1 _31627_ (
    .A1(\cpuregs[17] [6]),
    .A2(_22149_),
    .ZN(_23505_)
  );
  INV_X1 _31628_ (
    .A(_23505_),
    .ZN(_23506_)
  );
  AND2_X1 _31629_ (
    .A1(\cpuregs[21] [6]),
    .A2(_00008_[2]),
    .ZN(_23507_)
  );
  INV_X1 _31630_ (
    .A(_23507_),
    .ZN(_23508_)
  );
  AND2_X1 _31631_ (
    .A1(_22148_),
    .A2(_23508_),
    .ZN(_23509_)
  );
  AND2_X1 _31632_ (
    .A1(_23506_),
    .A2(_23509_),
    .ZN(_23510_)
  );
  INV_X1 _31633_ (
    .A(_23510_),
    .ZN(_23511_)
  );
  AND2_X1 _31634_ (
    .A1(\cpuregs[19] [6]),
    .A2(_22149_),
    .ZN(_23512_)
  );
  INV_X1 _31635_ (
    .A(_23512_),
    .ZN(_23513_)
  );
  AND2_X1 _31636_ (
    .A1(\cpuregs[23] [6]),
    .A2(_00008_[2]),
    .ZN(_23514_)
  );
  INV_X1 _31637_ (
    .A(_23514_),
    .ZN(_23515_)
  );
  AND2_X1 _31638_ (
    .A1(_00008_[1]),
    .A2(_23515_),
    .ZN(_23516_)
  );
  AND2_X1 _31639_ (
    .A1(_23513_),
    .A2(_23516_),
    .ZN(_23517_)
  );
  INV_X1 _31640_ (
    .A(_23517_),
    .ZN(_23518_)
  );
  AND2_X1 _31641_ (
    .A1(_23511_),
    .A2(_23518_),
    .ZN(_23519_)
  );
  INV_X1 _31642_ (
    .A(_23519_),
    .ZN(_23520_)
  );
  AND2_X1 _31643_ (
    .A1(_00008_[0]),
    .A2(_23520_),
    .ZN(_23521_)
  );
  INV_X1 _31644_ (
    .A(_23521_),
    .ZN(_23522_)
  );
  AND2_X1 _31645_ (
    .A1(\cpuregs[16] [6]),
    .A2(_22149_),
    .ZN(_23523_)
  );
  INV_X1 _31646_ (
    .A(_23523_),
    .ZN(_23524_)
  );
  AND2_X1 _31647_ (
    .A1(\cpuregs[20] [6]),
    .A2(_00008_[2]),
    .ZN(_23525_)
  );
  INV_X1 _31648_ (
    .A(_23525_),
    .ZN(_23526_)
  );
  AND2_X1 _31649_ (
    .A1(_22148_),
    .A2(_23526_),
    .ZN(_23527_)
  );
  AND2_X1 _31650_ (
    .A1(_23524_),
    .A2(_23527_),
    .ZN(_23528_)
  );
  INV_X1 _31651_ (
    .A(_23528_),
    .ZN(_23529_)
  );
  AND2_X1 _31652_ (
    .A1(\cpuregs[18] [6]),
    .A2(_22149_),
    .ZN(_23530_)
  );
  INV_X1 _31653_ (
    .A(_23530_),
    .ZN(_23531_)
  );
  AND2_X1 _31654_ (
    .A1(\cpuregs[22] [6]),
    .A2(_00008_[2]),
    .ZN(_23532_)
  );
  INV_X1 _31655_ (
    .A(_23532_),
    .ZN(_23533_)
  );
  AND2_X1 _31656_ (
    .A1(_00008_[1]),
    .A2(_23533_),
    .ZN(_23534_)
  );
  AND2_X1 _31657_ (
    .A1(_23531_),
    .A2(_23534_),
    .ZN(_23535_)
  );
  INV_X1 _31658_ (
    .A(_23535_),
    .ZN(_23536_)
  );
  AND2_X1 _31659_ (
    .A1(_23529_),
    .A2(_23536_),
    .ZN(_23537_)
  );
  INV_X1 _31660_ (
    .A(_23537_),
    .ZN(_23538_)
  );
  AND2_X1 _31661_ (
    .A1(_22147_),
    .A2(_23538_),
    .ZN(_23539_)
  );
  INV_X1 _31662_ (
    .A(_23539_),
    .ZN(_23540_)
  );
  AND2_X1 _31663_ (
    .A1(_23522_),
    .A2(_23540_),
    .ZN(_23541_)
  );
  INV_X1 _31664_ (
    .A(_23541_),
    .ZN(_23542_)
  );
  AND2_X1 _31665_ (
    .A1(_00008_[4]),
    .A2(_23542_),
    .ZN(_23543_)
  );
  INV_X1 _31666_ (
    .A(_23543_),
    .ZN(_23544_)
  );
  AND2_X1 _31667_ (
    .A1(_21785_),
    .A2(_00008_[2]),
    .ZN(_23545_)
  );
  INV_X1 _31668_ (
    .A(_23545_),
    .ZN(_23546_)
  );
  AND2_X1 _31669_ (
    .A1(_21493_),
    .A2(_22149_),
    .ZN(_23547_)
  );
  INV_X1 _31670_ (
    .A(_23547_),
    .ZN(_23548_)
  );
  AND2_X1 _31671_ (
    .A1(_00008_[0]),
    .A2(_23548_),
    .ZN(_23549_)
  );
  AND2_X1 _31672_ (
    .A1(_23546_),
    .A2(_23549_),
    .ZN(_23550_)
  );
  INV_X1 _31673_ (
    .A(_23550_),
    .ZN(_23551_)
  );
  AND2_X1 _31674_ (
    .A1(_21543_),
    .A2(_22149_),
    .ZN(_23552_)
  );
  INV_X1 _31675_ (
    .A(_23552_),
    .ZN(_23553_)
  );
  AND2_X1 _31676_ (
    .A1(_21810_),
    .A2(_00008_[2]),
    .ZN(_23554_)
  );
  INV_X1 _31677_ (
    .A(_23554_),
    .ZN(_23555_)
  );
  AND2_X1 _31678_ (
    .A1(_23553_),
    .A2(_23555_),
    .ZN(_23556_)
  );
  AND2_X1 _31679_ (
    .A1(_22147_),
    .A2(_23556_),
    .ZN(_23557_)
  );
  INV_X1 _31680_ (
    .A(_23557_),
    .ZN(_23558_)
  );
  AND2_X1 _31681_ (
    .A1(_23551_),
    .A2(_23558_),
    .ZN(_23559_)
  );
  AND2_X1 _31682_ (
    .A1(_00008_[1]),
    .A2(_23559_),
    .ZN(_23560_)
  );
  INV_X1 _31683_ (
    .A(_23560_),
    .ZN(_23561_)
  );
  AND2_X1 _31684_ (
    .A1(_21738_),
    .A2(_00008_[2]),
    .ZN(_23562_)
  );
  INV_X1 _31685_ (
    .A(_23562_),
    .ZN(_23563_)
  );
  AND2_X1 _31686_ (
    .A1(_21518_),
    .A2(_22149_),
    .ZN(_23564_)
  );
  INV_X1 _31687_ (
    .A(_23564_),
    .ZN(_23565_)
  );
  AND2_X1 _31688_ (
    .A1(_00008_[0]),
    .A2(_23565_),
    .ZN(_23566_)
  );
  AND2_X1 _31689_ (
    .A1(_23563_),
    .A2(_23566_),
    .ZN(_23567_)
  );
  INV_X1 _31690_ (
    .A(_23567_),
    .ZN(_23568_)
  );
  AND2_X1 _31691_ (
    .A1(_21959_),
    .A2(_22149_),
    .ZN(_23569_)
  );
  INV_X1 _31692_ (
    .A(_23569_),
    .ZN(_23570_)
  );
  AND2_X1 _31693_ (
    .A1(_21675_),
    .A2(_00008_[2]),
    .ZN(_23571_)
  );
  INV_X1 _31694_ (
    .A(_23571_),
    .ZN(_23572_)
  );
  AND2_X1 _31695_ (
    .A1(_23570_),
    .A2(_23572_),
    .ZN(_23573_)
  );
  AND2_X1 _31696_ (
    .A1(_22147_),
    .A2(_23573_),
    .ZN(_23574_)
  );
  INV_X1 _31697_ (
    .A(_23574_),
    .ZN(_23575_)
  );
  AND2_X1 _31698_ (
    .A1(_23568_),
    .A2(_23575_),
    .ZN(_23576_)
  );
  AND2_X1 _31699_ (
    .A1(_22148_),
    .A2(_23576_),
    .ZN(_23577_)
  );
  INV_X1 _31700_ (
    .A(_23577_),
    .ZN(_23578_)
  );
  AND2_X1 _31701_ (
    .A1(_23561_),
    .A2(_23578_),
    .ZN(_23579_)
  );
  INV_X1 _31702_ (
    .A(_23579_),
    .ZN(_23580_)
  );
  AND2_X1 _31703_ (
    .A1(_22151_),
    .A2(_23580_),
    .ZN(_23581_)
  );
  INV_X1 _31704_ (
    .A(_23581_),
    .ZN(_23582_)
  );
  AND2_X1 _31705_ (
    .A1(_23544_),
    .A2(_23582_),
    .ZN(_23583_)
  );
  INV_X1 _31706_ (
    .A(_23583_),
    .ZN(_23584_)
  );
  AND2_X1 _31707_ (
    .A1(_22150_),
    .A2(_23584_),
    .ZN(_23585_)
  );
  INV_X1 _31708_ (
    .A(_23585_),
    .ZN(_23586_)
  );
  AND2_X1 _31709_ (
    .A1(_22546_),
    .A2(_23504_),
    .ZN(_23587_)
  );
  AND2_X1 _31710_ (
    .A1(_23586_),
    .A2(_23587_),
    .ZN(_23588_)
  );
  INV_X1 _31711_ (
    .A(_23588_),
    .ZN(_23589_)
  );
  AND2_X1 _31712_ (
    .A1(_23427_),
    .A2(_23589_),
    .ZN(_23590_)
  );
  INV_X1 _31713_ (
    .A(_23590_),
    .ZN(_23591_)
  );
  AND2_X1 _31714_ (
    .A1(_22271_),
    .A2(_23591_),
    .ZN(_23592_)
  );
  INV_X1 _31715_ (
    .A(_23592_),
    .ZN(_23593_)
  );
  AND2_X1 _31716_ (
    .A1(reg_op1[5]),
    .A2(_22285_),
    .ZN(_23594_)
  );
  INV_X1 _31717_ (
    .A(_23594_),
    .ZN(_23595_)
  );
  AND2_X1 _31718_ (
    .A1(_22980_),
    .A2(_23595_),
    .ZN(_23596_)
  );
  AND2_X1 _31719_ (
    .A1(reg_op1[10]),
    .A2(_22290_),
    .ZN(_23597_)
  );
  INV_X1 _31720_ (
    .A(_23597_),
    .ZN(_23598_)
  );
  AND2_X1 _31721_ (
    .A1(_22975_),
    .A2(_23598_),
    .ZN(_23599_)
  );
  AND2_X1 _31722_ (
    .A1(_22559_),
    .A2(_23423_),
    .ZN(_23600_)
  );
  AND2_X1 _31723_ (
    .A1(_23425_),
    .A2(_23600_),
    .ZN(_23601_)
  );
  INV_X1 _31724_ (
    .A(_23601_),
    .ZN(_23602_)
  );
  AND2_X1 _31725_ (
    .A1(_22573_),
    .A2(_23599_),
    .ZN(_23603_)
  );
  INV_X1 _31726_ (
    .A(_23603_),
    .ZN(_23604_)
  );
  AND2_X1 _31727_ (
    .A1(_22572_),
    .A2(_23596_),
    .ZN(_23605_)
  );
  INV_X1 _31728_ (
    .A(_23605_),
    .ZN(_23606_)
  );
  AND2_X1 _31729_ (
    .A1(_22295_),
    .A2(_23604_),
    .ZN(_23607_)
  );
  AND2_X1 _31730_ (
    .A1(_23606_),
    .A2(_23607_),
    .ZN(_23608_)
  );
  INV_X1 _31731_ (
    .A(_23608_),
    .ZN(_23609_)
  );
  AND2_X1 _31732_ (
    .A1(_23593_),
    .A2(_23609_),
    .ZN(_23610_)
  );
  AND2_X1 _31733_ (
    .A1(_23602_),
    .A2(_23610_),
    .ZN(_23611_)
  );
  AND2_X1 _31734_ (
    .A1(_22333_),
    .A2(_23611_),
    .ZN(_23612_)
  );
  INV_X1 _31735_ (
    .A(_23612_),
    .ZN(_23613_)
  );
  AND2_X1 _31736_ (
    .A1(_23413_),
    .A2(_23613_),
    .ZN(_00063_)
  );
  AND2_X1 _31737_ (
    .A1(_23417_),
    .A2(_23423_),
    .ZN(_23614_)
  );
  INV_X1 _31738_ (
    .A(_23614_),
    .ZN(_23615_)
  );
  AND2_X1 _31739_ (
    .A1(reg_op1[7]),
    .A2(decoded_imm[7]),
    .ZN(_23616_)
  );
  INV_X1 _31740_ (
    .A(_23616_),
    .ZN(_23617_)
  );
  AND2_X1 _31741_ (
    .A1(_21174_),
    .A2(_22002_),
    .ZN(_23618_)
  );
  INV_X1 _31742_ (
    .A(_23618_),
    .ZN(_23619_)
  );
  AND2_X1 _31743_ (
    .A1(_23617_),
    .A2(_23619_),
    .ZN(_23620_)
  );
  INV_X1 _31744_ (
    .A(_23620_),
    .ZN(_23621_)
  );
  AND2_X1 _31745_ (
    .A1(_23614_),
    .A2(_23621_),
    .ZN(_23622_)
  );
  INV_X1 _31746_ (
    .A(_23622_),
    .ZN(_23623_)
  );
  AND2_X1 _31747_ (
    .A1(_23615_),
    .A2(_23620_),
    .ZN(_23624_)
  );
  INV_X1 _31748_ (
    .A(_23624_),
    .ZN(_23625_)
  );
  AND2_X1 _31749_ (
    .A1(_23623_),
    .A2(_23625_),
    .ZN(_23626_)
  );
  AND2_X1 _31750_ (
    .A1(_22559_),
    .A2(_23626_),
    .ZN(_23627_)
  );
  INV_X1 _31751_ (
    .A(_23627_),
    .ZN(_23628_)
  );
  AND2_X1 _31752_ (
    .A1(reg_pc[7]),
    .A2(_22335_),
    .ZN(_23629_)
  );
  INV_X1 _31753_ (
    .A(_23629_),
    .ZN(_23630_)
  );
  AND2_X1 _31754_ (
    .A1(_21700_),
    .A2(_22149_),
    .ZN(_23631_)
  );
  INV_X1 _31755_ (
    .A(_23631_),
    .ZN(_23632_)
  );
  AND2_X1 _31756_ (
    .A1(_21395_),
    .A2(_00008_[2]),
    .ZN(_23633_)
  );
  INV_X1 _31757_ (
    .A(_23633_),
    .ZN(_23634_)
  );
  AND2_X1 _31758_ (
    .A1(_23632_),
    .A2(_23634_),
    .ZN(_23635_)
  );
  AND2_X1 _31759_ (
    .A1(_22147_),
    .A2(_23635_),
    .ZN(_23636_)
  );
  INV_X1 _31760_ (
    .A(_23636_),
    .ZN(_23637_)
  );
  AND2_X1 _31761_ (
    .A1(_21403_),
    .A2(_00008_[2]),
    .ZN(_23638_)
  );
  INV_X1 _31762_ (
    .A(_23638_),
    .ZN(_23639_)
  );
  AND2_X1 _31763_ (
    .A1(_21585_),
    .A2(_22149_),
    .ZN(_23640_)
  );
  INV_X1 _31764_ (
    .A(_23640_),
    .ZN(_23641_)
  );
  AND2_X1 _31765_ (
    .A1(_00008_[0]),
    .A2(_23641_),
    .ZN(_23642_)
  );
  AND2_X1 _31766_ (
    .A1(_23639_),
    .A2(_23642_),
    .ZN(_23643_)
  );
  INV_X1 _31767_ (
    .A(_23643_),
    .ZN(_23644_)
  );
  AND2_X1 _31768_ (
    .A1(_23637_),
    .A2(_23644_),
    .ZN(_23645_)
  );
  AND2_X1 _31769_ (
    .A1(_00008_[1]),
    .A2(_23645_),
    .ZN(_23646_)
  );
  INV_X1 _31770_ (
    .A(_23646_),
    .ZN(_23647_)
  );
  AND2_X1 _31771_ (
    .A1(_21641_),
    .A2(_00008_[2]),
    .ZN(_23648_)
  );
  INV_X1 _31772_ (
    .A(_23648_),
    .ZN(_23649_)
  );
  AND2_X1 _31773_ (
    .A1(_21719_),
    .A2(_22149_),
    .ZN(_23650_)
  );
  INV_X1 _31774_ (
    .A(_23650_),
    .ZN(_23651_)
  );
  AND2_X1 _31775_ (
    .A1(_00008_[0]),
    .A2(_23651_),
    .ZN(_23652_)
  );
  AND2_X1 _31776_ (
    .A1(_23649_),
    .A2(_23652_),
    .ZN(_23653_)
  );
  INV_X1 _31777_ (
    .A(_23653_),
    .ZN(_23654_)
  );
  AND2_X1 _31778_ (
    .A1(_21727_),
    .A2(_22149_),
    .ZN(_23655_)
  );
  INV_X1 _31779_ (
    .A(_23655_),
    .ZN(_23656_)
  );
  AND2_X1 _31780_ (
    .A1(_21482_),
    .A2(_00008_[2]),
    .ZN(_23657_)
  );
  INV_X1 _31781_ (
    .A(_23657_),
    .ZN(_23658_)
  );
  AND2_X1 _31782_ (
    .A1(_23656_),
    .A2(_23658_),
    .ZN(_23659_)
  );
  AND2_X1 _31783_ (
    .A1(_22147_),
    .A2(_23659_),
    .ZN(_23660_)
  );
  INV_X1 _31784_ (
    .A(_23660_),
    .ZN(_23661_)
  );
  AND2_X1 _31785_ (
    .A1(_23654_),
    .A2(_23661_),
    .ZN(_23662_)
  );
  AND2_X1 _31786_ (
    .A1(_22148_),
    .A2(_23662_),
    .ZN(_23663_)
  );
  INV_X1 _31787_ (
    .A(_23663_),
    .ZN(_23664_)
  );
  AND2_X1 _31788_ (
    .A1(_23647_),
    .A2(_23664_),
    .ZN(_23665_)
  );
  AND2_X1 _31789_ (
    .A1(_21786_),
    .A2(_00008_[2]),
    .ZN(_23666_)
  );
  INV_X1 _31790_ (
    .A(_23666_),
    .ZN(_23667_)
  );
  AND2_X1 _31791_ (
    .A1(_21494_),
    .A2(_22149_),
    .ZN(_23668_)
  );
  INV_X1 _31792_ (
    .A(_23668_),
    .ZN(_23669_)
  );
  AND2_X1 _31793_ (
    .A1(_21544_),
    .A2(_22149_),
    .ZN(_23670_)
  );
  INV_X1 _31794_ (
    .A(_23670_),
    .ZN(_23671_)
  );
  AND2_X1 _31795_ (
    .A1(_21811_),
    .A2(_00008_[2]),
    .ZN(_23672_)
  );
  INV_X1 _31796_ (
    .A(_23672_),
    .ZN(_23673_)
  );
  AND2_X1 _31797_ (
    .A1(_23671_),
    .A2(_23673_),
    .ZN(_23674_)
  );
  AND2_X1 _31798_ (
    .A1(_00008_[0]),
    .A2(_23669_),
    .ZN(_23675_)
  );
  AND2_X1 _31799_ (
    .A1(_23667_),
    .A2(_23675_),
    .ZN(_23676_)
  );
  INV_X1 _31800_ (
    .A(_23676_),
    .ZN(_23677_)
  );
  AND2_X1 _31801_ (
    .A1(_22147_),
    .A2(_23674_),
    .ZN(_23678_)
  );
  INV_X1 _31802_ (
    .A(_23678_),
    .ZN(_23679_)
  );
  AND2_X1 _31803_ (
    .A1(_23677_),
    .A2(_23679_),
    .ZN(_23680_)
  );
  AND2_X1 _31804_ (
    .A1(_00008_[1]),
    .A2(_23680_),
    .ZN(_23681_)
  );
  INV_X1 _31805_ (
    .A(_23681_),
    .ZN(_23682_)
  );
  AND2_X1 _31806_ (
    .A1(_21519_),
    .A2(_22149_),
    .ZN(_23683_)
  );
  INV_X1 _31807_ (
    .A(_23683_),
    .ZN(_23684_)
  );
  AND2_X1 _31808_ (
    .A1(_21739_),
    .A2(_00008_[2]),
    .ZN(_23685_)
  );
  INV_X1 _31809_ (
    .A(_23685_),
    .ZN(_23686_)
  );
  AND2_X1 _31810_ (
    .A1(_21960_),
    .A2(_22149_),
    .ZN(_23687_)
  );
  INV_X1 _31811_ (
    .A(_23687_),
    .ZN(_23688_)
  );
  AND2_X1 _31812_ (
    .A1(_21676_),
    .A2(_00008_[2]),
    .ZN(_23689_)
  );
  INV_X1 _31813_ (
    .A(_23689_),
    .ZN(_23690_)
  );
  AND2_X1 _31814_ (
    .A1(_23688_),
    .A2(_23690_),
    .ZN(_23691_)
  );
  AND2_X1 _31815_ (
    .A1(_00008_[0]),
    .A2(_23684_),
    .ZN(_23692_)
  );
  AND2_X1 _31816_ (
    .A1(_23686_),
    .A2(_23692_),
    .ZN(_23693_)
  );
  INV_X1 _31817_ (
    .A(_23693_),
    .ZN(_23694_)
  );
  AND2_X1 _31818_ (
    .A1(_22147_),
    .A2(_23691_),
    .ZN(_23695_)
  );
  INV_X1 _31819_ (
    .A(_23695_),
    .ZN(_23696_)
  );
  AND2_X1 _31820_ (
    .A1(_23694_),
    .A2(_23696_),
    .ZN(_23697_)
  );
  AND2_X1 _31821_ (
    .A1(_22148_),
    .A2(_23697_),
    .ZN(_23698_)
  );
  INV_X1 _31822_ (
    .A(_23698_),
    .ZN(_23699_)
  );
  AND2_X1 _31823_ (
    .A1(_23682_),
    .A2(_23699_),
    .ZN(_23700_)
  );
  AND2_X1 _31824_ (
    .A1(_22151_),
    .A2(_23665_),
    .ZN(_23701_)
  );
  INV_X1 _31825_ (
    .A(_23701_),
    .ZN(_23702_)
  );
  AND2_X1 _31826_ (
    .A1(_21572_),
    .A2(_22149_),
    .ZN(_23703_)
  );
  INV_X1 _31827_ (
    .A(_23703_),
    .ZN(_23704_)
  );
  AND2_X1 _31828_ (
    .A1(_21910_),
    .A2(_00008_[2]),
    .ZN(_23705_)
  );
  INV_X1 _31829_ (
    .A(_23705_),
    .ZN(_23706_)
  );
  AND2_X1 _31830_ (
    .A1(_23704_),
    .A2(_23706_),
    .ZN(_23707_)
  );
  AND2_X1 _31831_ (
    .A1(_22147_),
    .A2(_23707_),
    .ZN(_23708_)
  );
  INV_X1 _31832_ (
    .A(_23708_),
    .ZN(_23709_)
  );
  AND2_X1 _31833_ (
    .A1(_21894_),
    .A2(_00008_[2]),
    .ZN(_23710_)
  );
  INV_X1 _31834_ (
    .A(_23710_),
    .ZN(_23711_)
  );
  AND2_X1 _31835_ (
    .A1(_21838_),
    .A2(_22149_),
    .ZN(_23712_)
  );
  INV_X1 _31836_ (
    .A(_23712_),
    .ZN(_23713_)
  );
  AND2_X1 _31837_ (
    .A1(_00008_[0]),
    .A2(_23713_),
    .ZN(_23714_)
  );
  AND2_X1 _31838_ (
    .A1(_23711_),
    .A2(_23714_),
    .ZN(_23715_)
  );
  INV_X1 _31839_ (
    .A(_23715_),
    .ZN(_23716_)
  );
  AND2_X1 _31840_ (
    .A1(_23709_),
    .A2(_23716_),
    .ZN(_23717_)
  );
  AND2_X1 _31841_ (
    .A1(_22148_),
    .A2(_23717_),
    .ZN(_23718_)
  );
  INV_X1 _31842_ (
    .A(_23718_),
    .ZN(_23719_)
  );
  AND2_X1 _31843_ (
    .A1(_21942_),
    .A2(_00008_[2]),
    .ZN(_23720_)
  );
  INV_X1 _31844_ (
    .A(_23720_),
    .ZN(_23721_)
  );
  AND2_X1 _31845_ (
    .A1(_21926_),
    .A2(_22149_),
    .ZN(_23722_)
  );
  INV_X1 _31846_ (
    .A(_23722_),
    .ZN(_23723_)
  );
  AND2_X1 _31847_ (
    .A1(_00008_[0]),
    .A2(_23723_),
    .ZN(_23724_)
  );
  AND2_X1 _31848_ (
    .A1(_23721_),
    .A2(_23724_),
    .ZN(_23725_)
  );
  INV_X1 _31849_ (
    .A(_23725_),
    .ZN(_23726_)
  );
  AND2_X1 _31850_ (
    .A1(_21870_),
    .A2(_22149_),
    .ZN(_23727_)
  );
  INV_X1 _31851_ (
    .A(_23727_),
    .ZN(_23728_)
  );
  AND2_X1 _31852_ (
    .A1(_21854_),
    .A2(_00008_[2]),
    .ZN(_23729_)
  );
  INV_X1 _31853_ (
    .A(_23729_),
    .ZN(_23730_)
  );
  AND2_X1 _31854_ (
    .A1(_23728_),
    .A2(_23730_),
    .ZN(_23731_)
  );
  AND2_X1 _31855_ (
    .A1(_22147_),
    .A2(_23731_),
    .ZN(_23732_)
  );
  INV_X1 _31856_ (
    .A(_23732_),
    .ZN(_23733_)
  );
  AND2_X1 _31857_ (
    .A1(_23726_),
    .A2(_23733_),
    .ZN(_23734_)
  );
  AND2_X1 _31858_ (
    .A1(_00008_[1]),
    .A2(_23734_),
    .ZN(_23735_)
  );
  INV_X1 _31859_ (
    .A(_23735_),
    .ZN(_23736_)
  );
  AND2_X1 _31860_ (
    .A1(_00008_[4]),
    .A2(_23736_),
    .ZN(_23737_)
  );
  AND2_X1 _31861_ (
    .A1(_23719_),
    .A2(_23737_),
    .ZN(_23738_)
  );
  INV_X1 _31862_ (
    .A(_23738_),
    .ZN(_23739_)
  );
  AND2_X1 _31863_ (
    .A1(_23702_),
    .A2(_23739_),
    .ZN(_23740_)
  );
  AND2_X1 _31864_ (
    .A1(_00008_[3]),
    .A2(_23740_),
    .ZN(_23741_)
  );
  INV_X1 _31865_ (
    .A(_23741_),
    .ZN(_23742_)
  );
  AND2_X1 _31866_ (
    .A1(_22151_),
    .A2(_23700_),
    .ZN(_23743_)
  );
  INV_X1 _31867_ (
    .A(_23743_),
    .ZN(_23744_)
  );
  AND2_X1 _31868_ (
    .A1(_21763_),
    .A2(_00008_[2]),
    .ZN(_23745_)
  );
  INV_X1 _31869_ (
    .A(_23745_),
    .ZN(_23746_)
  );
  AND2_X1 _31870_ (
    .A1(_21464_),
    .A2(_22149_),
    .ZN(_23747_)
  );
  INV_X1 _31871_ (
    .A(_23747_),
    .ZN(_23748_)
  );
  AND2_X1 _31872_ (
    .A1(_00008_[0]),
    .A2(_23748_),
    .ZN(_23749_)
  );
  AND2_X1 _31873_ (
    .A1(_23746_),
    .A2(_23749_),
    .ZN(_23750_)
  );
  INV_X1 _31874_ (
    .A(_23750_),
    .ZN(_23751_)
  );
  AND2_X1 _31875_ (
    .A1(_21442_),
    .A2(_22149_),
    .ZN(_23752_)
  );
  INV_X1 _31876_ (
    .A(_23752_),
    .ZN(_23753_)
  );
  AND2_X1 _31877_ (
    .A1(_21653_),
    .A2(_00008_[2]),
    .ZN(_23754_)
  );
  INV_X1 _31878_ (
    .A(_23754_),
    .ZN(_23755_)
  );
  AND2_X1 _31879_ (
    .A1(_23753_),
    .A2(_23755_),
    .ZN(_23756_)
  );
  AND2_X1 _31880_ (
    .A1(_22147_),
    .A2(_23756_),
    .ZN(_23757_)
  );
  INV_X1 _31881_ (
    .A(_23757_),
    .ZN(_23758_)
  );
  AND2_X1 _31882_ (
    .A1(_23751_),
    .A2(_23758_),
    .ZN(_23759_)
  );
  AND2_X1 _31883_ (
    .A1(_22148_),
    .A2(_23759_),
    .ZN(_23760_)
  );
  INV_X1 _31884_ (
    .A(_23760_),
    .ZN(_23761_)
  );
  AND2_X1 _31885_ (
    .A1(_21376_),
    .A2(_00008_[2]),
    .ZN(_23762_)
  );
  INV_X1 _31886_ (
    .A(_23762_),
    .ZN(_23763_)
  );
  AND2_X1 _31887_ (
    .A1(_21622_),
    .A2(_22149_),
    .ZN(_23764_)
  );
  INV_X1 _31888_ (
    .A(_23764_),
    .ZN(_23765_)
  );
  AND2_X1 _31889_ (
    .A1(_00008_[0]),
    .A2(_23765_),
    .ZN(_23766_)
  );
  AND2_X1 _31890_ (
    .A1(_23763_),
    .A2(_23766_),
    .ZN(_23767_)
  );
  INV_X1 _31891_ (
    .A(_23767_),
    .ZN(_23768_)
  );
  AND2_X1 _31892_ (
    .A1(_21596_),
    .A2(_22149_),
    .ZN(_23769_)
  );
  INV_X1 _31893_ (
    .A(_23769_),
    .ZN(_23770_)
  );
  AND2_X1 _31894_ (
    .A1(_21415_),
    .A2(_00008_[2]),
    .ZN(_23771_)
  );
  INV_X1 _31895_ (
    .A(_23771_),
    .ZN(_23772_)
  );
  AND2_X1 _31896_ (
    .A1(_23770_),
    .A2(_23772_),
    .ZN(_23773_)
  );
  AND2_X1 _31897_ (
    .A1(_22147_),
    .A2(_23773_),
    .ZN(_23774_)
  );
  INV_X1 _31898_ (
    .A(_23774_),
    .ZN(_23775_)
  );
  AND2_X1 _31899_ (
    .A1(_23768_),
    .A2(_23775_),
    .ZN(_23776_)
  );
  AND2_X1 _31900_ (
    .A1(_00008_[1]),
    .A2(_23776_),
    .ZN(_23777_)
  );
  INV_X1 _31901_ (
    .A(_23777_),
    .ZN(_23778_)
  );
  AND2_X1 _31902_ (
    .A1(_00008_[4]),
    .A2(_23778_),
    .ZN(_23779_)
  );
  AND2_X1 _31903_ (
    .A1(_23761_),
    .A2(_23779_),
    .ZN(_23780_)
  );
  INV_X1 _31904_ (
    .A(_23780_),
    .ZN(_23781_)
  );
  AND2_X1 _31905_ (
    .A1(_23744_),
    .A2(_23781_),
    .ZN(_23782_)
  );
  AND2_X1 _31906_ (
    .A1(_22150_),
    .A2(_23782_),
    .ZN(_23783_)
  );
  INV_X1 _31907_ (
    .A(_23783_),
    .ZN(_23784_)
  );
  AND2_X1 _31908_ (
    .A1(_22546_),
    .A2(_23784_),
    .ZN(_23785_)
  );
  AND2_X1 _31909_ (
    .A1(_23742_),
    .A2(_23785_),
    .ZN(_23786_)
  );
  INV_X1 _31910_ (
    .A(_23786_),
    .ZN(_23787_)
  );
  AND2_X1 _31911_ (
    .A1(_23630_),
    .A2(_23787_),
    .ZN(_23788_)
  );
  INV_X1 _31912_ (
    .A(_23788_),
    .ZN(_23789_)
  );
  AND2_X1 _31913_ (
    .A1(_22271_),
    .A2(_23789_),
    .ZN(_23790_)
  );
  INV_X1 _31914_ (
    .A(_23790_),
    .ZN(_23791_)
  );
  AND2_X1 _31915_ (
    .A1(reg_op1[6]),
    .A2(_22285_),
    .ZN(_23792_)
  );
  INV_X1 _31916_ (
    .A(_23792_),
    .ZN(_23793_)
  );
  AND2_X1 _31917_ (
    .A1(_23204_),
    .A2(_23793_),
    .ZN(_23794_)
  );
  AND2_X1 _31918_ (
    .A1(reg_op1[11]),
    .A2(_22290_),
    .ZN(_23795_)
  );
  INV_X1 _31919_ (
    .A(_23795_),
    .ZN(_23796_)
  );
  AND2_X1 _31920_ (
    .A1(_23195_),
    .A2(_23796_),
    .ZN(_23797_)
  );
  AND2_X1 _31921_ (
    .A1(_22573_),
    .A2(_23797_),
    .ZN(_23798_)
  );
  INV_X1 _31922_ (
    .A(_23798_),
    .ZN(_23799_)
  );
  AND2_X1 _31923_ (
    .A1(_22572_),
    .A2(_23794_),
    .ZN(_23800_)
  );
  INV_X1 _31924_ (
    .A(_23800_),
    .ZN(_23801_)
  );
  AND2_X1 _31925_ (
    .A1(_22295_),
    .A2(_23801_),
    .ZN(_23802_)
  );
  AND2_X1 _31926_ (
    .A1(_23799_),
    .A2(_23802_),
    .ZN(_23803_)
  );
  INV_X1 _31927_ (
    .A(_23803_),
    .ZN(_23804_)
  );
  AND2_X1 _31928_ (
    .A1(_22333_),
    .A2(_23804_),
    .ZN(_23805_)
  );
  AND2_X1 _31929_ (
    .A1(_23791_),
    .A2(_23805_),
    .ZN(_23806_)
  );
  AND2_X1 _31930_ (
    .A1(_23628_),
    .A2(_23806_),
    .ZN(_23807_)
  );
  INV_X1 _31931_ (
    .A(_23807_),
    .ZN(_23808_)
  );
  AND2_X1 _31932_ (
    .A1(_21174_),
    .A2(_22334_),
    .ZN(_23809_)
  );
  INV_X1 _31933_ (
    .A(_23809_),
    .ZN(_23810_)
  );
  AND2_X1 _31934_ (
    .A1(_23808_),
    .A2(_23810_),
    .ZN(_00064_)
  );
  AND2_X1 _31935_ (
    .A1(reg_op1[8]),
    .A2(decoded_imm[8]),
    .ZN(_23811_)
  );
  INV_X1 _31936_ (
    .A(_23811_),
    .ZN(_23812_)
  );
  AND2_X1 _31937_ (
    .A1(_21175_),
    .A2(_22001_),
    .ZN(_23813_)
  );
  INV_X1 _31938_ (
    .A(_23813_),
    .ZN(_23814_)
  );
  AND2_X1 _31939_ (
    .A1(_23812_),
    .A2(_23814_),
    .ZN(_23815_)
  );
  INV_X1 _31940_ (
    .A(_23815_),
    .ZN(_23816_)
  );
  AND2_X1 _31941_ (
    .A1(_23615_),
    .A2(_23619_),
    .ZN(_23817_)
  );
  INV_X1 _31942_ (
    .A(_23817_),
    .ZN(_23818_)
  );
  AND2_X1 _31943_ (
    .A1(_23614_),
    .A2(_23617_),
    .ZN(_23819_)
  );
  INV_X1 _31944_ (
    .A(_23819_),
    .ZN(_23820_)
  );
  AND2_X1 _31945_ (
    .A1(_23617_),
    .A2(_23818_),
    .ZN(_23821_)
  );
  AND2_X1 _31946_ (
    .A1(_23619_),
    .A2(_23820_),
    .ZN(_23822_)
  );
  AND2_X1 _31947_ (
    .A1(_23816_),
    .A2(_23821_),
    .ZN(_23823_)
  );
  INV_X1 _31948_ (
    .A(_23823_),
    .ZN(_23824_)
  );
  AND2_X1 _31949_ (
    .A1(_23815_),
    .A2(_23822_),
    .ZN(_23825_)
  );
  INV_X1 _31950_ (
    .A(_23825_),
    .ZN(_23826_)
  );
  AND2_X1 _31951_ (
    .A1(reg_pc[8]),
    .A2(_22335_),
    .ZN(_23827_)
  );
  INV_X1 _31952_ (
    .A(_23827_),
    .ZN(_23828_)
  );
  AND2_X1 _31953_ (
    .A1(\cpuregs[7] [8]),
    .A2(_00008_[2]),
    .ZN(_23829_)
  );
  INV_X1 _31954_ (
    .A(_23829_),
    .ZN(_23830_)
  );
  AND2_X1 _31955_ (
    .A1(\cpuregs[3] [8]),
    .A2(_22149_),
    .ZN(_23831_)
  );
  INV_X1 _31956_ (
    .A(_23831_),
    .ZN(_23832_)
  );
  AND2_X1 _31957_ (
    .A1(_23830_),
    .A2(_23832_),
    .ZN(_23833_)
  );
  AND2_X1 _31958_ (
    .A1(\cpuregs[6] [8]),
    .A2(_00008_[2]),
    .ZN(_23834_)
  );
  INV_X1 _31959_ (
    .A(_23834_),
    .ZN(_23835_)
  );
  AND2_X1 _31960_ (
    .A1(\cpuregs[2] [8]),
    .A2(_22149_),
    .ZN(_23836_)
  );
  INV_X1 _31961_ (
    .A(_23836_),
    .ZN(_23837_)
  );
  AND2_X1 _31962_ (
    .A1(_23835_),
    .A2(_23837_),
    .ZN(_23838_)
  );
  AND2_X1 _31963_ (
    .A1(_22147_),
    .A2(_23838_),
    .ZN(_23839_)
  );
  INV_X1 _31964_ (
    .A(_23839_),
    .ZN(_23840_)
  );
  AND2_X1 _31965_ (
    .A1(_00008_[0]),
    .A2(_23833_),
    .ZN(_23841_)
  );
  INV_X1 _31966_ (
    .A(_23841_),
    .ZN(_23842_)
  );
  AND2_X1 _31967_ (
    .A1(_23840_),
    .A2(_23842_),
    .ZN(_23843_)
  );
  INV_X1 _31968_ (
    .A(_23843_),
    .ZN(_23844_)
  );
  AND2_X1 _31969_ (
    .A1(\cpuregs[4] [8]),
    .A2(_00008_[2]),
    .ZN(_23845_)
  );
  INV_X1 _31970_ (
    .A(_23845_),
    .ZN(_23846_)
  );
  AND2_X1 _31971_ (
    .A1(\cpuregs[0] [8]),
    .A2(_22149_),
    .ZN(_23847_)
  );
  INV_X1 _31972_ (
    .A(_23847_),
    .ZN(_23848_)
  );
  AND2_X1 _31973_ (
    .A1(_23846_),
    .A2(_23848_),
    .ZN(_23849_)
  );
  AND2_X1 _31974_ (
    .A1(_22147_),
    .A2(_23849_),
    .ZN(_23850_)
  );
  INV_X1 _31975_ (
    .A(_23850_),
    .ZN(_23851_)
  );
  AND2_X1 _31976_ (
    .A1(\cpuregs[5] [8]),
    .A2(_00008_[2]),
    .ZN(_23852_)
  );
  INV_X1 _31977_ (
    .A(_23852_),
    .ZN(_23853_)
  );
  AND2_X1 _31978_ (
    .A1(\cpuregs[1] [8]),
    .A2(_22149_),
    .ZN(_23854_)
  );
  INV_X1 _31979_ (
    .A(_23854_),
    .ZN(_23855_)
  );
  AND2_X1 _31980_ (
    .A1(_00008_[0]),
    .A2(_23855_),
    .ZN(_23856_)
  );
  AND2_X1 _31981_ (
    .A1(_23853_),
    .A2(_23856_),
    .ZN(_23857_)
  );
  INV_X1 _31982_ (
    .A(_23857_),
    .ZN(_23858_)
  );
  AND2_X1 _31983_ (
    .A1(_23851_),
    .A2(_23858_),
    .ZN(_23859_)
  );
  INV_X1 _31984_ (
    .A(_23859_),
    .ZN(_23860_)
  );
  AND2_X1 _31985_ (
    .A1(\cpuregs[11] [8]),
    .A2(_22149_),
    .ZN(_23861_)
  );
  INV_X1 _31986_ (
    .A(_23861_),
    .ZN(_23862_)
  );
  AND2_X1 _31987_ (
    .A1(\cpuregs[15] [8]),
    .A2(_00008_[2]),
    .ZN(_23863_)
  );
  INV_X1 _31988_ (
    .A(_23863_),
    .ZN(_23864_)
  );
  AND2_X1 _31989_ (
    .A1(_23862_),
    .A2(_23864_),
    .ZN(_23865_)
  );
  INV_X1 _31990_ (
    .A(_23865_),
    .ZN(_23866_)
  );
  AND2_X1 _31991_ (
    .A1(_00008_[0]),
    .A2(_23866_),
    .ZN(_23867_)
  );
  INV_X1 _31992_ (
    .A(_23867_),
    .ZN(_23868_)
  );
  AND2_X1 _31993_ (
    .A1(\cpuregs[14] [8]),
    .A2(_00008_[2]),
    .ZN(_23869_)
  );
  INV_X1 _31994_ (
    .A(_23869_),
    .ZN(_23870_)
  );
  AND2_X1 _31995_ (
    .A1(\cpuregs[10] [8]),
    .A2(_22149_),
    .ZN(_23871_)
  );
  INV_X1 _31996_ (
    .A(_23871_),
    .ZN(_23872_)
  );
  AND2_X1 _31997_ (
    .A1(_23870_),
    .A2(_23872_),
    .ZN(_23873_)
  );
  INV_X1 _31998_ (
    .A(_23873_),
    .ZN(_23874_)
  );
  AND2_X1 _31999_ (
    .A1(_22147_),
    .A2(_23874_),
    .ZN(_23875_)
  );
  INV_X1 _32000_ (
    .A(_23875_),
    .ZN(_23876_)
  );
  AND2_X1 _32001_ (
    .A1(_23868_),
    .A2(_23876_),
    .ZN(_23877_)
  );
  AND2_X1 _32002_ (
    .A1(_21483_),
    .A2(_00008_[2]),
    .ZN(_23878_)
  );
  INV_X1 _32003_ (
    .A(_23878_),
    .ZN(_23879_)
  );
  AND2_X1 _32004_ (
    .A1(_21728_),
    .A2(_22149_),
    .ZN(_23880_)
  );
  INV_X1 _32005_ (
    .A(_23880_),
    .ZN(_23881_)
  );
  AND2_X1 _32006_ (
    .A1(_23879_),
    .A2(_23881_),
    .ZN(_23882_)
  );
  AND2_X1 _32007_ (
    .A1(_22147_),
    .A2(_23882_),
    .ZN(_23883_)
  );
  INV_X1 _32008_ (
    .A(_23883_),
    .ZN(_23884_)
  );
  AND2_X1 _32009_ (
    .A1(_21720_),
    .A2(_22149_),
    .ZN(_23885_)
  );
  INV_X1 _32010_ (
    .A(_23885_),
    .ZN(_23886_)
  );
  AND2_X1 _32011_ (
    .A1(_21642_),
    .A2(_00008_[2]),
    .ZN(_23887_)
  );
  INV_X1 _32012_ (
    .A(_23887_),
    .ZN(_23888_)
  );
  AND2_X1 _32013_ (
    .A1(_00008_[0]),
    .A2(_23888_),
    .ZN(_23889_)
  );
  AND2_X1 _32014_ (
    .A1(_23886_),
    .A2(_23889_),
    .ZN(_23890_)
  );
  INV_X1 _32015_ (
    .A(_23890_),
    .ZN(_23891_)
  );
  AND2_X1 _32016_ (
    .A1(_23884_),
    .A2(_23891_),
    .ZN(_23892_)
  );
  AND2_X1 _32017_ (
    .A1(_22150_),
    .A2(_23860_),
    .ZN(_23893_)
  );
  INV_X1 _32018_ (
    .A(_23893_),
    .ZN(_23894_)
  );
  AND2_X1 _32019_ (
    .A1(_00008_[3]),
    .A2(_23892_),
    .ZN(_23895_)
  );
  INV_X1 _32020_ (
    .A(_23895_),
    .ZN(_23896_)
  );
  AND2_X1 _32021_ (
    .A1(_22148_),
    .A2(_23896_),
    .ZN(_23897_)
  );
  AND2_X1 _32022_ (
    .A1(_23894_),
    .A2(_23897_),
    .ZN(_23898_)
  );
  INV_X1 _32023_ (
    .A(_23898_),
    .ZN(_23899_)
  );
  AND2_X1 _32024_ (
    .A1(_00008_[3]),
    .A2(_23877_),
    .ZN(_23900_)
  );
  INV_X1 _32025_ (
    .A(_23900_),
    .ZN(_23901_)
  );
  AND2_X1 _32026_ (
    .A1(_22150_),
    .A2(_23844_),
    .ZN(_23902_)
  );
  INV_X1 _32027_ (
    .A(_23902_),
    .ZN(_23903_)
  );
  AND2_X1 _32028_ (
    .A1(_23901_),
    .A2(_23903_),
    .ZN(_23904_)
  );
  AND2_X1 _32029_ (
    .A1(_00008_[1]),
    .A2(_23904_),
    .ZN(_23905_)
  );
  INV_X1 _32030_ (
    .A(_23905_),
    .ZN(_23906_)
  );
  AND2_X1 _32031_ (
    .A1(_22151_),
    .A2(_23906_),
    .ZN(_23907_)
  );
  AND2_X1 _32032_ (
    .A1(_23899_),
    .A2(_23907_),
    .ZN(_23908_)
  );
  INV_X1 _32033_ (
    .A(_23908_),
    .ZN(_23909_)
  );
  AND2_X1 _32034_ (
    .A1(\cpuregs[25] [8]),
    .A2(_22149_),
    .ZN(_23910_)
  );
  INV_X1 _32035_ (
    .A(_23910_),
    .ZN(_23911_)
  );
  AND2_X1 _32036_ (
    .A1(\cpuregs[29] [8]),
    .A2(_00008_[2]),
    .ZN(_23912_)
  );
  INV_X1 _32037_ (
    .A(_23912_),
    .ZN(_23913_)
  );
  AND2_X1 _32038_ (
    .A1(_22148_),
    .A2(_23913_),
    .ZN(_23914_)
  );
  AND2_X1 _32039_ (
    .A1(_23911_),
    .A2(_23914_),
    .ZN(_23915_)
  );
  INV_X1 _32040_ (
    .A(_23915_),
    .ZN(_23916_)
  );
  AND2_X1 _32041_ (
    .A1(\cpuregs[31] [8]),
    .A2(_00008_[2]),
    .ZN(_23917_)
  );
  INV_X1 _32042_ (
    .A(_23917_),
    .ZN(_23918_)
  );
  AND2_X1 _32043_ (
    .A1(\cpuregs[27] [8]),
    .A2(_22149_),
    .ZN(_23919_)
  );
  INV_X1 _32044_ (
    .A(_23919_),
    .ZN(_23920_)
  );
  AND2_X1 _32045_ (
    .A1(_00008_[1]),
    .A2(_23920_),
    .ZN(_23921_)
  );
  AND2_X1 _32046_ (
    .A1(_23918_),
    .A2(_23921_),
    .ZN(_23922_)
  );
  INV_X1 _32047_ (
    .A(_23922_),
    .ZN(_23923_)
  );
  AND2_X1 _32048_ (
    .A1(_23916_),
    .A2(_23923_),
    .ZN(_23924_)
  );
  INV_X1 _32049_ (
    .A(_23924_),
    .ZN(_23925_)
  );
  AND2_X1 _32050_ (
    .A1(_00008_[0]),
    .A2(_23925_),
    .ZN(_23926_)
  );
  INV_X1 _32051_ (
    .A(_23926_),
    .ZN(_23927_)
  );
  AND2_X1 _32052_ (
    .A1(\cpuregs[24] [8]),
    .A2(_22149_),
    .ZN(_23928_)
  );
  INV_X1 _32053_ (
    .A(_23928_),
    .ZN(_23929_)
  );
  AND2_X1 _32054_ (
    .A1(\cpuregs[28] [8]),
    .A2(_00008_[2]),
    .ZN(_23930_)
  );
  INV_X1 _32055_ (
    .A(_23930_),
    .ZN(_23931_)
  );
  AND2_X1 _32056_ (
    .A1(_22148_),
    .A2(_23931_),
    .ZN(_23932_)
  );
  AND2_X1 _32057_ (
    .A1(_23929_),
    .A2(_23932_),
    .ZN(_23933_)
  );
  INV_X1 _32058_ (
    .A(_23933_),
    .ZN(_23934_)
  );
  AND2_X1 _32059_ (
    .A1(\cpuregs[26] [8]),
    .A2(_22149_),
    .ZN(_23935_)
  );
  INV_X1 _32060_ (
    .A(_23935_),
    .ZN(_23936_)
  );
  AND2_X1 _32061_ (
    .A1(\cpuregs[30] [8]),
    .A2(_00008_[2]),
    .ZN(_23937_)
  );
  INV_X1 _32062_ (
    .A(_23937_),
    .ZN(_23938_)
  );
  AND2_X1 _32063_ (
    .A1(_00008_[1]),
    .A2(_23938_),
    .ZN(_23939_)
  );
  AND2_X1 _32064_ (
    .A1(_23936_),
    .A2(_23939_),
    .ZN(_23940_)
  );
  INV_X1 _32065_ (
    .A(_23940_),
    .ZN(_23941_)
  );
  AND2_X1 _32066_ (
    .A1(_23934_),
    .A2(_23941_),
    .ZN(_23942_)
  );
  INV_X1 _32067_ (
    .A(_23942_),
    .ZN(_23943_)
  );
  AND2_X1 _32068_ (
    .A1(_22147_),
    .A2(_23943_),
    .ZN(_23944_)
  );
  INV_X1 _32069_ (
    .A(_23944_),
    .ZN(_23945_)
  );
  AND2_X1 _32070_ (
    .A1(_23927_),
    .A2(_23945_),
    .ZN(_23946_)
  );
  INV_X1 _32071_ (
    .A(_23946_),
    .ZN(_23947_)
  );
  AND2_X1 _32072_ (
    .A1(_00008_[3]),
    .A2(_23947_),
    .ZN(_23948_)
  );
  INV_X1 _32073_ (
    .A(_23948_),
    .ZN(_23949_)
  );
  AND2_X1 _32074_ (
    .A1(\cpuregs[17] [8]),
    .A2(_22148_),
    .ZN(_23950_)
  );
  INV_X1 _32075_ (
    .A(_23950_),
    .ZN(_23951_)
  );
  AND2_X1 _32076_ (
    .A1(\cpuregs[19] [8]),
    .A2(_00008_[1]),
    .ZN(_23952_)
  );
  INV_X1 _32077_ (
    .A(_23952_),
    .ZN(_23953_)
  );
  AND2_X1 _32078_ (
    .A1(_22149_),
    .A2(_23953_),
    .ZN(_23954_)
  );
  AND2_X1 _32079_ (
    .A1(_23951_),
    .A2(_23954_),
    .ZN(_23955_)
  );
  INV_X1 _32080_ (
    .A(_23955_),
    .ZN(_23956_)
  );
  AND2_X1 _32081_ (
    .A1(\cpuregs[21] [8]),
    .A2(_22148_),
    .ZN(_23957_)
  );
  INV_X1 _32082_ (
    .A(_23957_),
    .ZN(_23958_)
  );
  AND2_X1 _32083_ (
    .A1(\cpuregs[23] [8]),
    .A2(_00008_[1]),
    .ZN(_23959_)
  );
  INV_X1 _32084_ (
    .A(_23959_),
    .ZN(_23960_)
  );
  AND2_X1 _32085_ (
    .A1(_00008_[2]),
    .A2(_23960_),
    .ZN(_23961_)
  );
  AND2_X1 _32086_ (
    .A1(_23958_),
    .A2(_23961_),
    .ZN(_23962_)
  );
  INV_X1 _32087_ (
    .A(_23962_),
    .ZN(_23963_)
  );
  AND2_X1 _32088_ (
    .A1(_23956_),
    .A2(_23963_),
    .ZN(_23964_)
  );
  INV_X1 _32089_ (
    .A(_23964_),
    .ZN(_23965_)
  );
  AND2_X1 _32090_ (
    .A1(_00008_[0]),
    .A2(_23965_),
    .ZN(_23966_)
  );
  INV_X1 _32091_ (
    .A(_23966_),
    .ZN(_23967_)
  );
  AND2_X1 _32092_ (
    .A1(\cpuregs[16] [8]),
    .A2(_22148_),
    .ZN(_23968_)
  );
  INV_X1 _32093_ (
    .A(_23968_),
    .ZN(_23969_)
  );
  AND2_X1 _32094_ (
    .A1(\cpuregs[18] [8]),
    .A2(_00008_[1]),
    .ZN(_23970_)
  );
  INV_X1 _32095_ (
    .A(_23970_),
    .ZN(_23971_)
  );
  AND2_X1 _32096_ (
    .A1(_22149_),
    .A2(_23971_),
    .ZN(_23972_)
  );
  AND2_X1 _32097_ (
    .A1(_23969_),
    .A2(_23972_),
    .ZN(_23973_)
  );
  INV_X1 _32098_ (
    .A(_23973_),
    .ZN(_23974_)
  );
  AND2_X1 _32099_ (
    .A1(\cpuregs[20] [8]),
    .A2(_22148_),
    .ZN(_23975_)
  );
  INV_X1 _32100_ (
    .A(_23975_),
    .ZN(_23976_)
  );
  AND2_X1 _32101_ (
    .A1(\cpuregs[22] [8]),
    .A2(_00008_[1]),
    .ZN(_23977_)
  );
  INV_X1 _32102_ (
    .A(_23977_),
    .ZN(_23978_)
  );
  AND2_X1 _32103_ (
    .A1(_00008_[2]),
    .A2(_23978_),
    .ZN(_23979_)
  );
  AND2_X1 _32104_ (
    .A1(_23976_),
    .A2(_23979_),
    .ZN(_23980_)
  );
  INV_X1 _32105_ (
    .A(_23980_),
    .ZN(_23981_)
  );
  AND2_X1 _32106_ (
    .A1(_23974_),
    .A2(_23981_),
    .ZN(_23982_)
  );
  INV_X1 _32107_ (
    .A(_23982_),
    .ZN(_23983_)
  );
  AND2_X1 _32108_ (
    .A1(_22147_),
    .A2(_23983_),
    .ZN(_23984_)
  );
  INV_X1 _32109_ (
    .A(_23984_),
    .ZN(_23985_)
  );
  AND2_X1 _32110_ (
    .A1(_23967_),
    .A2(_23985_),
    .ZN(_23986_)
  );
  INV_X1 _32111_ (
    .A(_23986_),
    .ZN(_23987_)
  );
  AND2_X1 _32112_ (
    .A1(_22150_),
    .A2(_23987_),
    .ZN(_23988_)
  );
  INV_X1 _32113_ (
    .A(_23988_),
    .ZN(_23989_)
  );
  AND2_X1 _32114_ (
    .A1(_23949_),
    .A2(_23989_),
    .ZN(_23990_)
  );
  INV_X1 _32115_ (
    .A(_23990_),
    .ZN(_23991_)
  );
  AND2_X1 _32116_ (
    .A1(_00008_[4]),
    .A2(_23991_),
    .ZN(_23992_)
  );
  INV_X1 _32117_ (
    .A(_23992_),
    .ZN(_23993_)
  );
  AND2_X1 _32118_ (
    .A1(_22546_),
    .A2(_23909_),
    .ZN(_23994_)
  );
  AND2_X1 _32119_ (
    .A1(_23993_),
    .A2(_23994_),
    .ZN(_23995_)
  );
  INV_X1 _32120_ (
    .A(_23995_),
    .ZN(_23996_)
  );
  AND2_X1 _32121_ (
    .A1(_23828_),
    .A2(_23996_),
    .ZN(_23997_)
  );
  INV_X1 _32122_ (
    .A(_23997_),
    .ZN(_23998_)
  );
  AND2_X1 _32123_ (
    .A1(_22271_),
    .A2(_23998_),
    .ZN(_23999_)
  );
  INV_X1 _32124_ (
    .A(_23999_),
    .ZN(_24000_)
  );
  AND2_X1 _32125_ (
    .A1(reg_op1[7]),
    .A2(_22285_),
    .ZN(_24001_)
  );
  INV_X1 _32126_ (
    .A(_24001_),
    .ZN(_24002_)
  );
  AND2_X1 _32127_ (
    .A1(_23393_),
    .A2(_24002_),
    .ZN(_24003_)
  );
  AND2_X1 _32128_ (
    .A1(reg_op1[12]),
    .A2(_22290_),
    .ZN(_24004_)
  );
  INV_X1 _32129_ (
    .A(_24004_),
    .ZN(_24005_)
  );
  AND2_X1 _32130_ (
    .A1(_23398_),
    .A2(_24005_),
    .ZN(_24006_)
  );
  AND2_X1 _32131_ (
    .A1(_21175_),
    .A2(_22334_),
    .ZN(_24007_)
  );
  INV_X1 _32132_ (
    .A(_24007_),
    .ZN(_24008_)
  );
  AND2_X1 _32133_ (
    .A1(_22559_),
    .A2(_23824_),
    .ZN(_24009_)
  );
  AND2_X1 _32134_ (
    .A1(_23826_),
    .A2(_24009_),
    .ZN(_24010_)
  );
  INV_X1 _32135_ (
    .A(_24010_),
    .ZN(_24011_)
  );
  AND2_X1 _32136_ (
    .A1(_22573_),
    .A2(_24006_),
    .ZN(_24012_)
  );
  INV_X1 _32137_ (
    .A(_24012_),
    .ZN(_24013_)
  );
  AND2_X1 _32138_ (
    .A1(_22572_),
    .A2(_24003_),
    .ZN(_24014_)
  );
  INV_X1 _32139_ (
    .A(_24014_),
    .ZN(_24015_)
  );
  AND2_X1 _32140_ (
    .A1(_22295_),
    .A2(_24015_),
    .ZN(_24016_)
  );
  AND2_X1 _32141_ (
    .A1(_24013_),
    .A2(_24016_),
    .ZN(_24017_)
  );
  INV_X1 _32142_ (
    .A(_24017_),
    .ZN(_24018_)
  );
  AND2_X1 _32143_ (
    .A1(_24000_),
    .A2(_24018_),
    .ZN(_24019_)
  );
  AND2_X1 _32144_ (
    .A1(_24011_),
    .A2(_24019_),
    .ZN(_24020_)
  );
  AND2_X1 _32145_ (
    .A1(_22333_),
    .A2(_24020_),
    .ZN(_24021_)
  );
  INV_X1 _32146_ (
    .A(_24021_),
    .ZN(_24022_)
  );
  AND2_X1 _32147_ (
    .A1(_24008_),
    .A2(_24022_),
    .ZN(_00065_)
  );
  AND2_X1 _32148_ (
    .A1(reg_op1[9]),
    .A2(decoded_imm[9]),
    .ZN(_24023_)
  );
  INV_X1 _32149_ (
    .A(_24023_),
    .ZN(_24024_)
  );
  AND2_X1 _32150_ (
    .A1(_21176_),
    .A2(_22000_),
    .ZN(_24025_)
  );
  INV_X1 _32151_ (
    .A(_24025_),
    .ZN(_24026_)
  );
  AND2_X1 _32152_ (
    .A1(_24024_),
    .A2(_24026_),
    .ZN(_24027_)
  );
  INV_X1 _32153_ (
    .A(_24027_),
    .ZN(_24028_)
  );
  AND2_X1 _32154_ (
    .A1(reg_pc[9]),
    .A2(_22335_),
    .ZN(_24029_)
  );
  INV_X1 _32155_ (
    .A(_24029_),
    .ZN(_24030_)
  );
  AND2_X1 _32156_ (
    .A1(_21443_),
    .A2(_22149_),
    .ZN(_24031_)
  );
  INV_X1 _32157_ (
    .A(_24031_),
    .ZN(_24032_)
  );
  AND2_X1 _32158_ (
    .A1(_21654_),
    .A2(_00008_[2]),
    .ZN(_24033_)
  );
  INV_X1 _32159_ (
    .A(_24033_),
    .ZN(_24034_)
  );
  AND2_X1 _32160_ (
    .A1(_24032_),
    .A2(_24034_),
    .ZN(_24035_)
  );
  AND2_X1 _32161_ (
    .A1(_22147_),
    .A2(_24035_),
    .ZN(_24036_)
  );
  INV_X1 _32162_ (
    .A(_24036_),
    .ZN(_24037_)
  );
  AND2_X1 _32163_ (
    .A1(_21764_),
    .A2(_00008_[2]),
    .ZN(_24038_)
  );
  INV_X1 _32164_ (
    .A(_24038_),
    .ZN(_24039_)
  );
  AND2_X1 _32165_ (
    .A1(_21465_),
    .A2(_22149_),
    .ZN(_24040_)
  );
  INV_X1 _32166_ (
    .A(_24040_),
    .ZN(_24041_)
  );
  AND2_X1 _32167_ (
    .A1(_00008_[0]),
    .A2(_24039_),
    .ZN(_24042_)
  );
  AND2_X1 _32168_ (
    .A1(_24041_),
    .A2(_24042_),
    .ZN(_24043_)
  );
  INV_X1 _32169_ (
    .A(_24043_),
    .ZN(_24044_)
  );
  AND2_X1 _32170_ (
    .A1(_24037_),
    .A2(_24044_),
    .ZN(_24045_)
  );
  AND2_X1 _32171_ (
    .A1(_22148_),
    .A2(_24045_),
    .ZN(_24046_)
  );
  INV_X1 _32172_ (
    .A(_24046_),
    .ZN(_24047_)
  );
  AND2_X1 _32173_ (
    .A1(_21597_),
    .A2(_22149_),
    .ZN(_24048_)
  );
  INV_X1 _32174_ (
    .A(_24048_),
    .ZN(_24049_)
  );
  AND2_X1 _32175_ (
    .A1(_21417_),
    .A2(_00008_[2]),
    .ZN(_24050_)
  );
  INV_X1 _32176_ (
    .A(_24050_),
    .ZN(_24051_)
  );
  AND2_X1 _32177_ (
    .A1(_24049_),
    .A2(_24051_),
    .ZN(_24052_)
  );
  AND2_X1 _32178_ (
    .A1(_22147_),
    .A2(_24052_),
    .ZN(_24053_)
  );
  INV_X1 _32179_ (
    .A(_24053_),
    .ZN(_24054_)
  );
  AND2_X1 _32180_ (
    .A1(_21377_),
    .A2(_00008_[2]),
    .ZN(_24055_)
  );
  INV_X1 _32181_ (
    .A(_24055_),
    .ZN(_24056_)
  );
  AND2_X1 _32182_ (
    .A1(_21623_),
    .A2(_22149_),
    .ZN(_24057_)
  );
  INV_X1 _32183_ (
    .A(_24057_),
    .ZN(_24058_)
  );
  AND2_X1 _32184_ (
    .A1(_00008_[0]),
    .A2(_24058_),
    .ZN(_24059_)
  );
  AND2_X1 _32185_ (
    .A1(_24056_),
    .A2(_24059_),
    .ZN(_24060_)
  );
  INV_X1 _32186_ (
    .A(_24060_),
    .ZN(_24061_)
  );
  AND2_X1 _32187_ (
    .A1(_24054_),
    .A2(_24061_),
    .ZN(_24062_)
  );
  AND2_X1 _32188_ (
    .A1(_00008_[1]),
    .A2(_24062_),
    .ZN(_24063_)
  );
  INV_X1 _32189_ (
    .A(_24063_),
    .ZN(_24064_)
  );
  AND2_X1 _32190_ (
    .A1(_24047_),
    .A2(_24064_),
    .ZN(_24065_)
  );
  AND2_X1 _32191_ (
    .A1(_21872_),
    .A2(_22149_),
    .ZN(_24066_)
  );
  INV_X1 _32192_ (
    .A(_24066_),
    .ZN(_24067_)
  );
  AND2_X1 _32193_ (
    .A1(_21855_),
    .A2(_00008_[2]),
    .ZN(_24068_)
  );
  INV_X1 _32194_ (
    .A(_24068_),
    .ZN(_24069_)
  );
  AND2_X1 _32195_ (
    .A1(_24067_),
    .A2(_24069_),
    .ZN(_24070_)
  );
  AND2_X1 _32196_ (
    .A1(_22147_),
    .A2(_24070_),
    .ZN(_24071_)
  );
  INV_X1 _32197_ (
    .A(_24071_),
    .ZN(_24072_)
  );
  AND2_X1 _32198_ (
    .A1(_21943_),
    .A2(_00008_[2]),
    .ZN(_24073_)
  );
  INV_X1 _32199_ (
    .A(_24073_),
    .ZN(_24074_)
  );
  AND2_X1 _32200_ (
    .A1(_21927_),
    .A2(_22149_),
    .ZN(_24075_)
  );
  INV_X1 _32201_ (
    .A(_24075_),
    .ZN(_24076_)
  );
  AND2_X1 _32202_ (
    .A1(_00008_[0]),
    .A2(_24076_),
    .ZN(_24077_)
  );
  AND2_X1 _32203_ (
    .A1(_24074_),
    .A2(_24077_),
    .ZN(_24078_)
  );
  INV_X1 _32204_ (
    .A(_24078_),
    .ZN(_24079_)
  );
  AND2_X1 _32205_ (
    .A1(_24072_),
    .A2(_24079_),
    .ZN(_24080_)
  );
  AND2_X1 _32206_ (
    .A1(_00008_[1]),
    .A2(_24080_),
    .ZN(_24081_)
  );
  INV_X1 _32207_ (
    .A(_24081_),
    .ZN(_24082_)
  );
  AND2_X1 _32208_ (
    .A1(_21895_),
    .A2(_00008_[2]),
    .ZN(_24083_)
  );
  INV_X1 _32209_ (
    .A(_24083_),
    .ZN(_24084_)
  );
  AND2_X1 _32210_ (
    .A1(_21839_),
    .A2(_22149_),
    .ZN(_24085_)
  );
  INV_X1 _32211_ (
    .A(_24085_),
    .ZN(_24086_)
  );
  AND2_X1 _32212_ (
    .A1(_00008_[0]),
    .A2(_24086_),
    .ZN(_24087_)
  );
  AND2_X1 _32213_ (
    .A1(_24084_),
    .A2(_24087_),
    .ZN(_24088_)
  );
  INV_X1 _32214_ (
    .A(_24088_),
    .ZN(_24089_)
  );
  AND2_X1 _32215_ (
    .A1(_21573_),
    .A2(_22149_),
    .ZN(_24090_)
  );
  INV_X1 _32216_ (
    .A(_24090_),
    .ZN(_24091_)
  );
  AND2_X1 _32217_ (
    .A1(_21911_),
    .A2(_00008_[2]),
    .ZN(_24092_)
  );
  INV_X1 _32218_ (
    .A(_24092_),
    .ZN(_24093_)
  );
  AND2_X1 _32219_ (
    .A1(_24091_),
    .A2(_24093_),
    .ZN(_24094_)
  );
  AND2_X1 _32220_ (
    .A1(_22147_),
    .A2(_24094_),
    .ZN(_24095_)
  );
  INV_X1 _32221_ (
    .A(_24095_),
    .ZN(_24096_)
  );
  AND2_X1 _32222_ (
    .A1(_24089_),
    .A2(_24096_),
    .ZN(_24097_)
  );
  AND2_X1 _32223_ (
    .A1(_22148_),
    .A2(_24097_),
    .ZN(_24098_)
  );
  INV_X1 _32224_ (
    .A(_24098_),
    .ZN(_24099_)
  );
  AND2_X1 _32225_ (
    .A1(_00008_[3]),
    .A2(_24082_),
    .ZN(_24100_)
  );
  AND2_X1 _32226_ (
    .A1(_24099_),
    .A2(_24100_),
    .ZN(_24101_)
  );
  INV_X1 _32227_ (
    .A(_24101_),
    .ZN(_24102_)
  );
  AND2_X1 _32228_ (
    .A1(_22150_),
    .A2(_24065_),
    .ZN(_24103_)
  );
  INV_X1 _32229_ (
    .A(_24103_),
    .ZN(_24104_)
  );
  AND2_X1 _32230_ (
    .A1(_00008_[4]),
    .A2(_24104_),
    .ZN(_24105_)
  );
  AND2_X1 _32231_ (
    .A1(_24102_),
    .A2(_24105_),
    .ZN(_24106_)
  );
  INV_X1 _32232_ (
    .A(_24106_),
    .ZN(_24107_)
  );
  AND2_X1 _32233_ (
    .A1(\cpuregs[10] [9]),
    .A2(_22149_),
    .ZN(_24108_)
  );
  INV_X1 _32234_ (
    .A(_24108_),
    .ZN(_24109_)
  );
  AND2_X1 _32235_ (
    .A1(\cpuregs[14] [9]),
    .A2(_00008_[2]),
    .ZN(_24110_)
  );
  INV_X1 _32236_ (
    .A(_24110_),
    .ZN(_24111_)
  );
  AND2_X1 _32237_ (
    .A1(_22147_),
    .A2(_24111_),
    .ZN(_24112_)
  );
  AND2_X1 _32238_ (
    .A1(_24109_),
    .A2(_24112_),
    .ZN(_24113_)
  );
  INV_X1 _32239_ (
    .A(_24113_),
    .ZN(_24114_)
  );
  AND2_X1 _32240_ (
    .A1(\cpuregs[15] [9]),
    .A2(_00008_[2]),
    .ZN(_24115_)
  );
  INV_X1 _32241_ (
    .A(_24115_),
    .ZN(_24116_)
  );
  AND2_X1 _32242_ (
    .A1(\cpuregs[11] [9]),
    .A2(_22149_),
    .ZN(_24117_)
  );
  INV_X1 _32243_ (
    .A(_24117_),
    .ZN(_24118_)
  );
  AND2_X1 _32244_ (
    .A1(_00008_[0]),
    .A2(_24118_),
    .ZN(_24119_)
  );
  AND2_X1 _32245_ (
    .A1(_24116_),
    .A2(_24119_),
    .ZN(_24120_)
  );
  INV_X1 _32246_ (
    .A(_24120_),
    .ZN(_24121_)
  );
  AND2_X1 _32247_ (
    .A1(_24114_),
    .A2(_24121_),
    .ZN(_24122_)
  );
  INV_X1 _32248_ (
    .A(_24122_),
    .ZN(_24123_)
  );
  AND2_X1 _32249_ (
    .A1(_00008_[3]),
    .A2(_24123_),
    .ZN(_24124_)
  );
  INV_X1 _32250_ (
    .A(_24124_),
    .ZN(_24125_)
  );
  AND2_X1 _32251_ (
    .A1(\cpuregs[2] [9]),
    .A2(_22149_),
    .ZN(_24126_)
  );
  INV_X1 _32252_ (
    .A(_24126_),
    .ZN(_24127_)
  );
  AND2_X1 _32253_ (
    .A1(\cpuregs[6] [9]),
    .A2(_00008_[2]),
    .ZN(_24128_)
  );
  INV_X1 _32254_ (
    .A(_24128_),
    .ZN(_24129_)
  );
  AND2_X1 _32255_ (
    .A1(_22147_),
    .A2(_24129_),
    .ZN(_24130_)
  );
  AND2_X1 _32256_ (
    .A1(_24127_),
    .A2(_24130_),
    .ZN(_24131_)
  );
  INV_X1 _32257_ (
    .A(_24131_),
    .ZN(_24132_)
  );
  AND2_X1 _32258_ (
    .A1(\cpuregs[3] [9]),
    .A2(_22149_),
    .ZN(_24133_)
  );
  INV_X1 _32259_ (
    .A(_24133_),
    .ZN(_24134_)
  );
  AND2_X1 _32260_ (
    .A1(\cpuregs[7] [9]),
    .A2(_00008_[2]),
    .ZN(_24135_)
  );
  INV_X1 _32261_ (
    .A(_24135_),
    .ZN(_24136_)
  );
  AND2_X1 _32262_ (
    .A1(_00008_[0]),
    .A2(_24136_),
    .ZN(_24137_)
  );
  AND2_X1 _32263_ (
    .A1(_24134_),
    .A2(_24137_),
    .ZN(_24138_)
  );
  INV_X1 _32264_ (
    .A(_24138_),
    .ZN(_24139_)
  );
  AND2_X1 _32265_ (
    .A1(_24132_),
    .A2(_24139_),
    .ZN(_24140_)
  );
  INV_X1 _32266_ (
    .A(_24140_),
    .ZN(_24141_)
  );
  AND2_X1 _32267_ (
    .A1(_22150_),
    .A2(_24141_),
    .ZN(_24142_)
  );
  INV_X1 _32268_ (
    .A(_24142_),
    .ZN(_24143_)
  );
  AND2_X1 _32269_ (
    .A1(\cpuregs[8] [9]),
    .A2(_22149_),
    .ZN(_24144_)
  );
  INV_X1 _32270_ (
    .A(_24144_),
    .ZN(_24145_)
  );
  AND2_X1 _32271_ (
    .A1(\cpuregs[12] [9]),
    .A2(_00008_[2]),
    .ZN(_24146_)
  );
  INV_X1 _32272_ (
    .A(_24146_),
    .ZN(_24147_)
  );
  AND2_X1 _32273_ (
    .A1(_22147_),
    .A2(_24147_),
    .ZN(_24148_)
  );
  AND2_X1 _32274_ (
    .A1(_24145_),
    .A2(_24148_),
    .ZN(_24149_)
  );
  INV_X1 _32275_ (
    .A(_24149_),
    .ZN(_24150_)
  );
  AND2_X1 _32276_ (
    .A1(\cpuregs[13] [9]),
    .A2(_00008_[2]),
    .ZN(_24151_)
  );
  INV_X1 _32277_ (
    .A(_24151_),
    .ZN(_24152_)
  );
  AND2_X1 _32278_ (
    .A1(\cpuregs[9] [9]),
    .A2(_22149_),
    .ZN(_24153_)
  );
  INV_X1 _32279_ (
    .A(_24153_),
    .ZN(_24154_)
  );
  AND2_X1 _32280_ (
    .A1(_00008_[0]),
    .A2(_24154_),
    .ZN(_24155_)
  );
  AND2_X1 _32281_ (
    .A1(_24152_),
    .A2(_24155_),
    .ZN(_24156_)
  );
  INV_X1 _32282_ (
    .A(_24156_),
    .ZN(_24157_)
  );
  AND2_X1 _32283_ (
    .A1(_24150_),
    .A2(_24157_),
    .ZN(_24158_)
  );
  AND2_X1 _32284_ (
    .A1(\cpuregs[0] [9]),
    .A2(_22149_),
    .ZN(_24159_)
  );
  INV_X1 _32285_ (
    .A(_24159_),
    .ZN(_24160_)
  );
  AND2_X1 _32286_ (
    .A1(\cpuregs[4] [9]),
    .A2(_00008_[2]),
    .ZN(_24161_)
  );
  INV_X1 _32287_ (
    .A(_24161_),
    .ZN(_24162_)
  );
  AND2_X1 _32288_ (
    .A1(_22147_),
    .A2(_24162_),
    .ZN(_24163_)
  );
  AND2_X1 _32289_ (
    .A1(_24160_),
    .A2(_24163_),
    .ZN(_24164_)
  );
  INV_X1 _32290_ (
    .A(_24164_),
    .ZN(_24165_)
  );
  AND2_X1 _32291_ (
    .A1(\cpuregs[1] [9]),
    .A2(_22149_),
    .ZN(_24166_)
  );
  INV_X1 _32292_ (
    .A(_24166_),
    .ZN(_24167_)
  );
  AND2_X1 _32293_ (
    .A1(\cpuregs[5] [9]),
    .A2(_00008_[2]),
    .ZN(_24168_)
  );
  INV_X1 _32294_ (
    .A(_24168_),
    .ZN(_24169_)
  );
  AND2_X1 _32295_ (
    .A1(_00008_[0]),
    .A2(_24169_),
    .ZN(_24170_)
  );
  AND2_X1 _32296_ (
    .A1(_24167_),
    .A2(_24170_),
    .ZN(_24171_)
  );
  INV_X1 _32297_ (
    .A(_24171_),
    .ZN(_24172_)
  );
  AND2_X1 _32298_ (
    .A1(_00008_[3]),
    .A2(_24158_),
    .ZN(_24173_)
  );
  INV_X1 _32299_ (
    .A(_24173_),
    .ZN(_24174_)
  );
  AND2_X1 _32300_ (
    .A1(_22150_),
    .A2(_24172_),
    .ZN(_24175_)
  );
  AND2_X1 _32301_ (
    .A1(_24165_),
    .A2(_24175_),
    .ZN(_24176_)
  );
  INV_X1 _32302_ (
    .A(_24176_),
    .ZN(_24177_)
  );
  AND2_X1 _32303_ (
    .A1(_24174_),
    .A2(_24177_),
    .ZN(_24178_)
  );
  INV_X1 _32304_ (
    .A(_24178_),
    .ZN(_24179_)
  );
  AND2_X1 _32305_ (
    .A1(_22148_),
    .A2(_24179_),
    .ZN(_24180_)
  );
  INV_X1 _32306_ (
    .A(_24180_),
    .ZN(_24181_)
  );
  AND2_X1 _32307_ (
    .A1(_00008_[1]),
    .A2(_24143_),
    .ZN(_24182_)
  );
  AND2_X1 _32308_ (
    .A1(_24125_),
    .A2(_24182_),
    .ZN(_24183_)
  );
  INV_X1 _32309_ (
    .A(_24183_),
    .ZN(_24184_)
  );
  AND2_X1 _32310_ (
    .A1(_22151_),
    .A2(_24184_),
    .ZN(_24185_)
  );
  AND2_X1 _32311_ (
    .A1(_24181_),
    .A2(_24185_),
    .ZN(_24186_)
  );
  INV_X1 _32312_ (
    .A(_24186_),
    .ZN(_24187_)
  );
  AND2_X1 _32313_ (
    .A1(_22546_),
    .A2(_24107_),
    .ZN(_24188_)
  );
  AND2_X1 _32314_ (
    .A1(_24187_),
    .A2(_24188_),
    .ZN(_24189_)
  );
  INV_X1 _32315_ (
    .A(_24189_),
    .ZN(_24190_)
  );
  AND2_X1 _32316_ (
    .A1(_24030_),
    .A2(_24190_),
    .ZN(_24191_)
  );
  INV_X1 _32317_ (
    .A(_24191_),
    .ZN(_24192_)
  );
  AND2_X1 _32318_ (
    .A1(_22271_),
    .A2(_24192_),
    .ZN(_24193_)
  );
  INV_X1 _32319_ (
    .A(_24193_),
    .ZN(_24194_)
  );
  AND2_X1 _32320_ (
    .A1(reg_op1[8]),
    .A2(_22285_),
    .ZN(_24195_)
  );
  INV_X1 _32321_ (
    .A(_24195_),
    .ZN(_24196_)
  );
  AND2_X1 _32322_ (
    .A1(_23598_),
    .A2(_24196_),
    .ZN(_24197_)
  );
  AND2_X1 _32323_ (
    .A1(reg_op1[13]),
    .A2(_22290_),
    .ZN(_24198_)
  );
  INV_X1 _32324_ (
    .A(_24198_),
    .ZN(_24199_)
  );
  AND2_X1 _32325_ (
    .A1(_23595_),
    .A2(_24199_),
    .ZN(_24200_)
  );
  AND2_X1 _32326_ (
    .A1(_21176_),
    .A2(_22334_),
    .ZN(_24201_)
  );
  INV_X1 _32327_ (
    .A(_24201_),
    .ZN(_24202_)
  );
  AND2_X1 _32328_ (
    .A1(_23812_),
    .A2(_24028_),
    .ZN(_24203_)
  );
  AND2_X1 _32329_ (
    .A1(_23826_),
    .A2(_24203_),
    .ZN(_24204_)
  );
  INV_X1 _32330_ (
    .A(_24204_),
    .ZN(_24205_)
  );
  AND2_X1 _32331_ (
    .A1(_23825_),
    .A2(_24027_),
    .ZN(_24206_)
  );
  INV_X1 _32332_ (
    .A(_24206_),
    .ZN(_24207_)
  );
  AND2_X1 _32333_ (
    .A1(_23811_),
    .A2(_24027_),
    .ZN(_24208_)
  );
  INV_X1 _32334_ (
    .A(_24208_),
    .ZN(_24209_)
  );
  AND2_X1 _32335_ (
    .A1(_22559_),
    .A2(_24209_),
    .ZN(_24210_)
  );
  AND2_X1 _32336_ (
    .A1(_24207_),
    .A2(_24210_),
    .ZN(_24211_)
  );
  AND2_X1 _32337_ (
    .A1(_24205_),
    .A2(_24211_),
    .ZN(_24212_)
  );
  INV_X1 _32338_ (
    .A(_24212_),
    .ZN(_24213_)
  );
  AND2_X1 _32339_ (
    .A1(_22573_),
    .A2(_24200_),
    .ZN(_24214_)
  );
  INV_X1 _32340_ (
    .A(_24214_),
    .ZN(_24215_)
  );
  AND2_X1 _32341_ (
    .A1(_22572_),
    .A2(_24197_),
    .ZN(_24216_)
  );
  INV_X1 _32342_ (
    .A(_24216_),
    .ZN(_24217_)
  );
  AND2_X1 _32343_ (
    .A1(_22295_),
    .A2(_24217_),
    .ZN(_24218_)
  );
  AND2_X1 _32344_ (
    .A1(_24215_),
    .A2(_24218_),
    .ZN(_24219_)
  );
  INV_X1 _32345_ (
    .A(_24219_),
    .ZN(_24220_)
  );
  AND2_X1 _32346_ (
    .A1(_24194_),
    .A2(_24220_),
    .ZN(_24221_)
  );
  AND2_X1 _32347_ (
    .A1(_24213_),
    .A2(_24221_),
    .ZN(_24222_)
  );
  AND2_X1 _32348_ (
    .A1(_22333_),
    .A2(_24222_),
    .ZN(_24223_)
  );
  INV_X1 _32349_ (
    .A(_24223_),
    .ZN(_24224_)
  );
  AND2_X1 _32350_ (
    .A1(_24202_),
    .A2(_24224_),
    .ZN(_00066_)
  );
  AND2_X1 _32351_ (
    .A1(_21177_),
    .A2(_22334_),
    .ZN(_24225_)
  );
  INV_X1 _32352_ (
    .A(_24225_),
    .ZN(_24226_)
  );
  AND2_X1 _32353_ (
    .A1(reg_pc[10]),
    .A2(_22335_),
    .ZN(_24227_)
  );
  INV_X1 _32354_ (
    .A(_24227_),
    .ZN(_24228_)
  );
  AND2_X1 _32355_ (
    .A1(_21547_),
    .A2(_22149_),
    .ZN(_24229_)
  );
  INV_X1 _32356_ (
    .A(_24229_),
    .ZN(_24230_)
  );
  AND2_X1 _32357_ (
    .A1(_21813_),
    .A2(_00008_[2]),
    .ZN(_24231_)
  );
  INV_X1 _32358_ (
    .A(_24231_),
    .ZN(_24232_)
  );
  AND2_X1 _32359_ (
    .A1(_24230_),
    .A2(_24232_),
    .ZN(_24233_)
  );
  AND2_X1 _32360_ (
    .A1(_22147_),
    .A2(_24233_),
    .ZN(_24234_)
  );
  INV_X1 _32361_ (
    .A(_24234_),
    .ZN(_24235_)
  );
  AND2_X1 _32362_ (
    .A1(\cpuregs[7] [10]),
    .A2(_00008_[2]),
    .ZN(_24236_)
  );
  INV_X1 _32363_ (
    .A(_24236_),
    .ZN(_24237_)
  );
  AND2_X1 _32364_ (
    .A1(\cpuregs[3] [10]),
    .A2(_22149_),
    .ZN(_24238_)
  );
  INV_X1 _32365_ (
    .A(_24238_),
    .ZN(_24239_)
  );
  AND2_X1 _32366_ (
    .A1(_24237_),
    .A2(_24239_),
    .ZN(_24240_)
  );
  INV_X1 _32367_ (
    .A(_24240_),
    .ZN(_24241_)
  );
  AND2_X1 _32368_ (
    .A1(_00008_[0]),
    .A2(_24241_),
    .ZN(_24242_)
  );
  INV_X1 _32369_ (
    .A(_24242_),
    .ZN(_24243_)
  );
  AND2_X1 _32370_ (
    .A1(\cpuregs[5] [10]),
    .A2(_00008_[2]),
    .ZN(_24244_)
  );
  INV_X1 _32371_ (
    .A(_24244_),
    .ZN(_24245_)
  );
  AND2_X1 _32372_ (
    .A1(\cpuregs[1] [10]),
    .A2(_22149_),
    .ZN(_24246_)
  );
  INV_X1 _32373_ (
    .A(_24246_),
    .ZN(_24247_)
  );
  AND2_X1 _32374_ (
    .A1(_24245_),
    .A2(_24247_),
    .ZN(_24248_)
  );
  INV_X1 _32375_ (
    .A(_24248_),
    .ZN(_24249_)
  );
  AND2_X1 _32376_ (
    .A1(_00008_[0]),
    .A2(_24249_),
    .ZN(_24250_)
  );
  INV_X1 _32377_ (
    .A(_24250_),
    .ZN(_24251_)
  );
  AND2_X1 _32378_ (
    .A1(\cpuregs[4] [10]),
    .A2(_00008_[2]),
    .ZN(_24252_)
  );
  INV_X1 _32379_ (
    .A(_24252_),
    .ZN(_24253_)
  );
  AND2_X1 _32380_ (
    .A1(\cpuregs[0] [10]),
    .A2(_22149_),
    .ZN(_24254_)
  );
  INV_X1 _32381_ (
    .A(_24254_),
    .ZN(_24255_)
  );
  AND2_X1 _32382_ (
    .A1(_24253_),
    .A2(_24255_),
    .ZN(_24256_)
  );
  INV_X1 _32383_ (
    .A(_24256_),
    .ZN(_24257_)
  );
  AND2_X1 _32384_ (
    .A1(_22147_),
    .A2(_24257_),
    .ZN(_24258_)
  );
  INV_X1 _32385_ (
    .A(_24258_),
    .ZN(_24259_)
  );
  AND2_X1 _32386_ (
    .A1(_24251_),
    .A2(_24259_),
    .ZN(_24260_)
  );
  AND2_X1 _32387_ (
    .A1(_00008_[1]),
    .A2(_24235_),
    .ZN(_24261_)
  );
  AND2_X1 _32388_ (
    .A1(_24243_),
    .A2(_24261_),
    .ZN(_24262_)
  );
  INV_X1 _32389_ (
    .A(_24262_),
    .ZN(_24263_)
  );
  AND2_X1 _32390_ (
    .A1(_22148_),
    .A2(_24260_),
    .ZN(_24264_)
  );
  INV_X1 _32391_ (
    .A(_24264_),
    .ZN(_24265_)
  );
  AND2_X1 _32392_ (
    .A1(_24263_),
    .A2(_24265_),
    .ZN(_24266_)
  );
  AND2_X1 _32393_ (
    .A1(_22151_),
    .A2(_24266_),
    .ZN(_24267_)
  );
  INV_X1 _32394_ (
    .A(_24267_),
    .ZN(_24268_)
  );
  AND2_X1 _32395_ (
    .A1(_21378_),
    .A2(_00008_[2]),
    .ZN(_24269_)
  );
  INV_X1 _32396_ (
    .A(_24269_),
    .ZN(_24270_)
  );
  AND2_X1 _32397_ (
    .A1(_21624_),
    .A2(_22149_),
    .ZN(_24271_)
  );
  INV_X1 _32398_ (
    .A(_24271_),
    .ZN(_24272_)
  );
  AND2_X1 _32399_ (
    .A1(_00008_[0]),
    .A2(_24272_),
    .ZN(_24273_)
  );
  AND2_X1 _32400_ (
    .A1(_24270_),
    .A2(_24273_),
    .ZN(_24274_)
  );
  INV_X1 _32401_ (
    .A(_24274_),
    .ZN(_24275_)
  );
  AND2_X1 _32402_ (
    .A1(_21598_),
    .A2(_22149_),
    .ZN(_24276_)
  );
  INV_X1 _32403_ (
    .A(_24276_),
    .ZN(_24277_)
  );
  AND2_X1 _32404_ (
    .A1(_21418_),
    .A2(_00008_[2]),
    .ZN(_24278_)
  );
  INV_X1 _32405_ (
    .A(_24278_),
    .ZN(_24279_)
  );
  AND2_X1 _32406_ (
    .A1(_24277_),
    .A2(_24279_),
    .ZN(_24280_)
  );
  AND2_X1 _32407_ (
    .A1(_22147_),
    .A2(_24280_),
    .ZN(_24281_)
  );
  INV_X1 _32408_ (
    .A(_24281_),
    .ZN(_24282_)
  );
  AND2_X1 _32409_ (
    .A1(_24275_),
    .A2(_24282_),
    .ZN(_24283_)
  );
  AND2_X1 _32410_ (
    .A1(_21765_),
    .A2(_00008_[2]),
    .ZN(_24284_)
  );
  INV_X1 _32411_ (
    .A(_24284_),
    .ZN(_24285_)
  );
  AND2_X1 _32412_ (
    .A1(_21466_),
    .A2(_22149_),
    .ZN(_24286_)
  );
  INV_X1 _32413_ (
    .A(_24286_),
    .ZN(_24287_)
  );
  AND2_X1 _32414_ (
    .A1(_00008_[0]),
    .A2(_24285_),
    .ZN(_24288_)
  );
  AND2_X1 _32415_ (
    .A1(_24287_),
    .A2(_24288_),
    .ZN(_24289_)
  );
  INV_X1 _32416_ (
    .A(_24289_),
    .ZN(_24290_)
  );
  AND2_X1 _32417_ (
    .A1(_21444_),
    .A2(_22149_),
    .ZN(_24291_)
  );
  INV_X1 _32418_ (
    .A(_24291_),
    .ZN(_24292_)
  );
  AND2_X1 _32419_ (
    .A1(_21655_),
    .A2(_00008_[2]),
    .ZN(_24293_)
  );
  INV_X1 _32420_ (
    .A(_24293_),
    .ZN(_24294_)
  );
  AND2_X1 _32421_ (
    .A1(_24292_),
    .A2(_24294_),
    .ZN(_24295_)
  );
  AND2_X1 _32422_ (
    .A1(_22147_),
    .A2(_24295_),
    .ZN(_24296_)
  );
  INV_X1 _32423_ (
    .A(_24296_),
    .ZN(_24297_)
  );
  AND2_X1 _32424_ (
    .A1(_24290_),
    .A2(_24297_),
    .ZN(_24298_)
  );
  AND2_X1 _32425_ (
    .A1(_22148_),
    .A2(_24298_),
    .ZN(_24299_)
  );
  INV_X1 _32426_ (
    .A(_24299_),
    .ZN(_24300_)
  );
  AND2_X1 _32427_ (
    .A1(_00008_[1]),
    .A2(_24283_),
    .ZN(_24301_)
  );
  INV_X1 _32428_ (
    .A(_24301_),
    .ZN(_24302_)
  );
  AND2_X1 _32429_ (
    .A1(_00008_[4]),
    .A2(_24300_),
    .ZN(_24303_)
  );
  AND2_X1 _32430_ (
    .A1(_24302_),
    .A2(_24303_),
    .ZN(_24304_)
  );
  INV_X1 _32431_ (
    .A(_24304_),
    .ZN(_24305_)
  );
  AND2_X1 _32432_ (
    .A1(_22150_),
    .A2(_24305_),
    .ZN(_24306_)
  );
  AND2_X1 _32433_ (
    .A1(_24268_),
    .A2(_24306_),
    .ZN(_24307_)
  );
  INV_X1 _32434_ (
    .A(_24307_),
    .ZN(_24308_)
  );
  AND2_X1 _32435_ (
    .A1(\cpuregs[29] [10]),
    .A2(_00008_[2]),
    .ZN(_24309_)
  );
  INV_X1 _32436_ (
    .A(_24309_),
    .ZN(_24310_)
  );
  AND2_X1 _32437_ (
    .A1(\cpuregs[25] [10]),
    .A2(_22149_),
    .ZN(_24311_)
  );
  INV_X1 _32438_ (
    .A(_24311_),
    .ZN(_24312_)
  );
  AND2_X1 _32439_ (
    .A1(_22148_),
    .A2(_24312_),
    .ZN(_24313_)
  );
  AND2_X1 _32440_ (
    .A1(_24310_),
    .A2(_24313_),
    .ZN(_24314_)
  );
  INV_X1 _32441_ (
    .A(_24314_),
    .ZN(_24315_)
  );
  AND2_X1 _32442_ (
    .A1(\cpuregs[27] [10]),
    .A2(_22149_),
    .ZN(_24316_)
  );
  INV_X1 _32443_ (
    .A(_24316_),
    .ZN(_24317_)
  );
  AND2_X1 _32444_ (
    .A1(\cpuregs[31] [10]),
    .A2(_00008_[2]),
    .ZN(_24318_)
  );
  INV_X1 _32445_ (
    .A(_24318_),
    .ZN(_24319_)
  );
  AND2_X1 _32446_ (
    .A1(_00008_[1]),
    .A2(_24319_),
    .ZN(_24320_)
  );
  AND2_X1 _32447_ (
    .A1(_24317_),
    .A2(_24320_),
    .ZN(_24321_)
  );
  INV_X1 _32448_ (
    .A(_24321_),
    .ZN(_24322_)
  );
  AND2_X1 _32449_ (
    .A1(_24315_),
    .A2(_24322_),
    .ZN(_24323_)
  );
  INV_X1 _32450_ (
    .A(_24323_),
    .ZN(_24324_)
  );
  AND2_X1 _32451_ (
    .A1(_00008_[0]),
    .A2(_24324_),
    .ZN(_24325_)
  );
  INV_X1 _32452_ (
    .A(_24325_),
    .ZN(_24326_)
  );
  AND2_X1 _32453_ (
    .A1(\cpuregs[24] [10]),
    .A2(_22149_),
    .ZN(_24327_)
  );
  INV_X1 _32454_ (
    .A(_24327_),
    .ZN(_24328_)
  );
  AND2_X1 _32455_ (
    .A1(\cpuregs[28] [10]),
    .A2(_00008_[2]),
    .ZN(_24329_)
  );
  INV_X1 _32456_ (
    .A(_24329_),
    .ZN(_24330_)
  );
  AND2_X1 _32457_ (
    .A1(_22148_),
    .A2(_24330_),
    .ZN(_24331_)
  );
  AND2_X1 _32458_ (
    .A1(_24328_),
    .A2(_24331_),
    .ZN(_24332_)
  );
  INV_X1 _32459_ (
    .A(_24332_),
    .ZN(_24333_)
  );
  AND2_X1 _32460_ (
    .A1(\cpuregs[26] [10]),
    .A2(_22149_),
    .ZN(_24334_)
  );
  INV_X1 _32461_ (
    .A(_24334_),
    .ZN(_24335_)
  );
  AND2_X1 _32462_ (
    .A1(\cpuregs[30] [10]),
    .A2(_00008_[2]),
    .ZN(_24336_)
  );
  INV_X1 _32463_ (
    .A(_24336_),
    .ZN(_24337_)
  );
  AND2_X1 _32464_ (
    .A1(_00008_[1]),
    .A2(_24337_),
    .ZN(_24338_)
  );
  AND2_X1 _32465_ (
    .A1(_24335_),
    .A2(_24338_),
    .ZN(_24339_)
  );
  INV_X1 _32466_ (
    .A(_24339_),
    .ZN(_24340_)
  );
  AND2_X1 _32467_ (
    .A1(_24333_),
    .A2(_24340_),
    .ZN(_24341_)
  );
  INV_X1 _32468_ (
    .A(_24341_),
    .ZN(_24342_)
  );
  AND2_X1 _32469_ (
    .A1(_22147_),
    .A2(_24342_),
    .ZN(_24343_)
  );
  INV_X1 _32470_ (
    .A(_24343_),
    .ZN(_24344_)
  );
  AND2_X1 _32471_ (
    .A1(_24326_),
    .A2(_24344_),
    .ZN(_24345_)
  );
  INV_X1 _32472_ (
    .A(_24345_),
    .ZN(_24346_)
  );
  AND2_X1 _32473_ (
    .A1(_00008_[4]),
    .A2(_24346_),
    .ZN(_24347_)
  );
  INV_X1 _32474_ (
    .A(_24347_),
    .ZN(_24348_)
  );
  AND2_X1 _32475_ (
    .A1(\cpuregs[9] [10]),
    .A2(_22148_),
    .ZN(_24349_)
  );
  INV_X1 _32476_ (
    .A(_24349_),
    .ZN(_24350_)
  );
  AND2_X1 _32477_ (
    .A1(\cpuregs[11] [10]),
    .A2(_00008_[1]),
    .ZN(_24351_)
  );
  INV_X1 _32478_ (
    .A(_24351_),
    .ZN(_24352_)
  );
  AND2_X1 _32479_ (
    .A1(_22149_),
    .A2(_24352_),
    .ZN(_24353_)
  );
  AND2_X1 _32480_ (
    .A1(_24350_),
    .A2(_24353_),
    .ZN(_24354_)
  );
  INV_X1 _32481_ (
    .A(_24354_),
    .ZN(_24355_)
  );
  AND2_X1 _32482_ (
    .A1(\cpuregs[13] [10]),
    .A2(_22148_),
    .ZN(_24356_)
  );
  INV_X1 _32483_ (
    .A(_24356_),
    .ZN(_24357_)
  );
  AND2_X1 _32484_ (
    .A1(\cpuregs[15] [10]),
    .A2(_00008_[1]),
    .ZN(_24358_)
  );
  INV_X1 _32485_ (
    .A(_24358_),
    .ZN(_24359_)
  );
  AND2_X1 _32486_ (
    .A1(_00008_[2]),
    .A2(_24359_),
    .ZN(_24360_)
  );
  AND2_X1 _32487_ (
    .A1(_24357_),
    .A2(_24360_),
    .ZN(_24361_)
  );
  INV_X1 _32488_ (
    .A(_24361_),
    .ZN(_24362_)
  );
  AND2_X1 _32489_ (
    .A1(_24355_),
    .A2(_24362_),
    .ZN(_24363_)
  );
  INV_X1 _32490_ (
    .A(_24363_),
    .ZN(_24364_)
  );
  AND2_X1 _32491_ (
    .A1(_00008_[0]),
    .A2(_24364_),
    .ZN(_24365_)
  );
  INV_X1 _32492_ (
    .A(_24365_),
    .ZN(_24366_)
  );
  AND2_X1 _32493_ (
    .A1(\cpuregs[8] [10]),
    .A2(_22148_),
    .ZN(_24367_)
  );
  INV_X1 _32494_ (
    .A(_24367_),
    .ZN(_24368_)
  );
  AND2_X1 _32495_ (
    .A1(\cpuregs[10] [10]),
    .A2(_00008_[1]),
    .ZN(_24369_)
  );
  INV_X1 _32496_ (
    .A(_24369_),
    .ZN(_24370_)
  );
  AND2_X1 _32497_ (
    .A1(_22149_),
    .A2(_24370_),
    .ZN(_24371_)
  );
  AND2_X1 _32498_ (
    .A1(_24368_),
    .A2(_24371_),
    .ZN(_24372_)
  );
  INV_X1 _32499_ (
    .A(_24372_),
    .ZN(_24373_)
  );
  AND2_X1 _32500_ (
    .A1(\cpuregs[12] [10]),
    .A2(_22148_),
    .ZN(_24374_)
  );
  INV_X1 _32501_ (
    .A(_24374_),
    .ZN(_24375_)
  );
  AND2_X1 _32502_ (
    .A1(\cpuregs[14] [10]),
    .A2(_00008_[1]),
    .ZN(_24376_)
  );
  INV_X1 _32503_ (
    .A(_24376_),
    .ZN(_24377_)
  );
  AND2_X1 _32504_ (
    .A1(_00008_[2]),
    .A2(_24377_),
    .ZN(_24378_)
  );
  AND2_X1 _32505_ (
    .A1(_24375_),
    .A2(_24378_),
    .ZN(_24379_)
  );
  INV_X1 _32506_ (
    .A(_24379_),
    .ZN(_24380_)
  );
  AND2_X1 _32507_ (
    .A1(_24373_),
    .A2(_24380_),
    .ZN(_24381_)
  );
  INV_X1 _32508_ (
    .A(_24381_),
    .ZN(_24382_)
  );
  AND2_X1 _32509_ (
    .A1(_22147_),
    .A2(_24382_),
    .ZN(_24383_)
  );
  INV_X1 _32510_ (
    .A(_24383_),
    .ZN(_24384_)
  );
  AND2_X1 _32511_ (
    .A1(_24366_),
    .A2(_24384_),
    .ZN(_24385_)
  );
  INV_X1 _32512_ (
    .A(_24385_),
    .ZN(_24386_)
  );
  AND2_X1 _32513_ (
    .A1(_22151_),
    .A2(_24386_),
    .ZN(_24387_)
  );
  INV_X1 _32514_ (
    .A(_24387_),
    .ZN(_24388_)
  );
  AND2_X1 _32515_ (
    .A1(_24348_),
    .A2(_24388_),
    .ZN(_24389_)
  );
  INV_X1 _32516_ (
    .A(_24389_),
    .ZN(_24390_)
  );
  AND2_X1 _32517_ (
    .A1(_00008_[3]),
    .A2(_24390_),
    .ZN(_24391_)
  );
  INV_X1 _32518_ (
    .A(_24391_),
    .ZN(_24392_)
  );
  AND2_X1 _32519_ (
    .A1(_22546_),
    .A2(_24308_),
    .ZN(_24393_)
  );
  AND2_X1 _32520_ (
    .A1(_24392_),
    .A2(_24393_),
    .ZN(_24394_)
  );
  INV_X1 _32521_ (
    .A(_24394_),
    .ZN(_24395_)
  );
  AND2_X1 _32522_ (
    .A1(_24228_),
    .A2(_24395_),
    .ZN(_24396_)
  );
  INV_X1 _32523_ (
    .A(_24396_),
    .ZN(_24397_)
  );
  AND2_X1 _32524_ (
    .A1(_22271_),
    .A2(_24397_),
    .ZN(_24398_)
  );
  INV_X1 _32525_ (
    .A(_24398_),
    .ZN(_24399_)
  );
  AND2_X1 _32526_ (
    .A1(reg_op1[9]),
    .A2(_22285_),
    .ZN(_24400_)
  );
  INV_X1 _32527_ (
    .A(_24400_),
    .ZN(_24401_)
  );
  AND2_X1 _32528_ (
    .A1(_23796_),
    .A2(_24401_),
    .ZN(_24402_)
  );
  AND2_X1 _32529_ (
    .A1(reg_op1[14]),
    .A2(_22290_),
    .ZN(_24403_)
  );
  INV_X1 _32530_ (
    .A(_24403_),
    .ZN(_24404_)
  );
  AND2_X1 _32531_ (
    .A1(_23793_),
    .A2(_24404_),
    .ZN(_24405_)
  );
  AND2_X1 _32532_ (
    .A1(_22572_),
    .A2(_24402_),
    .ZN(_24406_)
  );
  INV_X1 _32533_ (
    .A(_24406_),
    .ZN(_24407_)
  );
  AND2_X1 _32534_ (
    .A1(_22573_),
    .A2(_24405_),
    .ZN(_24408_)
  );
  INV_X1 _32535_ (
    .A(_24408_),
    .ZN(_24409_)
  );
  AND2_X1 _32536_ (
    .A1(_22295_),
    .A2(_24409_),
    .ZN(_24410_)
  );
  AND2_X1 _32537_ (
    .A1(_24407_),
    .A2(_24410_),
    .ZN(_24411_)
  );
  INV_X1 _32538_ (
    .A(_24411_),
    .ZN(_24412_)
  );
  AND2_X1 _32539_ (
    .A1(_22333_),
    .A2(_24399_),
    .ZN(_24413_)
  );
  AND2_X1 _32540_ (
    .A1(_24412_),
    .A2(_24413_),
    .ZN(_24414_)
  );
  AND2_X1 _32541_ (
    .A1(reg_op1[10]),
    .A2(decoded_imm[10]),
    .ZN(_24415_)
  );
  INV_X1 _32542_ (
    .A(_24415_),
    .ZN(_24416_)
  );
  AND2_X1 _32543_ (
    .A1(_21177_),
    .A2(_21999_),
    .ZN(_24417_)
  );
  INV_X1 _32544_ (
    .A(_24417_),
    .ZN(_24418_)
  );
  AND2_X1 _32545_ (
    .A1(_24416_),
    .A2(_24418_),
    .ZN(_24419_)
  );
  INV_X1 _32546_ (
    .A(_24419_),
    .ZN(_24420_)
  );
  AND2_X1 _32547_ (
    .A1(_24024_),
    .A2(_24209_),
    .ZN(_24421_)
  );
  AND2_X1 _32548_ (
    .A1(_24207_),
    .A2(_24421_),
    .ZN(_24422_)
  );
  INV_X1 _32549_ (
    .A(_24422_),
    .ZN(_24423_)
  );
  AND2_X1 _32550_ (
    .A1(_24419_),
    .A2(_24423_),
    .ZN(_24424_)
  );
  INV_X1 _32551_ (
    .A(_24424_),
    .ZN(_24425_)
  );
  AND2_X1 _32552_ (
    .A1(_24420_),
    .A2(_24422_),
    .ZN(_24426_)
  );
  INV_X1 _32553_ (
    .A(_24426_),
    .ZN(_24427_)
  );
  AND2_X1 _32554_ (
    .A1(_22559_),
    .A2(_24427_),
    .ZN(_24428_)
  );
  AND2_X1 _32555_ (
    .A1(_24425_),
    .A2(_24428_),
    .ZN(_24429_)
  );
  INV_X1 _32556_ (
    .A(_24429_),
    .ZN(_24430_)
  );
  AND2_X1 _32557_ (
    .A1(_24414_),
    .A2(_24430_),
    .ZN(_24431_)
  );
  INV_X1 _32558_ (
    .A(_24431_),
    .ZN(_24432_)
  );
  AND2_X1 _32559_ (
    .A1(_24226_),
    .A2(_24432_),
    .ZN(_00067_)
  );
  AND2_X1 _32560_ (
    .A1(_21178_),
    .A2(_22334_),
    .ZN(_24433_)
  );
  INV_X1 _32561_ (
    .A(_24433_),
    .ZN(_24434_)
  );
  AND2_X1 _32562_ (
    .A1(reg_op1[11]),
    .A2(decoded_imm[11]),
    .ZN(_24435_)
  );
  INV_X1 _32563_ (
    .A(_24435_),
    .ZN(_24436_)
  );
  AND2_X1 _32564_ (
    .A1(_21178_),
    .A2(_21998_),
    .ZN(_24437_)
  );
  INV_X1 _32565_ (
    .A(_24437_),
    .ZN(_24438_)
  );
  AND2_X1 _32566_ (
    .A1(_24436_),
    .A2(_24438_),
    .ZN(_24439_)
  );
  INV_X1 _32567_ (
    .A(_24439_),
    .ZN(_24440_)
  );
  AND2_X1 _32568_ (
    .A1(_24416_),
    .A2(_24440_),
    .ZN(_24441_)
  );
  AND2_X1 _32569_ (
    .A1(_24425_),
    .A2(_24441_),
    .ZN(_24442_)
  );
  INV_X1 _32570_ (
    .A(_24442_),
    .ZN(_24443_)
  );
  AND2_X1 _32571_ (
    .A1(_24424_),
    .A2(_24439_),
    .ZN(_24444_)
  );
  INV_X1 _32572_ (
    .A(_24444_),
    .ZN(_24445_)
  );
  AND2_X1 _32573_ (
    .A1(_24415_),
    .A2(_24439_),
    .ZN(_24446_)
  );
  INV_X1 _32574_ (
    .A(_24446_),
    .ZN(_24447_)
  );
  AND2_X1 _32575_ (
    .A1(_22559_),
    .A2(_24447_),
    .ZN(_24448_)
  );
  AND2_X1 _32576_ (
    .A1(_24445_),
    .A2(_24448_),
    .ZN(_24449_)
  );
  AND2_X1 _32577_ (
    .A1(_24443_),
    .A2(_24449_),
    .ZN(_24450_)
  );
  INV_X1 _32578_ (
    .A(_24450_),
    .ZN(_24451_)
  );
  AND2_X1 _32579_ (
    .A1(reg_pc[11]),
    .A2(_22335_),
    .ZN(_24452_)
  );
  INV_X1 _32580_ (
    .A(_24452_),
    .ZN(_24453_)
  );
  AND2_X1 _32581_ (
    .A1(\cpuregs[20] [11]),
    .A2(_00008_[2]),
    .ZN(_24454_)
  );
  INV_X1 _32582_ (
    .A(_24454_),
    .ZN(_24455_)
  );
  AND2_X1 _32583_ (
    .A1(\cpuregs[16] [11]),
    .A2(_22149_),
    .ZN(_24456_)
  );
  INV_X1 _32584_ (
    .A(_24456_),
    .ZN(_24457_)
  );
  AND2_X1 _32585_ (
    .A1(_24455_),
    .A2(_24457_),
    .ZN(_24458_)
  );
  INV_X1 _32586_ (
    .A(_24458_),
    .ZN(_24459_)
  );
  AND2_X1 _32587_ (
    .A1(_22147_),
    .A2(_24459_),
    .ZN(_24460_)
  );
  INV_X1 _32588_ (
    .A(_24460_),
    .ZN(_24461_)
  );
  AND2_X1 _32589_ (
    .A1(\cpuregs[21] [11]),
    .A2(_00008_[2]),
    .ZN(_24462_)
  );
  INV_X1 _32590_ (
    .A(_24462_),
    .ZN(_24463_)
  );
  AND2_X1 _32591_ (
    .A1(\cpuregs[17] [11]),
    .A2(_22149_),
    .ZN(_24464_)
  );
  INV_X1 _32592_ (
    .A(_24464_),
    .ZN(_24465_)
  );
  AND2_X1 _32593_ (
    .A1(_24463_),
    .A2(_24465_),
    .ZN(_24466_)
  );
  INV_X1 _32594_ (
    .A(_24466_),
    .ZN(_24467_)
  );
  AND2_X1 _32595_ (
    .A1(_00008_[0]),
    .A2(_24467_),
    .ZN(_24468_)
  );
  INV_X1 _32596_ (
    .A(_24468_),
    .ZN(_24469_)
  );
  AND2_X1 _32597_ (
    .A1(_24461_),
    .A2(_24469_),
    .ZN(_24470_)
  );
  AND2_X1 _32598_ (
    .A1(_22148_),
    .A2(_24470_),
    .ZN(_24471_)
  );
  INV_X1 _32599_ (
    .A(_24471_),
    .ZN(_24472_)
  );
  AND2_X1 _32600_ (
    .A1(\cpuregs[22] [11]),
    .A2(_00008_[2]),
    .ZN(_24473_)
  );
  INV_X1 _32601_ (
    .A(_24473_),
    .ZN(_24474_)
  );
  AND2_X1 _32602_ (
    .A1(\cpuregs[18] [11]),
    .A2(_22149_),
    .ZN(_24475_)
  );
  INV_X1 _32603_ (
    .A(_24475_),
    .ZN(_24476_)
  );
  AND2_X1 _32604_ (
    .A1(_24474_),
    .A2(_24476_),
    .ZN(_24477_)
  );
  INV_X1 _32605_ (
    .A(_24477_),
    .ZN(_24478_)
  );
  AND2_X1 _32606_ (
    .A1(_22147_),
    .A2(_24478_),
    .ZN(_24479_)
  );
  INV_X1 _32607_ (
    .A(_24479_),
    .ZN(_24480_)
  );
  AND2_X1 _32608_ (
    .A1(\cpuregs[23] [11]),
    .A2(_00008_[2]),
    .ZN(_24481_)
  );
  INV_X1 _32609_ (
    .A(_24481_),
    .ZN(_24482_)
  );
  AND2_X1 _32610_ (
    .A1(\cpuregs[19] [11]),
    .A2(_22149_),
    .ZN(_24483_)
  );
  INV_X1 _32611_ (
    .A(_24483_),
    .ZN(_24484_)
  );
  AND2_X1 _32612_ (
    .A1(_24482_),
    .A2(_24484_),
    .ZN(_24485_)
  );
  INV_X1 _32613_ (
    .A(_24485_),
    .ZN(_24486_)
  );
  AND2_X1 _32614_ (
    .A1(_00008_[0]),
    .A2(_24486_),
    .ZN(_24487_)
  );
  INV_X1 _32615_ (
    .A(_24487_),
    .ZN(_24488_)
  );
  AND2_X1 _32616_ (
    .A1(_24480_),
    .A2(_24488_),
    .ZN(_24489_)
  );
  AND2_X1 _32617_ (
    .A1(_00008_[1]),
    .A2(_24489_),
    .ZN(_24490_)
  );
  INV_X1 _32618_ (
    .A(_24490_),
    .ZN(_24491_)
  );
  AND2_X1 _32619_ (
    .A1(_24472_),
    .A2(_24491_),
    .ZN(_24492_)
  );
  AND2_X1 _32620_ (
    .A1(\cpuregs[27] [11]),
    .A2(_00008_[0]),
    .ZN(_24493_)
  );
  INV_X1 _32621_ (
    .A(_24493_),
    .ZN(_24494_)
  );
  AND2_X1 _32622_ (
    .A1(\cpuregs[26] [11]),
    .A2(_22147_),
    .ZN(_24495_)
  );
  INV_X1 _32623_ (
    .A(_24495_),
    .ZN(_24496_)
  );
  AND2_X1 _32624_ (
    .A1(_22149_),
    .A2(_24496_),
    .ZN(_24497_)
  );
  AND2_X1 _32625_ (
    .A1(_24494_),
    .A2(_24497_),
    .ZN(_24498_)
  );
  INV_X1 _32626_ (
    .A(_24498_),
    .ZN(_24499_)
  );
  AND2_X1 _32627_ (
    .A1(\cpuregs[31] [11]),
    .A2(_00008_[0]),
    .ZN(_24500_)
  );
  INV_X1 _32628_ (
    .A(_24500_),
    .ZN(_24501_)
  );
  AND2_X1 _32629_ (
    .A1(\cpuregs[30] [11]),
    .A2(_22147_),
    .ZN(_24502_)
  );
  INV_X1 _32630_ (
    .A(_24502_),
    .ZN(_24503_)
  );
  AND2_X1 _32631_ (
    .A1(_00008_[2]),
    .A2(_24503_),
    .ZN(_24504_)
  );
  AND2_X1 _32632_ (
    .A1(_24501_),
    .A2(_24504_),
    .ZN(_24505_)
  );
  INV_X1 _32633_ (
    .A(_24505_),
    .ZN(_24506_)
  );
  AND2_X1 _32634_ (
    .A1(_24499_),
    .A2(_24506_),
    .ZN(_24507_)
  );
  INV_X1 _32635_ (
    .A(_24507_),
    .ZN(_24508_)
  );
  AND2_X1 _32636_ (
    .A1(_00008_[1]),
    .A2(_24508_),
    .ZN(_24509_)
  );
  INV_X1 _32637_ (
    .A(_24509_),
    .ZN(_24510_)
  );
  AND2_X1 _32638_ (
    .A1(\cpuregs[25] [11]),
    .A2(_00008_[0]),
    .ZN(_24511_)
  );
  INV_X1 _32639_ (
    .A(_24511_),
    .ZN(_24512_)
  );
  AND2_X1 _32640_ (
    .A1(\cpuregs[24] [11]),
    .A2(_22147_),
    .ZN(_24513_)
  );
  INV_X1 _32641_ (
    .A(_24513_),
    .ZN(_24514_)
  );
  AND2_X1 _32642_ (
    .A1(_22149_),
    .A2(_24514_),
    .ZN(_24515_)
  );
  AND2_X1 _32643_ (
    .A1(_24512_),
    .A2(_24515_),
    .ZN(_24516_)
  );
  INV_X1 _32644_ (
    .A(_24516_),
    .ZN(_24517_)
  );
  AND2_X1 _32645_ (
    .A1(\cpuregs[29] [11]),
    .A2(_00008_[0]),
    .ZN(_24518_)
  );
  INV_X1 _32646_ (
    .A(_24518_),
    .ZN(_24519_)
  );
  AND2_X1 _32647_ (
    .A1(\cpuregs[28] [11]),
    .A2(_22147_),
    .ZN(_24520_)
  );
  INV_X1 _32648_ (
    .A(_24520_),
    .ZN(_24521_)
  );
  AND2_X1 _32649_ (
    .A1(_00008_[2]),
    .A2(_24521_),
    .ZN(_24522_)
  );
  AND2_X1 _32650_ (
    .A1(_24519_),
    .A2(_24522_),
    .ZN(_24523_)
  );
  INV_X1 _32651_ (
    .A(_24523_),
    .ZN(_24524_)
  );
  AND2_X1 _32652_ (
    .A1(_24517_),
    .A2(_24524_),
    .ZN(_24525_)
  );
  INV_X1 _32653_ (
    .A(_24525_),
    .ZN(_24526_)
  );
  AND2_X1 _32654_ (
    .A1(_22148_),
    .A2(_24526_),
    .ZN(_24527_)
  );
  INV_X1 _32655_ (
    .A(_24527_),
    .ZN(_24528_)
  );
  AND2_X1 _32656_ (
    .A1(_00008_[3]),
    .A2(_24510_),
    .ZN(_24529_)
  );
  AND2_X1 _32657_ (
    .A1(_24528_),
    .A2(_24529_),
    .ZN(_24530_)
  );
  INV_X1 _32658_ (
    .A(_24530_),
    .ZN(_24531_)
  );
  AND2_X1 _32659_ (
    .A1(_22150_),
    .A2(_24492_),
    .ZN(_24532_)
  );
  INV_X1 _32660_ (
    .A(_24532_),
    .ZN(_24533_)
  );
  AND2_X1 _32661_ (
    .A1(_00008_[4]),
    .A2(_24533_),
    .ZN(_24534_)
  );
  AND2_X1 _32662_ (
    .A1(_24531_),
    .A2(_24534_),
    .ZN(_24535_)
  );
  INV_X1 _32663_ (
    .A(_24535_),
    .ZN(_24536_)
  );
  AND2_X1 _32664_ (
    .A1(\cpuregs[10] [11]),
    .A2(_22149_),
    .ZN(_24537_)
  );
  INV_X1 _32665_ (
    .A(_24537_),
    .ZN(_24538_)
  );
  AND2_X1 _32666_ (
    .A1(\cpuregs[14] [11]),
    .A2(_00008_[2]),
    .ZN(_24539_)
  );
  INV_X1 _32667_ (
    .A(_24539_),
    .ZN(_24540_)
  );
  AND2_X1 _32668_ (
    .A1(_22147_),
    .A2(_24540_),
    .ZN(_24541_)
  );
  AND2_X1 _32669_ (
    .A1(_24538_),
    .A2(_24541_),
    .ZN(_24542_)
  );
  INV_X1 _32670_ (
    .A(_24542_),
    .ZN(_24543_)
  );
  AND2_X1 _32671_ (
    .A1(\cpuregs[15] [11]),
    .A2(_00008_[2]),
    .ZN(_24544_)
  );
  INV_X1 _32672_ (
    .A(_24544_),
    .ZN(_24545_)
  );
  AND2_X1 _32673_ (
    .A1(\cpuregs[11] [11]),
    .A2(_22149_),
    .ZN(_24546_)
  );
  INV_X1 _32674_ (
    .A(_24546_),
    .ZN(_24547_)
  );
  AND2_X1 _32675_ (
    .A1(_00008_[0]),
    .A2(_24547_),
    .ZN(_24548_)
  );
  AND2_X1 _32676_ (
    .A1(_24545_),
    .A2(_24548_),
    .ZN(_24549_)
  );
  INV_X1 _32677_ (
    .A(_24549_),
    .ZN(_24550_)
  );
  AND2_X1 _32678_ (
    .A1(_24543_),
    .A2(_24550_),
    .ZN(_24551_)
  );
  INV_X1 _32679_ (
    .A(_24551_),
    .ZN(_24552_)
  );
  AND2_X1 _32680_ (
    .A1(_00008_[3]),
    .A2(_24552_),
    .ZN(_24553_)
  );
  INV_X1 _32681_ (
    .A(_24553_),
    .ZN(_24554_)
  );
  AND2_X1 _32682_ (
    .A1(\cpuregs[2] [11]),
    .A2(_22149_),
    .ZN(_24555_)
  );
  INV_X1 _32683_ (
    .A(_24555_),
    .ZN(_24556_)
  );
  AND2_X1 _32684_ (
    .A1(\cpuregs[6] [11]),
    .A2(_00008_[2]),
    .ZN(_24557_)
  );
  INV_X1 _32685_ (
    .A(_24557_),
    .ZN(_24558_)
  );
  AND2_X1 _32686_ (
    .A1(_22147_),
    .A2(_24558_),
    .ZN(_24559_)
  );
  AND2_X1 _32687_ (
    .A1(_24556_),
    .A2(_24559_),
    .ZN(_24560_)
  );
  INV_X1 _32688_ (
    .A(_24560_),
    .ZN(_24561_)
  );
  AND2_X1 _32689_ (
    .A1(\cpuregs[3] [11]),
    .A2(_22149_),
    .ZN(_24562_)
  );
  INV_X1 _32690_ (
    .A(_24562_),
    .ZN(_24563_)
  );
  AND2_X1 _32691_ (
    .A1(\cpuregs[7] [11]),
    .A2(_00008_[2]),
    .ZN(_24564_)
  );
  INV_X1 _32692_ (
    .A(_24564_),
    .ZN(_24565_)
  );
  AND2_X1 _32693_ (
    .A1(_00008_[0]),
    .A2(_24565_),
    .ZN(_24566_)
  );
  AND2_X1 _32694_ (
    .A1(_24563_),
    .A2(_24566_),
    .ZN(_24567_)
  );
  INV_X1 _32695_ (
    .A(_24567_),
    .ZN(_24568_)
  );
  AND2_X1 _32696_ (
    .A1(_24561_),
    .A2(_24568_),
    .ZN(_24569_)
  );
  INV_X1 _32697_ (
    .A(_24569_),
    .ZN(_24570_)
  );
  AND2_X1 _32698_ (
    .A1(_22150_),
    .A2(_24570_),
    .ZN(_24571_)
  );
  INV_X1 _32699_ (
    .A(_24571_),
    .ZN(_24572_)
  );
  AND2_X1 _32700_ (
    .A1(\cpuregs[8] [11]),
    .A2(_22149_),
    .ZN(_24573_)
  );
  INV_X1 _32701_ (
    .A(_24573_),
    .ZN(_24574_)
  );
  AND2_X1 _32702_ (
    .A1(\cpuregs[12] [11]),
    .A2(_00008_[2]),
    .ZN(_24575_)
  );
  INV_X1 _32703_ (
    .A(_24575_),
    .ZN(_24576_)
  );
  AND2_X1 _32704_ (
    .A1(_22147_),
    .A2(_24576_),
    .ZN(_24577_)
  );
  AND2_X1 _32705_ (
    .A1(_24574_),
    .A2(_24577_),
    .ZN(_24578_)
  );
  INV_X1 _32706_ (
    .A(_24578_),
    .ZN(_24579_)
  );
  AND2_X1 _32707_ (
    .A1(\cpuregs[13] [11]),
    .A2(_00008_[2]),
    .ZN(_24580_)
  );
  INV_X1 _32708_ (
    .A(_24580_),
    .ZN(_24581_)
  );
  AND2_X1 _32709_ (
    .A1(\cpuregs[9] [11]),
    .A2(_22149_),
    .ZN(_24582_)
  );
  INV_X1 _32710_ (
    .A(_24582_),
    .ZN(_24583_)
  );
  AND2_X1 _32711_ (
    .A1(_00008_[0]),
    .A2(_24583_),
    .ZN(_24584_)
  );
  AND2_X1 _32712_ (
    .A1(_24581_),
    .A2(_24584_),
    .ZN(_24585_)
  );
  INV_X1 _32713_ (
    .A(_24585_),
    .ZN(_24586_)
  );
  AND2_X1 _32714_ (
    .A1(_24579_),
    .A2(_24586_),
    .ZN(_24587_)
  );
  AND2_X1 _32715_ (
    .A1(\cpuregs[0] [11]),
    .A2(_22149_),
    .ZN(_24588_)
  );
  INV_X1 _32716_ (
    .A(_24588_),
    .ZN(_24589_)
  );
  AND2_X1 _32717_ (
    .A1(\cpuregs[4] [11]),
    .A2(_00008_[2]),
    .ZN(_24590_)
  );
  INV_X1 _32718_ (
    .A(_24590_),
    .ZN(_24591_)
  );
  AND2_X1 _32719_ (
    .A1(_22147_),
    .A2(_24591_),
    .ZN(_24592_)
  );
  AND2_X1 _32720_ (
    .A1(_24589_),
    .A2(_24592_),
    .ZN(_24593_)
  );
  INV_X1 _32721_ (
    .A(_24593_),
    .ZN(_24594_)
  );
  AND2_X1 _32722_ (
    .A1(\cpuregs[1] [11]),
    .A2(_22149_),
    .ZN(_24595_)
  );
  INV_X1 _32723_ (
    .A(_24595_),
    .ZN(_24596_)
  );
  AND2_X1 _32724_ (
    .A1(\cpuregs[5] [11]),
    .A2(_00008_[2]),
    .ZN(_24597_)
  );
  INV_X1 _32725_ (
    .A(_24597_),
    .ZN(_24598_)
  );
  AND2_X1 _32726_ (
    .A1(_00008_[0]),
    .A2(_24598_),
    .ZN(_24599_)
  );
  AND2_X1 _32727_ (
    .A1(_24596_),
    .A2(_24599_),
    .ZN(_24600_)
  );
  INV_X1 _32728_ (
    .A(_24600_),
    .ZN(_24601_)
  );
  AND2_X1 _32729_ (
    .A1(_00008_[3]),
    .A2(_24587_),
    .ZN(_24602_)
  );
  INV_X1 _32730_ (
    .A(_24602_),
    .ZN(_24603_)
  );
  AND2_X1 _32731_ (
    .A1(_22150_),
    .A2(_24601_),
    .ZN(_24604_)
  );
  AND2_X1 _32732_ (
    .A1(_24594_),
    .A2(_24604_),
    .ZN(_24605_)
  );
  INV_X1 _32733_ (
    .A(_24605_),
    .ZN(_24606_)
  );
  AND2_X1 _32734_ (
    .A1(_24603_),
    .A2(_24606_),
    .ZN(_24607_)
  );
  INV_X1 _32735_ (
    .A(_24607_),
    .ZN(_24608_)
  );
  AND2_X1 _32736_ (
    .A1(_22148_),
    .A2(_24608_),
    .ZN(_24609_)
  );
  INV_X1 _32737_ (
    .A(_24609_),
    .ZN(_24610_)
  );
  AND2_X1 _32738_ (
    .A1(_00008_[1]),
    .A2(_24572_),
    .ZN(_24611_)
  );
  AND2_X1 _32739_ (
    .A1(_24554_),
    .A2(_24611_),
    .ZN(_24612_)
  );
  INV_X1 _32740_ (
    .A(_24612_),
    .ZN(_24613_)
  );
  AND2_X1 _32741_ (
    .A1(_22151_),
    .A2(_24613_),
    .ZN(_24614_)
  );
  AND2_X1 _32742_ (
    .A1(_24610_),
    .A2(_24614_),
    .ZN(_24615_)
  );
  INV_X1 _32743_ (
    .A(_24615_),
    .ZN(_24616_)
  );
  AND2_X1 _32744_ (
    .A1(_22546_),
    .A2(_24536_),
    .ZN(_24617_)
  );
  AND2_X1 _32745_ (
    .A1(_24616_),
    .A2(_24617_),
    .ZN(_24618_)
  );
  INV_X1 _32746_ (
    .A(_24618_),
    .ZN(_24619_)
  );
  AND2_X1 _32747_ (
    .A1(_24453_),
    .A2(_24619_),
    .ZN(_24620_)
  );
  INV_X1 _32748_ (
    .A(_24620_),
    .ZN(_24621_)
  );
  AND2_X1 _32749_ (
    .A1(_22271_),
    .A2(_24621_),
    .ZN(_24622_)
  );
  INV_X1 _32750_ (
    .A(_24622_),
    .ZN(_24623_)
  );
  AND2_X1 _32751_ (
    .A1(reg_op1[10]),
    .A2(_22285_),
    .ZN(_24624_)
  );
  INV_X1 _32752_ (
    .A(_24624_),
    .ZN(_24625_)
  );
  AND2_X1 _32753_ (
    .A1(_24005_),
    .A2(_24625_),
    .ZN(_24626_)
  );
  AND2_X1 _32754_ (
    .A1(reg_op1[15]),
    .A2(_22290_),
    .ZN(_24627_)
  );
  INV_X1 _32755_ (
    .A(_24627_),
    .ZN(_24628_)
  );
  AND2_X1 _32756_ (
    .A1(_24002_),
    .A2(_24628_),
    .ZN(_24629_)
  );
  AND2_X1 _32757_ (
    .A1(_22573_),
    .A2(_24629_),
    .ZN(_24630_)
  );
  INV_X1 _32758_ (
    .A(_24630_),
    .ZN(_24631_)
  );
  AND2_X1 _32759_ (
    .A1(_22572_),
    .A2(_24626_),
    .ZN(_24632_)
  );
  INV_X1 _32760_ (
    .A(_24632_),
    .ZN(_24633_)
  );
  AND2_X1 _32761_ (
    .A1(_22295_),
    .A2(_24631_),
    .ZN(_24634_)
  );
  AND2_X1 _32762_ (
    .A1(_24633_),
    .A2(_24634_),
    .ZN(_24635_)
  );
  INV_X1 _32763_ (
    .A(_24635_),
    .ZN(_24636_)
  );
  AND2_X1 _32764_ (
    .A1(_24623_),
    .A2(_24636_),
    .ZN(_24637_)
  );
  AND2_X1 _32765_ (
    .A1(_24451_),
    .A2(_24637_),
    .ZN(_24638_)
  );
  AND2_X1 _32766_ (
    .A1(_22333_),
    .A2(_24638_),
    .ZN(_24639_)
  );
  INV_X1 _32767_ (
    .A(_24639_),
    .ZN(_24640_)
  );
  AND2_X1 _32768_ (
    .A1(_24434_),
    .A2(_24640_),
    .ZN(_00068_)
  );
  AND2_X1 _32769_ (
    .A1(_21179_),
    .A2(_22334_),
    .ZN(_24641_)
  );
  INV_X1 _32770_ (
    .A(_24641_),
    .ZN(_24642_)
  );
  AND2_X1 _32771_ (
    .A1(reg_pc[12]),
    .A2(_22335_),
    .ZN(_24643_)
  );
  INV_X1 _32772_ (
    .A(_24643_),
    .ZN(_24644_)
  );
  AND2_X1 _32773_ (
    .A1(_21599_),
    .A2(_22149_),
    .ZN(_24645_)
  );
  INV_X1 _32774_ (
    .A(_24645_),
    .ZN(_24646_)
  );
  AND2_X1 _32775_ (
    .A1(_21419_),
    .A2(_00008_[2]),
    .ZN(_24647_)
  );
  INV_X1 _32776_ (
    .A(_24647_),
    .ZN(_24648_)
  );
  AND2_X1 _32777_ (
    .A1(_24646_),
    .A2(_24648_),
    .ZN(_24649_)
  );
  AND2_X1 _32778_ (
    .A1(_22147_),
    .A2(_24649_),
    .ZN(_24650_)
  );
  INV_X1 _32779_ (
    .A(_24650_),
    .ZN(_24651_)
  );
  AND2_X1 _32780_ (
    .A1(_21379_),
    .A2(_00008_[2]),
    .ZN(_24652_)
  );
  INV_X1 _32781_ (
    .A(_24652_),
    .ZN(_24653_)
  );
  AND2_X1 _32782_ (
    .A1(_21625_),
    .A2(_22149_),
    .ZN(_24654_)
  );
  INV_X1 _32783_ (
    .A(_24654_),
    .ZN(_24655_)
  );
  AND2_X1 _32784_ (
    .A1(_00008_[0]),
    .A2(_24655_),
    .ZN(_24656_)
  );
  AND2_X1 _32785_ (
    .A1(_24653_),
    .A2(_24656_),
    .ZN(_24657_)
  );
  INV_X1 _32786_ (
    .A(_24657_),
    .ZN(_24658_)
  );
  AND2_X1 _32787_ (
    .A1(_24651_),
    .A2(_24658_),
    .ZN(_24659_)
  );
  AND2_X1 _32788_ (
    .A1(_00008_[1]),
    .A2(_24659_),
    .ZN(_24660_)
  );
  INV_X1 _32789_ (
    .A(_24660_),
    .ZN(_24661_)
  );
  AND2_X1 _32790_ (
    .A1(_21445_),
    .A2(_22149_),
    .ZN(_24662_)
  );
  INV_X1 _32791_ (
    .A(_24662_),
    .ZN(_24663_)
  );
  AND2_X1 _32792_ (
    .A1(_21656_),
    .A2(_00008_[2]),
    .ZN(_24664_)
  );
  INV_X1 _32793_ (
    .A(_24664_),
    .ZN(_24665_)
  );
  AND2_X1 _32794_ (
    .A1(_24663_),
    .A2(_24665_),
    .ZN(_24666_)
  );
  AND2_X1 _32795_ (
    .A1(_22147_),
    .A2(_24666_),
    .ZN(_24667_)
  );
  INV_X1 _32796_ (
    .A(_24667_),
    .ZN(_24668_)
  );
  AND2_X1 _32797_ (
    .A1(_21766_),
    .A2(_00008_[2]),
    .ZN(_24669_)
  );
  INV_X1 _32798_ (
    .A(_24669_),
    .ZN(_24670_)
  );
  AND2_X1 _32799_ (
    .A1(_21467_),
    .A2(_22149_),
    .ZN(_24671_)
  );
  INV_X1 _32800_ (
    .A(_24671_),
    .ZN(_24672_)
  );
  AND2_X1 _32801_ (
    .A1(_00008_[0]),
    .A2(_24670_),
    .ZN(_24673_)
  );
  AND2_X1 _32802_ (
    .A1(_24672_),
    .A2(_24673_),
    .ZN(_24674_)
  );
  INV_X1 _32803_ (
    .A(_24674_),
    .ZN(_24675_)
  );
  AND2_X1 _32804_ (
    .A1(_24668_),
    .A2(_24675_),
    .ZN(_24676_)
  );
  AND2_X1 _32805_ (
    .A1(_22148_),
    .A2(_24676_),
    .ZN(_24677_)
  );
  INV_X1 _32806_ (
    .A(_24677_),
    .ZN(_24678_)
  );
  AND2_X1 _32807_ (
    .A1(\cpuregs[27] [12]),
    .A2(_00008_[0]),
    .ZN(_24679_)
  );
  INV_X1 _32808_ (
    .A(_24679_),
    .ZN(_24680_)
  );
  AND2_X1 _32809_ (
    .A1(\cpuregs[26] [12]),
    .A2(_22147_),
    .ZN(_24681_)
  );
  INV_X1 _32810_ (
    .A(_24681_),
    .ZN(_24682_)
  );
  AND2_X1 _32811_ (
    .A1(_22149_),
    .A2(_24682_),
    .ZN(_24683_)
  );
  AND2_X1 _32812_ (
    .A1(_24680_),
    .A2(_24683_),
    .ZN(_24684_)
  );
  INV_X1 _32813_ (
    .A(_24684_),
    .ZN(_24685_)
  );
  AND2_X1 _32814_ (
    .A1(\cpuregs[31] [12]),
    .A2(_00008_[0]),
    .ZN(_24686_)
  );
  INV_X1 _32815_ (
    .A(_24686_),
    .ZN(_24687_)
  );
  AND2_X1 _32816_ (
    .A1(\cpuregs[30] [12]),
    .A2(_22147_),
    .ZN(_24688_)
  );
  INV_X1 _32817_ (
    .A(_24688_),
    .ZN(_24689_)
  );
  AND2_X1 _32818_ (
    .A1(_00008_[2]),
    .A2(_24689_),
    .ZN(_24690_)
  );
  AND2_X1 _32819_ (
    .A1(_24687_),
    .A2(_24690_),
    .ZN(_24691_)
  );
  INV_X1 _32820_ (
    .A(_24691_),
    .ZN(_24692_)
  );
  AND2_X1 _32821_ (
    .A1(_24685_),
    .A2(_24692_),
    .ZN(_24693_)
  );
  INV_X1 _32822_ (
    .A(_24693_),
    .ZN(_24694_)
  );
  AND2_X1 _32823_ (
    .A1(_00008_[1]),
    .A2(_24694_),
    .ZN(_24695_)
  );
  INV_X1 _32824_ (
    .A(_24695_),
    .ZN(_24696_)
  );
  AND2_X1 _32825_ (
    .A1(\cpuregs[25] [12]),
    .A2(_00008_[0]),
    .ZN(_24697_)
  );
  INV_X1 _32826_ (
    .A(_24697_),
    .ZN(_24698_)
  );
  AND2_X1 _32827_ (
    .A1(\cpuregs[24] [12]),
    .A2(_22147_),
    .ZN(_24699_)
  );
  INV_X1 _32828_ (
    .A(_24699_),
    .ZN(_24700_)
  );
  AND2_X1 _32829_ (
    .A1(_22149_),
    .A2(_24700_),
    .ZN(_24701_)
  );
  AND2_X1 _32830_ (
    .A1(_24698_),
    .A2(_24701_),
    .ZN(_24702_)
  );
  INV_X1 _32831_ (
    .A(_24702_),
    .ZN(_24703_)
  );
  AND2_X1 _32832_ (
    .A1(\cpuregs[29] [12]),
    .A2(_00008_[0]),
    .ZN(_24704_)
  );
  INV_X1 _32833_ (
    .A(_24704_),
    .ZN(_24705_)
  );
  AND2_X1 _32834_ (
    .A1(\cpuregs[28] [12]),
    .A2(_22147_),
    .ZN(_24706_)
  );
  INV_X1 _32835_ (
    .A(_24706_),
    .ZN(_24707_)
  );
  AND2_X1 _32836_ (
    .A1(_00008_[2]),
    .A2(_24707_),
    .ZN(_24708_)
  );
  AND2_X1 _32837_ (
    .A1(_24705_),
    .A2(_24708_),
    .ZN(_24709_)
  );
  INV_X1 _32838_ (
    .A(_24709_),
    .ZN(_24710_)
  );
  AND2_X1 _32839_ (
    .A1(_24703_),
    .A2(_24710_),
    .ZN(_24711_)
  );
  INV_X1 _32840_ (
    .A(_24711_),
    .ZN(_24712_)
  );
  AND2_X1 _32841_ (
    .A1(_22148_),
    .A2(_24712_),
    .ZN(_24713_)
  );
  INV_X1 _32842_ (
    .A(_24713_),
    .ZN(_24714_)
  );
  AND2_X1 _32843_ (
    .A1(_00008_[3]),
    .A2(_24696_),
    .ZN(_24715_)
  );
  AND2_X1 _32844_ (
    .A1(_24714_),
    .A2(_24715_),
    .ZN(_24716_)
  );
  INV_X1 _32845_ (
    .A(_24716_),
    .ZN(_24717_)
  );
  AND2_X1 _32846_ (
    .A1(_22150_),
    .A2(_24678_),
    .ZN(_24718_)
  );
  AND2_X1 _32847_ (
    .A1(_24661_),
    .A2(_24718_),
    .ZN(_24719_)
  );
  INV_X1 _32848_ (
    .A(_24719_),
    .ZN(_24720_)
  );
  AND2_X1 _32849_ (
    .A1(_00008_[4]),
    .A2(_24720_),
    .ZN(_24721_)
  );
  AND2_X1 _32850_ (
    .A1(_24717_),
    .A2(_24721_),
    .ZN(_24722_)
  );
  INV_X1 _32851_ (
    .A(_24722_),
    .ZN(_24723_)
  );
  AND2_X1 _32852_ (
    .A1(\cpuregs[10] [12]),
    .A2(_22149_),
    .ZN(_24724_)
  );
  INV_X1 _32853_ (
    .A(_24724_),
    .ZN(_24725_)
  );
  AND2_X1 _32854_ (
    .A1(\cpuregs[14] [12]),
    .A2(_00008_[2]),
    .ZN(_24726_)
  );
  INV_X1 _32855_ (
    .A(_24726_),
    .ZN(_24727_)
  );
  AND2_X1 _32856_ (
    .A1(_22147_),
    .A2(_24727_),
    .ZN(_24728_)
  );
  AND2_X1 _32857_ (
    .A1(_24725_),
    .A2(_24728_),
    .ZN(_24729_)
  );
  INV_X1 _32858_ (
    .A(_24729_),
    .ZN(_24730_)
  );
  AND2_X1 _32859_ (
    .A1(\cpuregs[15] [12]),
    .A2(_00008_[2]),
    .ZN(_24731_)
  );
  INV_X1 _32860_ (
    .A(_24731_),
    .ZN(_24732_)
  );
  AND2_X1 _32861_ (
    .A1(\cpuregs[11] [12]),
    .A2(_22149_),
    .ZN(_24733_)
  );
  INV_X1 _32862_ (
    .A(_24733_),
    .ZN(_24734_)
  );
  AND2_X1 _32863_ (
    .A1(_00008_[0]),
    .A2(_24734_),
    .ZN(_24735_)
  );
  AND2_X1 _32864_ (
    .A1(_24732_),
    .A2(_24735_),
    .ZN(_24736_)
  );
  INV_X1 _32865_ (
    .A(_24736_),
    .ZN(_24737_)
  );
  AND2_X1 _32866_ (
    .A1(_24730_),
    .A2(_24737_),
    .ZN(_24738_)
  );
  AND2_X1 _32867_ (
    .A1(\cpuregs[2] [12]),
    .A2(_22149_),
    .ZN(_24739_)
  );
  INV_X1 _32868_ (
    .A(_24739_),
    .ZN(_24740_)
  );
  AND2_X1 _32869_ (
    .A1(\cpuregs[6] [12]),
    .A2(_00008_[2]),
    .ZN(_24741_)
  );
  INV_X1 _32870_ (
    .A(_24741_),
    .ZN(_24742_)
  );
  AND2_X1 _32871_ (
    .A1(_22147_),
    .A2(_24742_),
    .ZN(_24743_)
  );
  AND2_X1 _32872_ (
    .A1(_24740_),
    .A2(_24743_),
    .ZN(_24744_)
  );
  INV_X1 _32873_ (
    .A(_24744_),
    .ZN(_24745_)
  );
  AND2_X1 _32874_ (
    .A1(\cpuregs[3] [12]),
    .A2(_22149_),
    .ZN(_24746_)
  );
  INV_X1 _32875_ (
    .A(_24746_),
    .ZN(_24747_)
  );
  AND2_X1 _32876_ (
    .A1(\cpuregs[7] [12]),
    .A2(_00008_[2]),
    .ZN(_24748_)
  );
  INV_X1 _32877_ (
    .A(_24748_),
    .ZN(_24749_)
  );
  AND2_X1 _32878_ (
    .A1(_00008_[0]),
    .A2(_24749_),
    .ZN(_24750_)
  );
  AND2_X1 _32879_ (
    .A1(_24747_),
    .A2(_24750_),
    .ZN(_24751_)
  );
  INV_X1 _32880_ (
    .A(_24751_),
    .ZN(_24752_)
  );
  AND2_X1 _32881_ (
    .A1(_00008_[3]),
    .A2(_24738_),
    .ZN(_24753_)
  );
  INV_X1 _32882_ (
    .A(_24753_),
    .ZN(_24754_)
  );
  AND2_X1 _32883_ (
    .A1(_22150_),
    .A2(_24752_),
    .ZN(_24755_)
  );
  AND2_X1 _32884_ (
    .A1(_24745_),
    .A2(_24755_),
    .ZN(_24756_)
  );
  INV_X1 _32885_ (
    .A(_24756_),
    .ZN(_24757_)
  );
  AND2_X1 _32886_ (
    .A1(_24754_),
    .A2(_24757_),
    .ZN(_24758_)
  );
  INV_X1 _32887_ (
    .A(_24758_),
    .ZN(_24759_)
  );
  AND2_X1 _32888_ (
    .A1(\cpuregs[8] [12]),
    .A2(_22149_),
    .ZN(_24760_)
  );
  INV_X1 _32889_ (
    .A(_24760_),
    .ZN(_24761_)
  );
  AND2_X1 _32890_ (
    .A1(\cpuregs[12] [12]),
    .A2(_00008_[2]),
    .ZN(_24762_)
  );
  INV_X1 _32891_ (
    .A(_24762_),
    .ZN(_24763_)
  );
  AND2_X1 _32892_ (
    .A1(_22147_),
    .A2(_24763_),
    .ZN(_24764_)
  );
  AND2_X1 _32893_ (
    .A1(_24761_),
    .A2(_24764_),
    .ZN(_24765_)
  );
  INV_X1 _32894_ (
    .A(_24765_),
    .ZN(_24766_)
  );
  AND2_X1 _32895_ (
    .A1(\cpuregs[13] [12]),
    .A2(_00008_[2]),
    .ZN(_24767_)
  );
  INV_X1 _32896_ (
    .A(_24767_),
    .ZN(_24768_)
  );
  AND2_X1 _32897_ (
    .A1(\cpuregs[9] [12]),
    .A2(_22149_),
    .ZN(_24769_)
  );
  INV_X1 _32898_ (
    .A(_24769_),
    .ZN(_24770_)
  );
  AND2_X1 _32899_ (
    .A1(_00008_[0]),
    .A2(_24770_),
    .ZN(_24771_)
  );
  AND2_X1 _32900_ (
    .A1(_24768_),
    .A2(_24771_),
    .ZN(_24772_)
  );
  INV_X1 _32901_ (
    .A(_24772_),
    .ZN(_24773_)
  );
  AND2_X1 _32902_ (
    .A1(_24766_),
    .A2(_24773_),
    .ZN(_24774_)
  );
  AND2_X1 _32903_ (
    .A1(\cpuregs[0] [12]),
    .A2(_22149_),
    .ZN(_24775_)
  );
  INV_X1 _32904_ (
    .A(_24775_),
    .ZN(_24776_)
  );
  AND2_X1 _32905_ (
    .A1(\cpuregs[4] [12]),
    .A2(_00008_[2]),
    .ZN(_24777_)
  );
  INV_X1 _32906_ (
    .A(_24777_),
    .ZN(_24778_)
  );
  AND2_X1 _32907_ (
    .A1(_22147_),
    .A2(_24778_),
    .ZN(_24779_)
  );
  AND2_X1 _32908_ (
    .A1(_24776_),
    .A2(_24779_),
    .ZN(_24780_)
  );
  INV_X1 _32909_ (
    .A(_24780_),
    .ZN(_24781_)
  );
  AND2_X1 _32910_ (
    .A1(\cpuregs[1] [12]),
    .A2(_22149_),
    .ZN(_24782_)
  );
  INV_X1 _32911_ (
    .A(_24782_),
    .ZN(_24783_)
  );
  AND2_X1 _32912_ (
    .A1(\cpuregs[5] [12]),
    .A2(_00008_[2]),
    .ZN(_24784_)
  );
  INV_X1 _32913_ (
    .A(_24784_),
    .ZN(_24785_)
  );
  AND2_X1 _32914_ (
    .A1(_00008_[0]),
    .A2(_24785_),
    .ZN(_24786_)
  );
  AND2_X1 _32915_ (
    .A1(_24783_),
    .A2(_24786_),
    .ZN(_24787_)
  );
  INV_X1 _32916_ (
    .A(_24787_),
    .ZN(_24788_)
  );
  AND2_X1 _32917_ (
    .A1(_00008_[3]),
    .A2(_24774_),
    .ZN(_24789_)
  );
  INV_X1 _32918_ (
    .A(_24789_),
    .ZN(_24790_)
  );
  AND2_X1 _32919_ (
    .A1(_22150_),
    .A2(_24788_),
    .ZN(_24791_)
  );
  AND2_X1 _32920_ (
    .A1(_24781_),
    .A2(_24791_),
    .ZN(_24792_)
  );
  INV_X1 _32921_ (
    .A(_24792_),
    .ZN(_24793_)
  );
  AND2_X1 _32922_ (
    .A1(_24790_),
    .A2(_24793_),
    .ZN(_24794_)
  );
  INV_X1 _32923_ (
    .A(_24794_),
    .ZN(_24795_)
  );
  AND2_X1 _32924_ (
    .A1(_22148_),
    .A2(_24795_),
    .ZN(_24796_)
  );
  INV_X1 _32925_ (
    .A(_24796_),
    .ZN(_24797_)
  );
  AND2_X1 _32926_ (
    .A1(_00008_[1]),
    .A2(_24759_),
    .ZN(_24798_)
  );
  INV_X1 _32927_ (
    .A(_24798_),
    .ZN(_24799_)
  );
  AND2_X1 _32928_ (
    .A1(_24797_),
    .A2(_24799_),
    .ZN(_24800_)
  );
  AND2_X1 _32929_ (
    .A1(_22151_),
    .A2(_24800_),
    .ZN(_24801_)
  );
  INV_X1 _32930_ (
    .A(_24801_),
    .ZN(_24802_)
  );
  AND2_X1 _32931_ (
    .A1(_22546_),
    .A2(_24723_),
    .ZN(_24803_)
  );
  AND2_X1 _32932_ (
    .A1(_24802_),
    .A2(_24803_),
    .ZN(_24804_)
  );
  INV_X1 _32933_ (
    .A(_24804_),
    .ZN(_24805_)
  );
  AND2_X1 _32934_ (
    .A1(_24644_),
    .A2(_24805_),
    .ZN(_24806_)
  );
  INV_X1 _32935_ (
    .A(_24806_),
    .ZN(_24807_)
  );
  AND2_X1 _32936_ (
    .A1(_22271_),
    .A2(_24807_),
    .ZN(_24808_)
  );
  INV_X1 _32937_ (
    .A(_24808_),
    .ZN(_24809_)
  );
  AND2_X1 _32938_ (
    .A1(reg_op1[11]),
    .A2(_22285_),
    .ZN(_24810_)
  );
  INV_X1 _32939_ (
    .A(_24810_),
    .ZN(_24811_)
  );
  AND2_X1 _32940_ (
    .A1(_24199_),
    .A2(_24811_),
    .ZN(_24812_)
  );
  AND2_X1 _32941_ (
    .A1(reg_op1[16]),
    .A2(_22290_),
    .ZN(_24813_)
  );
  INV_X1 _32942_ (
    .A(_24813_),
    .ZN(_24814_)
  );
  AND2_X1 _32943_ (
    .A1(_24196_),
    .A2(_24814_),
    .ZN(_24815_)
  );
  AND2_X1 _32944_ (
    .A1(_22572_),
    .A2(_24812_),
    .ZN(_24816_)
  );
  INV_X1 _32945_ (
    .A(_24816_),
    .ZN(_24817_)
  );
  AND2_X1 _32946_ (
    .A1(_22573_),
    .A2(_24815_),
    .ZN(_24818_)
  );
  INV_X1 _32947_ (
    .A(_24818_),
    .ZN(_24819_)
  );
  AND2_X1 _32948_ (
    .A1(_22295_),
    .A2(_24819_),
    .ZN(_24820_)
  );
  AND2_X1 _32949_ (
    .A1(_24817_),
    .A2(_24820_),
    .ZN(_24821_)
  );
  INV_X1 _32950_ (
    .A(_24821_),
    .ZN(_24822_)
  );
  AND2_X1 _32951_ (
    .A1(_22333_),
    .A2(_24822_),
    .ZN(_24823_)
  );
  AND2_X1 _32952_ (
    .A1(_24809_),
    .A2(_24823_),
    .ZN(_24824_)
  );
  AND2_X1 _32953_ (
    .A1(_24436_),
    .A2(_24447_),
    .ZN(_24825_)
  );
  AND2_X1 _32954_ (
    .A1(_24445_),
    .A2(_24825_),
    .ZN(_24826_)
  );
  INV_X1 _32955_ (
    .A(_24826_),
    .ZN(_24827_)
  );
  AND2_X1 _32956_ (
    .A1(reg_op1[12]),
    .A2(decoded_imm[12]),
    .ZN(_24828_)
  );
  INV_X1 _32957_ (
    .A(_24828_),
    .ZN(_24829_)
  );
  AND2_X1 _32958_ (
    .A1(_21179_),
    .A2(_21997_),
    .ZN(_24830_)
  );
  INV_X1 _32959_ (
    .A(_24830_),
    .ZN(_24831_)
  );
  AND2_X1 _32960_ (
    .A1(_24829_),
    .A2(_24831_),
    .ZN(_24832_)
  );
  INV_X1 _32961_ (
    .A(_24832_),
    .ZN(_24833_)
  );
  AND2_X1 _32962_ (
    .A1(_24827_),
    .A2(_24832_),
    .ZN(_24834_)
  );
  INV_X1 _32963_ (
    .A(_24834_),
    .ZN(_24835_)
  );
  AND2_X1 _32964_ (
    .A1(_24826_),
    .A2(_24833_),
    .ZN(_24836_)
  );
  INV_X1 _32965_ (
    .A(_24836_),
    .ZN(_24837_)
  );
  AND2_X1 _32966_ (
    .A1(_22559_),
    .A2(_24837_),
    .ZN(_24838_)
  );
  AND2_X1 _32967_ (
    .A1(_24835_),
    .A2(_24838_),
    .ZN(_24839_)
  );
  INV_X1 _32968_ (
    .A(_24839_),
    .ZN(_24840_)
  );
  AND2_X1 _32969_ (
    .A1(_24824_),
    .A2(_24840_),
    .ZN(_24841_)
  );
  INV_X1 _32970_ (
    .A(_24841_),
    .ZN(_24842_)
  );
  AND2_X1 _32971_ (
    .A1(_24642_),
    .A2(_24842_),
    .ZN(_00069_)
  );
  AND2_X1 _32972_ (
    .A1(_21180_),
    .A2(_22334_),
    .ZN(_24843_)
  );
  INV_X1 _32973_ (
    .A(_24843_),
    .ZN(_24844_)
  );
  AND2_X1 _32974_ (
    .A1(reg_pc[13]),
    .A2(_22335_),
    .ZN(_24845_)
  );
  INV_X1 _32975_ (
    .A(_24845_),
    .ZN(_24846_)
  );
  AND2_X1 _32976_ (
    .A1(_21446_),
    .A2(_22149_),
    .ZN(_24847_)
  );
  INV_X1 _32977_ (
    .A(_24847_),
    .ZN(_24848_)
  );
  AND2_X1 _32978_ (
    .A1(_21657_),
    .A2(_00008_[2]),
    .ZN(_24849_)
  );
  INV_X1 _32979_ (
    .A(_24849_),
    .ZN(_24850_)
  );
  AND2_X1 _32980_ (
    .A1(_24848_),
    .A2(_24850_),
    .ZN(_24851_)
  );
  AND2_X1 _32981_ (
    .A1(_22147_),
    .A2(_24851_),
    .ZN(_24852_)
  );
  INV_X1 _32982_ (
    .A(_24852_),
    .ZN(_24853_)
  );
  AND2_X1 _32983_ (
    .A1(_21767_),
    .A2(_00008_[2]),
    .ZN(_24854_)
  );
  INV_X1 _32984_ (
    .A(_24854_),
    .ZN(_24855_)
  );
  AND2_X1 _32985_ (
    .A1(_21468_),
    .A2(_22149_),
    .ZN(_24856_)
  );
  INV_X1 _32986_ (
    .A(_24856_),
    .ZN(_24857_)
  );
  AND2_X1 _32987_ (
    .A1(_00008_[0]),
    .A2(_24855_),
    .ZN(_24858_)
  );
  AND2_X1 _32988_ (
    .A1(_24857_),
    .A2(_24858_),
    .ZN(_24859_)
  );
  INV_X1 _32989_ (
    .A(_24859_),
    .ZN(_24860_)
  );
  AND2_X1 _32990_ (
    .A1(_24853_),
    .A2(_24860_),
    .ZN(_24861_)
  );
  AND2_X1 _32991_ (
    .A1(_22148_),
    .A2(_24861_),
    .ZN(_24862_)
  );
  INV_X1 _32992_ (
    .A(_24862_),
    .ZN(_24863_)
  );
  AND2_X1 _32993_ (
    .A1(_21600_),
    .A2(_22149_),
    .ZN(_24864_)
  );
  INV_X1 _32994_ (
    .A(_24864_),
    .ZN(_24865_)
  );
  AND2_X1 _32995_ (
    .A1(_21420_),
    .A2(_00008_[2]),
    .ZN(_24866_)
  );
  INV_X1 _32996_ (
    .A(_24866_),
    .ZN(_24867_)
  );
  AND2_X1 _32997_ (
    .A1(_24865_),
    .A2(_24867_),
    .ZN(_24868_)
  );
  AND2_X1 _32998_ (
    .A1(_22147_),
    .A2(_24868_),
    .ZN(_24869_)
  );
  INV_X1 _32999_ (
    .A(_24869_),
    .ZN(_24870_)
  );
  AND2_X1 _33000_ (
    .A1(_21380_),
    .A2(_00008_[2]),
    .ZN(_24871_)
  );
  INV_X1 _33001_ (
    .A(_24871_),
    .ZN(_24872_)
  );
  AND2_X1 _33002_ (
    .A1(_21626_),
    .A2(_22149_),
    .ZN(_24873_)
  );
  INV_X1 _33003_ (
    .A(_24873_),
    .ZN(_24874_)
  );
  AND2_X1 _33004_ (
    .A1(_00008_[0]),
    .A2(_24874_),
    .ZN(_24875_)
  );
  AND2_X1 _33005_ (
    .A1(_24872_),
    .A2(_24875_),
    .ZN(_24876_)
  );
  INV_X1 _33006_ (
    .A(_24876_),
    .ZN(_24877_)
  );
  AND2_X1 _33007_ (
    .A1(_24870_),
    .A2(_24877_),
    .ZN(_24878_)
  );
  AND2_X1 _33008_ (
    .A1(_00008_[1]),
    .A2(_24878_),
    .ZN(_24879_)
  );
  INV_X1 _33009_ (
    .A(_24879_),
    .ZN(_24880_)
  );
  AND2_X1 _33010_ (
    .A1(_24863_),
    .A2(_24880_),
    .ZN(_24881_)
  );
  AND2_X1 _33011_ (
    .A1(_21876_),
    .A2(_22149_),
    .ZN(_24882_)
  );
  INV_X1 _33012_ (
    .A(_24882_),
    .ZN(_24883_)
  );
  AND2_X1 _33013_ (
    .A1(_21856_),
    .A2(_00008_[2]),
    .ZN(_24884_)
  );
  INV_X1 _33014_ (
    .A(_24884_),
    .ZN(_24885_)
  );
  AND2_X1 _33015_ (
    .A1(_24883_),
    .A2(_24885_),
    .ZN(_24886_)
  );
  AND2_X1 _33016_ (
    .A1(_22147_),
    .A2(_24886_),
    .ZN(_24887_)
  );
  INV_X1 _33017_ (
    .A(_24887_),
    .ZN(_24888_)
  );
  AND2_X1 _33018_ (
    .A1(_21944_),
    .A2(_00008_[2]),
    .ZN(_24889_)
  );
  INV_X1 _33019_ (
    .A(_24889_),
    .ZN(_24890_)
  );
  AND2_X1 _33020_ (
    .A1(_21928_),
    .A2(_22149_),
    .ZN(_24891_)
  );
  INV_X1 _33021_ (
    .A(_24891_),
    .ZN(_24892_)
  );
  AND2_X1 _33022_ (
    .A1(_00008_[0]),
    .A2(_24892_),
    .ZN(_24893_)
  );
  AND2_X1 _33023_ (
    .A1(_24890_),
    .A2(_24893_),
    .ZN(_24894_)
  );
  INV_X1 _33024_ (
    .A(_24894_),
    .ZN(_24895_)
  );
  AND2_X1 _33025_ (
    .A1(_24888_),
    .A2(_24895_),
    .ZN(_24896_)
  );
  AND2_X1 _33026_ (
    .A1(_00008_[1]),
    .A2(_24896_),
    .ZN(_24897_)
  );
  INV_X1 _33027_ (
    .A(_24897_),
    .ZN(_24898_)
  );
  AND2_X1 _33028_ (
    .A1(_21896_),
    .A2(_00008_[2]),
    .ZN(_24899_)
  );
  INV_X1 _33029_ (
    .A(_24899_),
    .ZN(_24900_)
  );
  AND2_X1 _33030_ (
    .A1(_21840_),
    .A2(_22149_),
    .ZN(_24901_)
  );
  INV_X1 _33031_ (
    .A(_24901_),
    .ZN(_24902_)
  );
  AND2_X1 _33032_ (
    .A1(_00008_[0]),
    .A2(_24902_),
    .ZN(_24903_)
  );
  AND2_X1 _33033_ (
    .A1(_24900_),
    .A2(_24903_),
    .ZN(_24904_)
  );
  INV_X1 _33034_ (
    .A(_24904_),
    .ZN(_24905_)
  );
  AND2_X1 _33035_ (
    .A1(_21574_),
    .A2(_22149_),
    .ZN(_24906_)
  );
  INV_X1 _33036_ (
    .A(_24906_),
    .ZN(_24907_)
  );
  AND2_X1 _33037_ (
    .A1(_21912_),
    .A2(_00008_[2]),
    .ZN(_24908_)
  );
  INV_X1 _33038_ (
    .A(_24908_),
    .ZN(_24909_)
  );
  AND2_X1 _33039_ (
    .A1(_24907_),
    .A2(_24909_),
    .ZN(_24910_)
  );
  AND2_X1 _33040_ (
    .A1(_22147_),
    .A2(_24910_),
    .ZN(_24911_)
  );
  INV_X1 _33041_ (
    .A(_24911_),
    .ZN(_24912_)
  );
  AND2_X1 _33042_ (
    .A1(_24905_),
    .A2(_24912_),
    .ZN(_24913_)
  );
  AND2_X1 _33043_ (
    .A1(_22148_),
    .A2(_24913_),
    .ZN(_24914_)
  );
  INV_X1 _33044_ (
    .A(_24914_),
    .ZN(_24915_)
  );
  AND2_X1 _33045_ (
    .A1(_00008_[3]),
    .A2(_24898_),
    .ZN(_24916_)
  );
  AND2_X1 _33046_ (
    .A1(_24915_),
    .A2(_24916_),
    .ZN(_24917_)
  );
  INV_X1 _33047_ (
    .A(_24917_),
    .ZN(_24918_)
  );
  AND2_X1 _33048_ (
    .A1(_22150_),
    .A2(_24881_),
    .ZN(_24919_)
  );
  INV_X1 _33049_ (
    .A(_24919_),
    .ZN(_24920_)
  );
  AND2_X1 _33050_ (
    .A1(_00008_[4]),
    .A2(_24920_),
    .ZN(_24921_)
  );
  AND2_X1 _33051_ (
    .A1(_24918_),
    .A2(_24921_),
    .ZN(_24922_)
  );
  INV_X1 _33052_ (
    .A(_24922_),
    .ZN(_24923_)
  );
  AND2_X1 _33053_ (
    .A1(\cpuregs[9] [13]),
    .A2(_22149_),
    .ZN(_24924_)
  );
  INV_X1 _33054_ (
    .A(_24924_),
    .ZN(_24925_)
  );
  AND2_X1 _33055_ (
    .A1(\cpuregs[13] [13]),
    .A2(_00008_[2]),
    .ZN(_24926_)
  );
  INV_X1 _33056_ (
    .A(_24926_),
    .ZN(_24927_)
  );
  AND2_X1 _33057_ (
    .A1(_22148_),
    .A2(_24927_),
    .ZN(_24928_)
  );
  AND2_X1 _33058_ (
    .A1(_24925_),
    .A2(_24928_),
    .ZN(_24929_)
  );
  INV_X1 _33059_ (
    .A(_24929_),
    .ZN(_24930_)
  );
  AND2_X1 _33060_ (
    .A1(\cpuregs[15] [13]),
    .A2(_00008_[2]),
    .ZN(_24931_)
  );
  INV_X1 _33061_ (
    .A(_24931_),
    .ZN(_24932_)
  );
  AND2_X1 _33062_ (
    .A1(\cpuregs[11] [13]),
    .A2(_22149_),
    .ZN(_24933_)
  );
  INV_X1 _33063_ (
    .A(_24933_),
    .ZN(_24934_)
  );
  AND2_X1 _33064_ (
    .A1(_00008_[1]),
    .A2(_24934_),
    .ZN(_24935_)
  );
  AND2_X1 _33065_ (
    .A1(_24932_),
    .A2(_24935_),
    .ZN(_24936_)
  );
  INV_X1 _33066_ (
    .A(_24936_),
    .ZN(_24937_)
  );
  AND2_X1 _33067_ (
    .A1(_24930_),
    .A2(_24937_),
    .ZN(_24938_)
  );
  INV_X1 _33068_ (
    .A(_24938_),
    .ZN(_24939_)
  );
  AND2_X1 _33069_ (
    .A1(_00008_[0]),
    .A2(_24939_),
    .ZN(_24940_)
  );
  INV_X1 _33070_ (
    .A(_24940_),
    .ZN(_24941_)
  );
  AND2_X1 _33071_ (
    .A1(\cpuregs[8] [13]),
    .A2(_22149_),
    .ZN(_24942_)
  );
  INV_X1 _33072_ (
    .A(_24942_),
    .ZN(_24943_)
  );
  AND2_X1 _33073_ (
    .A1(\cpuregs[12] [13]),
    .A2(_00008_[2]),
    .ZN(_24944_)
  );
  INV_X1 _33074_ (
    .A(_24944_),
    .ZN(_24945_)
  );
  AND2_X1 _33075_ (
    .A1(_22148_),
    .A2(_24945_),
    .ZN(_24946_)
  );
  AND2_X1 _33076_ (
    .A1(_24943_),
    .A2(_24946_),
    .ZN(_24947_)
  );
  INV_X1 _33077_ (
    .A(_24947_),
    .ZN(_24948_)
  );
  AND2_X1 _33078_ (
    .A1(\cpuregs[10] [13]),
    .A2(_22149_),
    .ZN(_24949_)
  );
  INV_X1 _33079_ (
    .A(_24949_),
    .ZN(_24950_)
  );
  AND2_X1 _33080_ (
    .A1(\cpuregs[14] [13]),
    .A2(_00008_[2]),
    .ZN(_24951_)
  );
  INV_X1 _33081_ (
    .A(_24951_),
    .ZN(_24952_)
  );
  AND2_X1 _33082_ (
    .A1(_00008_[1]),
    .A2(_24952_),
    .ZN(_24953_)
  );
  AND2_X1 _33083_ (
    .A1(_24950_),
    .A2(_24953_),
    .ZN(_24954_)
  );
  INV_X1 _33084_ (
    .A(_24954_),
    .ZN(_24955_)
  );
  AND2_X1 _33085_ (
    .A1(_24948_),
    .A2(_24955_),
    .ZN(_24956_)
  );
  INV_X1 _33086_ (
    .A(_24956_),
    .ZN(_24957_)
  );
  AND2_X1 _33087_ (
    .A1(_22147_),
    .A2(_24957_),
    .ZN(_24958_)
  );
  INV_X1 _33088_ (
    .A(_24958_),
    .ZN(_24959_)
  );
  AND2_X1 _33089_ (
    .A1(_24941_),
    .A2(_24959_),
    .ZN(_24960_)
  );
  INV_X1 _33090_ (
    .A(_24960_),
    .ZN(_24961_)
  );
  AND2_X1 _33091_ (
    .A1(_00008_[3]),
    .A2(_24961_),
    .ZN(_24962_)
  );
  INV_X1 _33092_ (
    .A(_24962_),
    .ZN(_24963_)
  );
  AND2_X1 _33093_ (
    .A1(_21789_),
    .A2(_00008_[2]),
    .ZN(_24964_)
  );
  INV_X1 _33094_ (
    .A(_24964_),
    .ZN(_24965_)
  );
  AND2_X1 _33095_ (
    .A1(_21497_),
    .A2(_22149_),
    .ZN(_24966_)
  );
  INV_X1 _33096_ (
    .A(_24966_),
    .ZN(_24967_)
  );
  AND2_X1 _33097_ (
    .A1(_00008_[0]),
    .A2(_24967_),
    .ZN(_24968_)
  );
  AND2_X1 _33098_ (
    .A1(_24965_),
    .A2(_24968_),
    .ZN(_24969_)
  );
  INV_X1 _33099_ (
    .A(_24969_),
    .ZN(_24970_)
  );
  AND2_X1 _33100_ (
    .A1(_21550_),
    .A2(_22149_),
    .ZN(_24971_)
  );
  INV_X1 _33101_ (
    .A(_24971_),
    .ZN(_24972_)
  );
  AND2_X1 _33102_ (
    .A1(_21816_),
    .A2(_00008_[2]),
    .ZN(_24973_)
  );
  INV_X1 _33103_ (
    .A(_24973_),
    .ZN(_24974_)
  );
  AND2_X1 _33104_ (
    .A1(_24972_),
    .A2(_24974_),
    .ZN(_24975_)
  );
  AND2_X1 _33105_ (
    .A1(_22147_),
    .A2(_24975_),
    .ZN(_24976_)
  );
  INV_X1 _33106_ (
    .A(_24976_),
    .ZN(_24977_)
  );
  AND2_X1 _33107_ (
    .A1(_24970_),
    .A2(_24977_),
    .ZN(_24978_)
  );
  AND2_X1 _33108_ (
    .A1(_00008_[1]),
    .A2(_24978_),
    .ZN(_24979_)
  );
  INV_X1 _33109_ (
    .A(_24979_),
    .ZN(_24980_)
  );
  AND2_X1 _33110_ (
    .A1(_21742_),
    .A2(_00008_[2]),
    .ZN(_24981_)
  );
  INV_X1 _33111_ (
    .A(_24981_),
    .ZN(_24982_)
  );
  AND2_X1 _33112_ (
    .A1(_21522_),
    .A2(_22149_),
    .ZN(_24983_)
  );
  INV_X1 _33113_ (
    .A(_24983_),
    .ZN(_24984_)
  );
  AND2_X1 _33114_ (
    .A1(_00008_[0]),
    .A2(_24984_),
    .ZN(_24985_)
  );
  AND2_X1 _33115_ (
    .A1(_24982_),
    .A2(_24985_),
    .ZN(_24986_)
  );
  INV_X1 _33116_ (
    .A(_24986_),
    .ZN(_24987_)
  );
  AND2_X1 _33117_ (
    .A1(_21963_),
    .A2(_22149_),
    .ZN(_24988_)
  );
  INV_X1 _33118_ (
    .A(_24988_),
    .ZN(_24989_)
  );
  AND2_X1 _33119_ (
    .A1(_21679_),
    .A2(_00008_[2]),
    .ZN(_24990_)
  );
  INV_X1 _33120_ (
    .A(_24990_),
    .ZN(_24991_)
  );
  AND2_X1 _33121_ (
    .A1(_24989_),
    .A2(_24991_),
    .ZN(_24992_)
  );
  AND2_X1 _33122_ (
    .A1(_22147_),
    .A2(_24992_),
    .ZN(_24993_)
  );
  INV_X1 _33123_ (
    .A(_24993_),
    .ZN(_24994_)
  );
  AND2_X1 _33124_ (
    .A1(_24987_),
    .A2(_24994_),
    .ZN(_24995_)
  );
  AND2_X1 _33125_ (
    .A1(_22148_),
    .A2(_24995_),
    .ZN(_24996_)
  );
  INV_X1 _33126_ (
    .A(_24996_),
    .ZN(_24997_)
  );
  AND2_X1 _33127_ (
    .A1(_24980_),
    .A2(_24997_),
    .ZN(_24998_)
  );
  INV_X1 _33128_ (
    .A(_24998_),
    .ZN(_24999_)
  );
  AND2_X1 _33129_ (
    .A1(_22150_),
    .A2(_24999_),
    .ZN(_25000_)
  );
  INV_X1 _33130_ (
    .A(_25000_),
    .ZN(_25001_)
  );
  AND2_X1 _33131_ (
    .A1(_24963_),
    .A2(_25001_),
    .ZN(_25002_)
  );
  INV_X1 _33132_ (
    .A(_25002_),
    .ZN(_25003_)
  );
  AND2_X1 _33133_ (
    .A1(_22151_),
    .A2(_25003_),
    .ZN(_25004_)
  );
  INV_X1 _33134_ (
    .A(_25004_),
    .ZN(_25005_)
  );
  AND2_X1 _33135_ (
    .A1(_22546_),
    .A2(_24923_),
    .ZN(_25006_)
  );
  AND2_X1 _33136_ (
    .A1(_25005_),
    .A2(_25006_),
    .ZN(_25007_)
  );
  INV_X1 _33137_ (
    .A(_25007_),
    .ZN(_25008_)
  );
  AND2_X1 _33138_ (
    .A1(_24846_),
    .A2(_25008_),
    .ZN(_25009_)
  );
  INV_X1 _33139_ (
    .A(_25009_),
    .ZN(_25010_)
  );
  AND2_X1 _33140_ (
    .A1(_22271_),
    .A2(_25010_),
    .ZN(_25011_)
  );
  INV_X1 _33141_ (
    .A(_25011_),
    .ZN(_25012_)
  );
  AND2_X1 _33142_ (
    .A1(reg_op1[12]),
    .A2(_22285_),
    .ZN(_25013_)
  );
  INV_X1 _33143_ (
    .A(_25013_),
    .ZN(_25014_)
  );
  AND2_X1 _33144_ (
    .A1(_24404_),
    .A2(_25014_),
    .ZN(_25015_)
  );
  AND2_X1 _33145_ (
    .A1(reg_op1[17]),
    .A2(_22290_),
    .ZN(_25016_)
  );
  INV_X1 _33146_ (
    .A(_25016_),
    .ZN(_25017_)
  );
  AND2_X1 _33147_ (
    .A1(_24401_),
    .A2(_25017_),
    .ZN(_25018_)
  );
  AND2_X1 _33148_ (
    .A1(_22572_),
    .A2(_25015_),
    .ZN(_25019_)
  );
  INV_X1 _33149_ (
    .A(_25019_),
    .ZN(_25020_)
  );
  AND2_X1 _33150_ (
    .A1(_22573_),
    .A2(_25018_),
    .ZN(_25021_)
  );
  INV_X1 _33151_ (
    .A(_25021_),
    .ZN(_25022_)
  );
  AND2_X1 _33152_ (
    .A1(_22295_),
    .A2(_25022_),
    .ZN(_25023_)
  );
  AND2_X1 _33153_ (
    .A1(_25020_),
    .A2(_25023_),
    .ZN(_25024_)
  );
  INV_X1 _33154_ (
    .A(_25024_),
    .ZN(_25025_)
  );
  AND2_X1 _33155_ (
    .A1(_22333_),
    .A2(_25025_),
    .ZN(_25026_)
  );
  AND2_X1 _33156_ (
    .A1(_25012_),
    .A2(_25026_),
    .ZN(_25027_)
  );
  AND2_X1 _33157_ (
    .A1(reg_op1[13]),
    .A2(decoded_imm[13]),
    .ZN(_25028_)
  );
  INV_X1 _33158_ (
    .A(_25028_),
    .ZN(_25029_)
  );
  AND2_X1 _33159_ (
    .A1(_21180_),
    .A2(_21996_),
    .ZN(_25030_)
  );
  INV_X1 _33160_ (
    .A(_25030_),
    .ZN(_25031_)
  );
  AND2_X1 _33161_ (
    .A1(_25029_),
    .A2(_25031_),
    .ZN(_25032_)
  );
  INV_X1 _33162_ (
    .A(_25032_),
    .ZN(_25033_)
  );
  AND2_X1 _33163_ (
    .A1(_24829_),
    .A2(_24835_),
    .ZN(_25034_)
  );
  INV_X1 _33164_ (
    .A(_25034_),
    .ZN(_25035_)
  );
  AND2_X1 _33165_ (
    .A1(_25032_),
    .A2(_25035_),
    .ZN(_25036_)
  );
  INV_X1 _33166_ (
    .A(_25036_),
    .ZN(_25037_)
  );
  AND2_X1 _33167_ (
    .A1(_25033_),
    .A2(_25034_),
    .ZN(_25038_)
  );
  INV_X1 _33168_ (
    .A(_25038_),
    .ZN(_25039_)
  );
  AND2_X1 _33169_ (
    .A1(_22559_),
    .A2(_25039_),
    .ZN(_25040_)
  );
  AND2_X1 _33170_ (
    .A1(_25037_),
    .A2(_25040_),
    .ZN(_25041_)
  );
  INV_X1 _33171_ (
    .A(_25041_),
    .ZN(_25042_)
  );
  AND2_X1 _33172_ (
    .A1(_25027_),
    .A2(_25042_),
    .ZN(_25043_)
  );
  INV_X1 _33173_ (
    .A(_25043_),
    .ZN(_25044_)
  );
  AND2_X1 _33174_ (
    .A1(_24844_),
    .A2(_25044_),
    .ZN(_00070_)
  );
  AND2_X1 _33175_ (
    .A1(_21181_),
    .A2(_22334_),
    .ZN(_25045_)
  );
  INV_X1 _33176_ (
    .A(_25045_),
    .ZN(_25046_)
  );
  AND2_X1 _33177_ (
    .A1(reg_pc[14]),
    .A2(_22335_),
    .ZN(_25047_)
  );
  INV_X1 _33178_ (
    .A(_25047_),
    .ZN(_25048_)
  );
  AND2_X1 _33179_ (
    .A1(\cpuregs[20] [14]),
    .A2(_00008_[2]),
    .ZN(_25049_)
  );
  INV_X1 _33180_ (
    .A(_25049_),
    .ZN(_25050_)
  );
  AND2_X1 _33181_ (
    .A1(\cpuregs[16] [14]),
    .A2(_22149_),
    .ZN(_25051_)
  );
  INV_X1 _33182_ (
    .A(_25051_),
    .ZN(_25052_)
  );
  AND2_X1 _33183_ (
    .A1(_25050_),
    .A2(_25052_),
    .ZN(_25053_)
  );
  AND2_X1 _33184_ (
    .A1(\cpuregs[21] [14]),
    .A2(_00008_[2]),
    .ZN(_25054_)
  );
  INV_X1 _33185_ (
    .A(_25054_),
    .ZN(_25055_)
  );
  AND2_X1 _33186_ (
    .A1(\cpuregs[17] [14]),
    .A2(_22149_),
    .ZN(_25056_)
  );
  INV_X1 _33187_ (
    .A(_25056_),
    .ZN(_25057_)
  );
  AND2_X1 _33188_ (
    .A1(_22147_),
    .A2(_25053_),
    .ZN(_25058_)
  );
  INV_X1 _33189_ (
    .A(_25058_),
    .ZN(_25059_)
  );
  AND2_X1 _33190_ (
    .A1(_00008_[0]),
    .A2(_25055_),
    .ZN(_25060_)
  );
  AND2_X1 _33191_ (
    .A1(_25057_),
    .A2(_25060_),
    .ZN(_25061_)
  );
  INV_X1 _33192_ (
    .A(_25061_),
    .ZN(_25062_)
  );
  AND2_X1 _33193_ (
    .A1(_25059_),
    .A2(_25062_),
    .ZN(_25063_)
  );
  INV_X1 _33194_ (
    .A(_25063_),
    .ZN(_25064_)
  );
  AND2_X1 _33195_ (
    .A1(_22150_),
    .A2(_25064_),
    .ZN(_25065_)
  );
  INV_X1 _33196_ (
    .A(_25065_),
    .ZN(_25066_)
  );
  AND2_X1 _33197_ (
    .A1(\cpuregs[28] [14]),
    .A2(_00008_[2]),
    .ZN(_25067_)
  );
  INV_X1 _33198_ (
    .A(_25067_),
    .ZN(_25068_)
  );
  AND2_X1 _33199_ (
    .A1(\cpuregs[24] [14]),
    .A2(_22149_),
    .ZN(_25069_)
  );
  INV_X1 _33200_ (
    .A(_25069_),
    .ZN(_25070_)
  );
  AND2_X1 _33201_ (
    .A1(_25068_),
    .A2(_25070_),
    .ZN(_25071_)
  );
  INV_X1 _33202_ (
    .A(_25071_),
    .ZN(_25072_)
  );
  AND2_X1 _33203_ (
    .A1(_22147_),
    .A2(_25072_),
    .ZN(_25073_)
  );
  INV_X1 _33204_ (
    .A(_25073_),
    .ZN(_25074_)
  );
  AND2_X1 _33205_ (
    .A1(\cpuregs[29] [14]),
    .A2(_00008_[2]),
    .ZN(_25075_)
  );
  INV_X1 _33206_ (
    .A(_25075_),
    .ZN(_25076_)
  );
  AND2_X1 _33207_ (
    .A1(\cpuregs[25] [14]),
    .A2(_22149_),
    .ZN(_25077_)
  );
  INV_X1 _33208_ (
    .A(_25077_),
    .ZN(_25078_)
  );
  AND2_X1 _33209_ (
    .A1(_25076_),
    .A2(_25078_),
    .ZN(_25079_)
  );
  INV_X1 _33210_ (
    .A(_25079_),
    .ZN(_25080_)
  );
  AND2_X1 _33211_ (
    .A1(_00008_[0]),
    .A2(_25080_),
    .ZN(_25081_)
  );
  INV_X1 _33212_ (
    .A(_25081_),
    .ZN(_25082_)
  );
  AND2_X1 _33213_ (
    .A1(_25074_),
    .A2(_25082_),
    .ZN(_25083_)
  );
  AND2_X1 _33214_ (
    .A1(_00008_[3]),
    .A2(_25083_),
    .ZN(_25084_)
  );
  INV_X1 _33215_ (
    .A(_25084_),
    .ZN(_25085_)
  );
  AND2_X1 _33216_ (
    .A1(\cpuregs[27] [14]),
    .A2(_00008_[0]),
    .ZN(_25086_)
  );
  INV_X1 _33217_ (
    .A(_25086_),
    .ZN(_25087_)
  );
  AND2_X1 _33218_ (
    .A1(\cpuregs[26] [14]),
    .A2(_22147_),
    .ZN(_25088_)
  );
  INV_X1 _33219_ (
    .A(_25088_),
    .ZN(_25089_)
  );
  AND2_X1 _33220_ (
    .A1(_22149_),
    .A2(_25089_),
    .ZN(_25090_)
  );
  AND2_X1 _33221_ (
    .A1(_25087_),
    .A2(_25090_),
    .ZN(_25091_)
  );
  INV_X1 _33222_ (
    .A(_25091_),
    .ZN(_25092_)
  );
  AND2_X1 _33223_ (
    .A1(\cpuregs[31] [14]),
    .A2(_00008_[0]),
    .ZN(_25093_)
  );
  INV_X1 _33224_ (
    .A(_25093_),
    .ZN(_25094_)
  );
  AND2_X1 _33225_ (
    .A1(\cpuregs[30] [14]),
    .A2(_22147_),
    .ZN(_25095_)
  );
  INV_X1 _33226_ (
    .A(_25095_),
    .ZN(_25096_)
  );
  AND2_X1 _33227_ (
    .A1(_00008_[2]),
    .A2(_25096_),
    .ZN(_25097_)
  );
  AND2_X1 _33228_ (
    .A1(_25094_),
    .A2(_25097_),
    .ZN(_25098_)
  );
  INV_X1 _33229_ (
    .A(_25098_),
    .ZN(_25099_)
  );
  AND2_X1 _33230_ (
    .A1(_25092_),
    .A2(_25099_),
    .ZN(_25100_)
  );
  INV_X1 _33231_ (
    .A(_25100_),
    .ZN(_25101_)
  );
  AND2_X1 _33232_ (
    .A1(_00008_[3]),
    .A2(_25101_),
    .ZN(_25102_)
  );
  INV_X1 _33233_ (
    .A(_25102_),
    .ZN(_25103_)
  );
  AND2_X1 _33234_ (
    .A1(\cpuregs[22] [14]),
    .A2(_00008_[2]),
    .ZN(_25104_)
  );
  INV_X1 _33235_ (
    .A(_25104_),
    .ZN(_25105_)
  );
  AND2_X1 _33236_ (
    .A1(\cpuregs[18] [14]),
    .A2(_22149_),
    .ZN(_25106_)
  );
  INV_X1 _33237_ (
    .A(_25106_),
    .ZN(_25107_)
  );
  AND2_X1 _33238_ (
    .A1(_22147_),
    .A2(_25107_),
    .ZN(_25108_)
  );
  AND2_X1 _33239_ (
    .A1(_25105_),
    .A2(_25108_),
    .ZN(_25109_)
  );
  INV_X1 _33240_ (
    .A(_25109_),
    .ZN(_25110_)
  );
  AND2_X1 _33241_ (
    .A1(\cpuregs[19] [14]),
    .A2(_22149_),
    .ZN(_25111_)
  );
  INV_X1 _33242_ (
    .A(_25111_),
    .ZN(_25112_)
  );
  AND2_X1 _33243_ (
    .A1(\cpuregs[23] [14]),
    .A2(_00008_[2]),
    .ZN(_25113_)
  );
  INV_X1 _33244_ (
    .A(_25113_),
    .ZN(_25114_)
  );
  AND2_X1 _33245_ (
    .A1(_00008_[0]),
    .A2(_25114_),
    .ZN(_25115_)
  );
  AND2_X1 _33246_ (
    .A1(_25112_),
    .A2(_25115_),
    .ZN(_25116_)
  );
  INV_X1 _33247_ (
    .A(_25116_),
    .ZN(_25117_)
  );
  AND2_X1 _33248_ (
    .A1(_25110_),
    .A2(_25117_),
    .ZN(_25118_)
  );
  INV_X1 _33249_ (
    .A(_25118_),
    .ZN(_25119_)
  );
  AND2_X1 _33250_ (
    .A1(_22150_),
    .A2(_25119_),
    .ZN(_25120_)
  );
  INV_X1 _33251_ (
    .A(_25120_),
    .ZN(_25121_)
  );
  AND2_X1 _33252_ (
    .A1(_25103_),
    .A2(_25121_),
    .ZN(_25122_)
  );
  AND2_X1 _33253_ (
    .A1(_00008_[1]),
    .A2(_25122_),
    .ZN(_25123_)
  );
  INV_X1 _33254_ (
    .A(_25123_),
    .ZN(_25124_)
  );
  AND2_X1 _33255_ (
    .A1(_22148_),
    .A2(_25085_),
    .ZN(_25125_)
  );
  AND2_X1 _33256_ (
    .A1(_25066_),
    .A2(_25125_),
    .ZN(_25126_)
  );
  INV_X1 _33257_ (
    .A(_25126_),
    .ZN(_25127_)
  );
  AND2_X1 _33258_ (
    .A1(_00008_[4]),
    .A2(_25127_),
    .ZN(_25128_)
  );
  AND2_X1 _33259_ (
    .A1(_25124_),
    .A2(_25128_),
    .ZN(_25129_)
  );
  INV_X1 _33260_ (
    .A(_25129_),
    .ZN(_25130_)
  );
  AND2_X1 _33261_ (
    .A1(\cpuregs[9] [14]),
    .A2(_22149_),
    .ZN(_25131_)
  );
  INV_X1 _33262_ (
    .A(_25131_),
    .ZN(_25132_)
  );
  AND2_X1 _33263_ (
    .A1(\cpuregs[13] [14]),
    .A2(_00008_[2]),
    .ZN(_25133_)
  );
  INV_X1 _33264_ (
    .A(_25133_),
    .ZN(_25134_)
  );
  AND2_X1 _33265_ (
    .A1(_22148_),
    .A2(_25134_),
    .ZN(_25135_)
  );
  AND2_X1 _33266_ (
    .A1(_25132_),
    .A2(_25135_),
    .ZN(_25136_)
  );
  INV_X1 _33267_ (
    .A(_25136_),
    .ZN(_25137_)
  );
  AND2_X1 _33268_ (
    .A1(\cpuregs[15] [14]),
    .A2(_00008_[2]),
    .ZN(_25138_)
  );
  INV_X1 _33269_ (
    .A(_25138_),
    .ZN(_25139_)
  );
  AND2_X1 _33270_ (
    .A1(\cpuregs[11] [14]),
    .A2(_22149_),
    .ZN(_25140_)
  );
  INV_X1 _33271_ (
    .A(_25140_),
    .ZN(_25141_)
  );
  AND2_X1 _33272_ (
    .A1(_00008_[1]),
    .A2(_25141_),
    .ZN(_25142_)
  );
  AND2_X1 _33273_ (
    .A1(_25139_),
    .A2(_25142_),
    .ZN(_25143_)
  );
  INV_X1 _33274_ (
    .A(_25143_),
    .ZN(_25144_)
  );
  AND2_X1 _33275_ (
    .A1(_25137_),
    .A2(_25144_),
    .ZN(_25145_)
  );
  INV_X1 _33276_ (
    .A(_25145_),
    .ZN(_25146_)
  );
  AND2_X1 _33277_ (
    .A1(_00008_[0]),
    .A2(_25146_),
    .ZN(_25147_)
  );
  INV_X1 _33278_ (
    .A(_25147_),
    .ZN(_25148_)
  );
  AND2_X1 _33279_ (
    .A1(\cpuregs[8] [14]),
    .A2(_22149_),
    .ZN(_25149_)
  );
  INV_X1 _33280_ (
    .A(_25149_),
    .ZN(_25150_)
  );
  AND2_X1 _33281_ (
    .A1(\cpuregs[12] [14]),
    .A2(_00008_[2]),
    .ZN(_25151_)
  );
  INV_X1 _33282_ (
    .A(_25151_),
    .ZN(_25152_)
  );
  AND2_X1 _33283_ (
    .A1(_22148_),
    .A2(_25152_),
    .ZN(_25153_)
  );
  AND2_X1 _33284_ (
    .A1(_25150_),
    .A2(_25153_),
    .ZN(_25154_)
  );
  INV_X1 _33285_ (
    .A(_25154_),
    .ZN(_25155_)
  );
  AND2_X1 _33286_ (
    .A1(\cpuregs[10] [14]),
    .A2(_22149_),
    .ZN(_25156_)
  );
  INV_X1 _33287_ (
    .A(_25156_),
    .ZN(_25157_)
  );
  AND2_X1 _33288_ (
    .A1(\cpuregs[14] [14]),
    .A2(_00008_[2]),
    .ZN(_25158_)
  );
  INV_X1 _33289_ (
    .A(_25158_),
    .ZN(_25159_)
  );
  AND2_X1 _33290_ (
    .A1(_00008_[1]),
    .A2(_25159_),
    .ZN(_25160_)
  );
  AND2_X1 _33291_ (
    .A1(_25157_),
    .A2(_25160_),
    .ZN(_25161_)
  );
  INV_X1 _33292_ (
    .A(_25161_),
    .ZN(_25162_)
  );
  AND2_X1 _33293_ (
    .A1(_25155_),
    .A2(_25162_),
    .ZN(_25163_)
  );
  INV_X1 _33294_ (
    .A(_25163_),
    .ZN(_25164_)
  );
  AND2_X1 _33295_ (
    .A1(_22147_),
    .A2(_25164_),
    .ZN(_25165_)
  );
  INV_X1 _33296_ (
    .A(_25165_),
    .ZN(_25166_)
  );
  AND2_X1 _33297_ (
    .A1(_25148_),
    .A2(_25166_),
    .ZN(_25167_)
  );
  INV_X1 _33298_ (
    .A(_25167_),
    .ZN(_25168_)
  );
  AND2_X1 _33299_ (
    .A1(_00008_[3]),
    .A2(_25168_),
    .ZN(_25169_)
  );
  INV_X1 _33300_ (
    .A(_25169_),
    .ZN(_25170_)
  );
  AND2_X1 _33301_ (
    .A1(_21743_),
    .A2(_00008_[2]),
    .ZN(_25171_)
  );
  INV_X1 _33302_ (
    .A(_25171_),
    .ZN(_25172_)
  );
  AND2_X1 _33303_ (
    .A1(_21523_),
    .A2(_22149_),
    .ZN(_25173_)
  );
  INV_X1 _33304_ (
    .A(_25173_),
    .ZN(_25174_)
  );
  AND2_X1 _33305_ (
    .A1(_00008_[0]),
    .A2(_25174_),
    .ZN(_25175_)
  );
  AND2_X1 _33306_ (
    .A1(_25172_),
    .A2(_25175_),
    .ZN(_25176_)
  );
  INV_X1 _33307_ (
    .A(_25176_),
    .ZN(_25177_)
  );
  AND2_X1 _33308_ (
    .A1(_21964_),
    .A2(_22149_),
    .ZN(_25178_)
  );
  INV_X1 _33309_ (
    .A(_25178_),
    .ZN(_25179_)
  );
  AND2_X1 _33310_ (
    .A1(_21680_),
    .A2(_00008_[2]),
    .ZN(_25180_)
  );
  INV_X1 _33311_ (
    .A(_25180_),
    .ZN(_25181_)
  );
  AND2_X1 _33312_ (
    .A1(_25179_),
    .A2(_25181_),
    .ZN(_25182_)
  );
  AND2_X1 _33313_ (
    .A1(_22147_),
    .A2(_25182_),
    .ZN(_25183_)
  );
  INV_X1 _33314_ (
    .A(_25183_),
    .ZN(_25184_)
  );
  AND2_X1 _33315_ (
    .A1(_25177_),
    .A2(_25184_),
    .ZN(_25185_)
  );
  AND2_X1 _33316_ (
    .A1(_22148_),
    .A2(_25185_),
    .ZN(_25186_)
  );
  INV_X1 _33317_ (
    .A(_25186_),
    .ZN(_25187_)
  );
  AND2_X1 _33318_ (
    .A1(_21790_),
    .A2(_00008_[2]),
    .ZN(_25188_)
  );
  INV_X1 _33319_ (
    .A(_25188_),
    .ZN(_25189_)
  );
  AND2_X1 _33320_ (
    .A1(_21498_),
    .A2(_22149_),
    .ZN(_25190_)
  );
  INV_X1 _33321_ (
    .A(_25190_),
    .ZN(_25191_)
  );
  AND2_X1 _33322_ (
    .A1(_00008_[0]),
    .A2(_25191_),
    .ZN(_25192_)
  );
  AND2_X1 _33323_ (
    .A1(_25189_),
    .A2(_25192_),
    .ZN(_25193_)
  );
  INV_X1 _33324_ (
    .A(_25193_),
    .ZN(_25194_)
  );
  AND2_X1 _33325_ (
    .A1(_21551_),
    .A2(_22149_),
    .ZN(_25195_)
  );
  INV_X1 _33326_ (
    .A(_25195_),
    .ZN(_25196_)
  );
  AND2_X1 _33327_ (
    .A1(_21817_),
    .A2(_00008_[2]),
    .ZN(_25197_)
  );
  INV_X1 _33328_ (
    .A(_25197_),
    .ZN(_25198_)
  );
  AND2_X1 _33329_ (
    .A1(_25196_),
    .A2(_25198_),
    .ZN(_25199_)
  );
  AND2_X1 _33330_ (
    .A1(_22147_),
    .A2(_25199_),
    .ZN(_25200_)
  );
  INV_X1 _33331_ (
    .A(_25200_),
    .ZN(_25201_)
  );
  AND2_X1 _33332_ (
    .A1(_25194_),
    .A2(_25201_),
    .ZN(_25202_)
  );
  AND2_X1 _33333_ (
    .A1(_00008_[1]),
    .A2(_25202_),
    .ZN(_25203_)
  );
  INV_X1 _33334_ (
    .A(_25203_),
    .ZN(_25204_)
  );
  AND2_X1 _33335_ (
    .A1(_25187_),
    .A2(_25204_),
    .ZN(_25205_)
  );
  INV_X1 _33336_ (
    .A(_25205_),
    .ZN(_25206_)
  );
  AND2_X1 _33337_ (
    .A1(_22150_),
    .A2(_25206_),
    .ZN(_25207_)
  );
  INV_X1 _33338_ (
    .A(_25207_),
    .ZN(_25208_)
  );
  AND2_X1 _33339_ (
    .A1(_25170_),
    .A2(_25208_),
    .ZN(_25209_)
  );
  INV_X1 _33340_ (
    .A(_25209_),
    .ZN(_25210_)
  );
  AND2_X1 _33341_ (
    .A1(_22151_),
    .A2(_25210_),
    .ZN(_25211_)
  );
  INV_X1 _33342_ (
    .A(_25211_),
    .ZN(_25212_)
  );
  AND2_X1 _33343_ (
    .A1(_22546_),
    .A2(_25130_),
    .ZN(_25213_)
  );
  AND2_X1 _33344_ (
    .A1(_25212_),
    .A2(_25213_),
    .ZN(_25214_)
  );
  INV_X1 _33345_ (
    .A(_25214_),
    .ZN(_25215_)
  );
  AND2_X1 _33346_ (
    .A1(_25048_),
    .A2(_25215_),
    .ZN(_25216_)
  );
  INV_X1 _33347_ (
    .A(_25216_),
    .ZN(_25217_)
  );
  AND2_X1 _33348_ (
    .A1(_22271_),
    .A2(_25217_),
    .ZN(_25218_)
  );
  INV_X1 _33349_ (
    .A(_25218_),
    .ZN(_25219_)
  );
  AND2_X1 _33350_ (
    .A1(reg_op1[13]),
    .A2(_22285_),
    .ZN(_25220_)
  );
  INV_X1 _33351_ (
    .A(_25220_),
    .ZN(_25221_)
  );
  AND2_X1 _33352_ (
    .A1(_24628_),
    .A2(_25221_),
    .ZN(_25222_)
  );
  AND2_X1 _33353_ (
    .A1(reg_op1[18]),
    .A2(_22290_),
    .ZN(_25223_)
  );
  INV_X1 _33354_ (
    .A(_25223_),
    .ZN(_25224_)
  );
  AND2_X1 _33355_ (
    .A1(_24625_),
    .A2(_25224_),
    .ZN(_25225_)
  );
  AND2_X1 _33356_ (
    .A1(_22572_),
    .A2(_25222_),
    .ZN(_25226_)
  );
  INV_X1 _33357_ (
    .A(_25226_),
    .ZN(_25227_)
  );
  AND2_X1 _33358_ (
    .A1(_22573_),
    .A2(_25225_),
    .ZN(_25228_)
  );
  INV_X1 _33359_ (
    .A(_25228_),
    .ZN(_25229_)
  );
  AND2_X1 _33360_ (
    .A1(_22295_),
    .A2(_25229_),
    .ZN(_25230_)
  );
  AND2_X1 _33361_ (
    .A1(_25227_),
    .A2(_25230_),
    .ZN(_25231_)
  );
  INV_X1 _33362_ (
    .A(_25231_),
    .ZN(_25232_)
  );
  AND2_X1 _33363_ (
    .A1(_22333_),
    .A2(_25232_),
    .ZN(_25233_)
  );
  AND2_X1 _33364_ (
    .A1(_25219_),
    .A2(_25233_),
    .ZN(_25234_)
  );
  AND2_X1 _33365_ (
    .A1(_25029_),
    .A2(_25037_),
    .ZN(_25235_)
  );
  INV_X1 _33366_ (
    .A(_25235_),
    .ZN(_25236_)
  );
  AND2_X1 _33367_ (
    .A1(reg_op1[14]),
    .A2(decoded_imm[14]),
    .ZN(_25237_)
  );
  INV_X1 _33368_ (
    .A(_25237_),
    .ZN(_25238_)
  );
  AND2_X1 _33369_ (
    .A1(_21181_),
    .A2(_21995_),
    .ZN(_25239_)
  );
  INV_X1 _33370_ (
    .A(_25239_),
    .ZN(_25240_)
  );
  AND2_X1 _33371_ (
    .A1(_25238_),
    .A2(_25240_),
    .ZN(_25241_)
  );
  INV_X1 _33372_ (
    .A(_25241_),
    .ZN(_25242_)
  );
  AND2_X1 _33373_ (
    .A1(_25236_),
    .A2(_25241_),
    .ZN(_25243_)
  );
  INV_X1 _33374_ (
    .A(_25243_),
    .ZN(_25244_)
  );
  AND2_X1 _33375_ (
    .A1(_25235_),
    .A2(_25242_),
    .ZN(_25245_)
  );
  INV_X1 _33376_ (
    .A(_25245_),
    .ZN(_25246_)
  );
  AND2_X1 _33377_ (
    .A1(_22559_),
    .A2(_25246_),
    .ZN(_25247_)
  );
  AND2_X1 _33378_ (
    .A1(_25244_),
    .A2(_25247_),
    .ZN(_25248_)
  );
  INV_X1 _33379_ (
    .A(_25248_),
    .ZN(_25249_)
  );
  AND2_X1 _33380_ (
    .A1(_25234_),
    .A2(_25249_),
    .ZN(_25250_)
  );
  INV_X1 _33381_ (
    .A(_25250_),
    .ZN(_25251_)
  );
  AND2_X1 _33382_ (
    .A1(_25046_),
    .A2(_25251_),
    .ZN(_00071_)
  );
  AND2_X1 _33383_ (
    .A1(_21182_),
    .A2(_22334_),
    .ZN(_25252_)
  );
  INV_X1 _33384_ (
    .A(_25252_),
    .ZN(_25253_)
  );
  AND2_X1 _33385_ (
    .A1(reg_pc[15]),
    .A2(_22335_),
    .ZN(_25254_)
  );
  INV_X1 _33386_ (
    .A(_25254_),
    .ZN(_25255_)
  );
  AND2_X1 _33387_ (
    .A1(\cpuregs[12] [15]),
    .A2(_00008_[2]),
    .ZN(_25256_)
  );
  INV_X1 _33388_ (
    .A(_25256_),
    .ZN(_25257_)
  );
  AND2_X1 _33389_ (
    .A1(\cpuregs[8] [15]),
    .A2(_22149_),
    .ZN(_25258_)
  );
  INV_X1 _33390_ (
    .A(_25258_),
    .ZN(_25259_)
  );
  AND2_X1 _33391_ (
    .A1(_25257_),
    .A2(_25259_),
    .ZN(_25260_)
  );
  INV_X1 _33392_ (
    .A(_25260_),
    .ZN(_25261_)
  );
  AND2_X1 _33393_ (
    .A1(_22147_),
    .A2(_25261_),
    .ZN(_25262_)
  );
  INV_X1 _33394_ (
    .A(_25262_),
    .ZN(_25263_)
  );
  AND2_X1 _33395_ (
    .A1(\cpuregs[13] [15]),
    .A2(_00008_[2]),
    .ZN(_25264_)
  );
  INV_X1 _33396_ (
    .A(_25264_),
    .ZN(_25265_)
  );
  AND2_X1 _33397_ (
    .A1(\cpuregs[9] [15]),
    .A2(_22149_),
    .ZN(_25266_)
  );
  INV_X1 _33398_ (
    .A(_25266_),
    .ZN(_25267_)
  );
  AND2_X1 _33399_ (
    .A1(_25265_),
    .A2(_25267_),
    .ZN(_25268_)
  );
  INV_X1 _33400_ (
    .A(_25268_),
    .ZN(_25269_)
  );
  AND2_X1 _33401_ (
    .A1(_00008_[0]),
    .A2(_25269_),
    .ZN(_25270_)
  );
  INV_X1 _33402_ (
    .A(_25270_),
    .ZN(_25271_)
  );
  AND2_X1 _33403_ (
    .A1(_25263_),
    .A2(_25271_),
    .ZN(_25272_)
  );
  AND2_X1 _33404_ (
    .A1(_22148_),
    .A2(_25272_),
    .ZN(_25273_)
  );
  INV_X1 _33405_ (
    .A(_25273_),
    .ZN(_25274_)
  );
  AND2_X1 _33406_ (
    .A1(_21706_),
    .A2(_22149_),
    .ZN(_25275_)
  );
  INV_X1 _33407_ (
    .A(_25275_),
    .ZN(_25276_)
  );
  AND2_X1 _33408_ (
    .A1(_21396_),
    .A2(_00008_[2]),
    .ZN(_25277_)
  );
  INV_X1 _33409_ (
    .A(_25277_),
    .ZN(_25278_)
  );
  AND2_X1 _33410_ (
    .A1(_25276_),
    .A2(_25278_),
    .ZN(_25279_)
  );
  AND2_X1 _33411_ (
    .A1(_22147_),
    .A2(_25279_),
    .ZN(_25280_)
  );
  INV_X1 _33412_ (
    .A(_25280_),
    .ZN(_25281_)
  );
  AND2_X1 _33413_ (
    .A1(\cpuregs[11] [15]),
    .A2(_22149_),
    .ZN(_25282_)
  );
  INV_X1 _33414_ (
    .A(_25282_),
    .ZN(_25283_)
  );
  AND2_X1 _33415_ (
    .A1(\cpuregs[15] [15]),
    .A2(_00008_[2]),
    .ZN(_25284_)
  );
  INV_X1 _33416_ (
    .A(_25284_),
    .ZN(_25285_)
  );
  AND2_X1 _33417_ (
    .A1(_25283_),
    .A2(_25285_),
    .ZN(_25286_)
  );
  INV_X1 _33418_ (
    .A(_25286_),
    .ZN(_25287_)
  );
  AND2_X1 _33419_ (
    .A1(_00008_[0]),
    .A2(_25287_),
    .ZN(_25288_)
  );
  INV_X1 _33420_ (
    .A(_25288_),
    .ZN(_25289_)
  );
  AND2_X1 _33421_ (
    .A1(_25281_),
    .A2(_25289_),
    .ZN(_25290_)
  );
  AND2_X1 _33422_ (
    .A1(_00008_[1]),
    .A2(_25290_),
    .ZN(_25291_)
  );
  INV_X1 _33423_ (
    .A(_25291_),
    .ZN(_25292_)
  );
  AND2_X1 _33424_ (
    .A1(_25274_),
    .A2(_25292_),
    .ZN(_25293_)
  );
  AND2_X1 _33425_ (
    .A1(_21877_),
    .A2(_22149_),
    .ZN(_25294_)
  );
  INV_X1 _33426_ (
    .A(_25294_),
    .ZN(_25295_)
  );
  AND2_X1 _33427_ (
    .A1(_21857_),
    .A2(_00008_[2]),
    .ZN(_25296_)
  );
  INV_X1 _33428_ (
    .A(_25296_),
    .ZN(_25297_)
  );
  AND2_X1 _33429_ (
    .A1(_25295_),
    .A2(_25297_),
    .ZN(_25298_)
  );
  AND2_X1 _33430_ (
    .A1(_22147_),
    .A2(_25298_),
    .ZN(_25299_)
  );
  INV_X1 _33431_ (
    .A(_25299_),
    .ZN(_25300_)
  );
  AND2_X1 _33432_ (
    .A1(_21945_),
    .A2(_00008_[2]),
    .ZN(_25301_)
  );
  INV_X1 _33433_ (
    .A(_25301_),
    .ZN(_25302_)
  );
  AND2_X1 _33434_ (
    .A1(_21929_),
    .A2(_22149_),
    .ZN(_25303_)
  );
  INV_X1 _33435_ (
    .A(_25303_),
    .ZN(_25304_)
  );
  AND2_X1 _33436_ (
    .A1(_00008_[0]),
    .A2(_25304_),
    .ZN(_25305_)
  );
  AND2_X1 _33437_ (
    .A1(_25302_),
    .A2(_25305_),
    .ZN(_25306_)
  );
  INV_X1 _33438_ (
    .A(_25306_),
    .ZN(_25307_)
  );
  AND2_X1 _33439_ (
    .A1(_25300_),
    .A2(_25307_),
    .ZN(_25308_)
  );
  AND2_X1 _33440_ (
    .A1(_00008_[1]),
    .A2(_25308_),
    .ZN(_25309_)
  );
  INV_X1 _33441_ (
    .A(_25309_),
    .ZN(_25310_)
  );
  AND2_X1 _33442_ (
    .A1(_21897_),
    .A2(_00008_[2]),
    .ZN(_25311_)
  );
  INV_X1 _33443_ (
    .A(_25311_),
    .ZN(_25312_)
  );
  AND2_X1 _33444_ (
    .A1(_21841_),
    .A2(_22149_),
    .ZN(_25313_)
  );
  INV_X1 _33445_ (
    .A(_25313_),
    .ZN(_25314_)
  );
  AND2_X1 _33446_ (
    .A1(_00008_[0]),
    .A2(_25314_),
    .ZN(_25315_)
  );
  AND2_X1 _33447_ (
    .A1(_25312_),
    .A2(_25315_),
    .ZN(_25316_)
  );
  INV_X1 _33448_ (
    .A(_25316_),
    .ZN(_25317_)
  );
  AND2_X1 _33449_ (
    .A1(_21575_),
    .A2(_22149_),
    .ZN(_25318_)
  );
  INV_X1 _33450_ (
    .A(_25318_),
    .ZN(_25319_)
  );
  AND2_X1 _33451_ (
    .A1(_21913_),
    .A2(_00008_[2]),
    .ZN(_25320_)
  );
  INV_X1 _33452_ (
    .A(_25320_),
    .ZN(_25321_)
  );
  AND2_X1 _33453_ (
    .A1(_25319_),
    .A2(_25321_),
    .ZN(_25322_)
  );
  AND2_X1 _33454_ (
    .A1(_22147_),
    .A2(_25322_),
    .ZN(_25323_)
  );
  INV_X1 _33455_ (
    .A(_25323_),
    .ZN(_25324_)
  );
  AND2_X1 _33456_ (
    .A1(_25317_),
    .A2(_25324_),
    .ZN(_25325_)
  );
  AND2_X1 _33457_ (
    .A1(_22148_),
    .A2(_25325_),
    .ZN(_25326_)
  );
  INV_X1 _33458_ (
    .A(_25326_),
    .ZN(_25327_)
  );
  AND2_X1 _33459_ (
    .A1(_00008_[4]),
    .A2(_25310_),
    .ZN(_25328_)
  );
  AND2_X1 _33460_ (
    .A1(_25327_),
    .A2(_25328_),
    .ZN(_25329_)
  );
  INV_X1 _33461_ (
    .A(_25329_),
    .ZN(_25330_)
  );
  AND2_X1 _33462_ (
    .A1(_22151_),
    .A2(_25293_),
    .ZN(_25331_)
  );
  INV_X1 _33463_ (
    .A(_25331_),
    .ZN(_25332_)
  );
  AND2_X1 _33464_ (
    .A1(_25330_),
    .A2(_25332_),
    .ZN(_25333_)
  );
  AND2_X1 _33465_ (
    .A1(_00008_[3]),
    .A2(_25333_),
    .ZN(_25334_)
  );
  INV_X1 _33466_ (
    .A(_25334_),
    .ZN(_25335_)
  );
  AND2_X1 _33467_ (
    .A1(_21447_),
    .A2(_22149_),
    .ZN(_25336_)
  );
  INV_X1 _33468_ (
    .A(_25336_),
    .ZN(_25337_)
  );
  AND2_X1 _33469_ (
    .A1(_21658_),
    .A2(_00008_[2]),
    .ZN(_25338_)
  );
  INV_X1 _33470_ (
    .A(_25338_),
    .ZN(_25339_)
  );
  AND2_X1 _33471_ (
    .A1(_25337_),
    .A2(_25339_),
    .ZN(_25340_)
  );
  AND2_X1 _33472_ (
    .A1(_22147_),
    .A2(_25340_),
    .ZN(_25341_)
  );
  INV_X1 _33473_ (
    .A(_25341_),
    .ZN(_25342_)
  );
  AND2_X1 _33474_ (
    .A1(_21768_),
    .A2(_00008_[2]),
    .ZN(_25343_)
  );
  INV_X1 _33475_ (
    .A(_25343_),
    .ZN(_25344_)
  );
  AND2_X1 _33476_ (
    .A1(_21469_),
    .A2(_22149_),
    .ZN(_25345_)
  );
  INV_X1 _33477_ (
    .A(_25345_),
    .ZN(_25346_)
  );
  AND2_X1 _33478_ (
    .A1(_00008_[0]),
    .A2(_25346_),
    .ZN(_25347_)
  );
  AND2_X1 _33479_ (
    .A1(_25344_),
    .A2(_25347_),
    .ZN(_25348_)
  );
  INV_X1 _33480_ (
    .A(_25348_),
    .ZN(_25349_)
  );
  AND2_X1 _33481_ (
    .A1(_25342_),
    .A2(_25349_),
    .ZN(_25350_)
  );
  AND2_X1 _33482_ (
    .A1(_22148_),
    .A2(_25350_),
    .ZN(_25351_)
  );
  INV_X1 _33483_ (
    .A(_25351_),
    .ZN(_25352_)
  );
  AND2_X1 _33484_ (
    .A1(_21602_),
    .A2(_22149_),
    .ZN(_25353_)
  );
  INV_X1 _33485_ (
    .A(_25353_),
    .ZN(_25354_)
  );
  AND2_X1 _33486_ (
    .A1(_21422_),
    .A2(_00008_[2]),
    .ZN(_25355_)
  );
  INV_X1 _33487_ (
    .A(_25355_),
    .ZN(_25356_)
  );
  AND2_X1 _33488_ (
    .A1(_25354_),
    .A2(_25356_),
    .ZN(_25357_)
  );
  AND2_X1 _33489_ (
    .A1(_22147_),
    .A2(_25357_),
    .ZN(_25358_)
  );
  INV_X1 _33490_ (
    .A(_25358_),
    .ZN(_25359_)
  );
  AND2_X1 _33491_ (
    .A1(_21381_),
    .A2(_00008_[2]),
    .ZN(_25360_)
  );
  INV_X1 _33492_ (
    .A(_25360_),
    .ZN(_25361_)
  );
  AND2_X1 _33493_ (
    .A1(_21627_),
    .A2(_22149_),
    .ZN(_25362_)
  );
  INV_X1 _33494_ (
    .A(_25362_),
    .ZN(_25363_)
  );
  AND2_X1 _33495_ (
    .A1(_00008_[0]),
    .A2(_25363_),
    .ZN(_25364_)
  );
  AND2_X1 _33496_ (
    .A1(_25361_),
    .A2(_25364_),
    .ZN(_25365_)
  );
  INV_X1 _33497_ (
    .A(_25365_),
    .ZN(_25366_)
  );
  AND2_X1 _33498_ (
    .A1(_25359_),
    .A2(_25366_),
    .ZN(_25367_)
  );
  AND2_X1 _33499_ (
    .A1(_00008_[1]),
    .A2(_25367_),
    .ZN(_25368_)
  );
  INV_X1 _33500_ (
    .A(_25368_),
    .ZN(_25369_)
  );
  AND2_X1 _33501_ (
    .A1(_21791_),
    .A2(_00008_[2]),
    .ZN(_25370_)
  );
  INV_X1 _33502_ (
    .A(_25370_),
    .ZN(_25371_)
  );
  AND2_X1 _33503_ (
    .A1(_21499_),
    .A2(_22149_),
    .ZN(_25372_)
  );
  INV_X1 _33504_ (
    .A(_25372_),
    .ZN(_25373_)
  );
  AND2_X1 _33505_ (
    .A1(_00008_[0]),
    .A2(_25373_),
    .ZN(_25374_)
  );
  AND2_X1 _33506_ (
    .A1(_25371_),
    .A2(_25374_),
    .ZN(_25375_)
  );
  INV_X1 _33507_ (
    .A(_25375_),
    .ZN(_25376_)
  );
  AND2_X1 _33508_ (
    .A1(_21552_),
    .A2(_22149_),
    .ZN(_25377_)
  );
  INV_X1 _33509_ (
    .A(_25377_),
    .ZN(_25378_)
  );
  AND2_X1 _33510_ (
    .A1(_21818_),
    .A2(_00008_[2]),
    .ZN(_25379_)
  );
  INV_X1 _33511_ (
    .A(_25379_),
    .ZN(_25380_)
  );
  AND2_X1 _33512_ (
    .A1(_25378_),
    .A2(_25380_),
    .ZN(_25381_)
  );
  AND2_X1 _33513_ (
    .A1(_22147_),
    .A2(_25381_),
    .ZN(_25382_)
  );
  INV_X1 _33514_ (
    .A(_25382_),
    .ZN(_25383_)
  );
  AND2_X1 _33515_ (
    .A1(_25376_),
    .A2(_25383_),
    .ZN(_25384_)
  );
  AND2_X1 _33516_ (
    .A1(_00008_[1]),
    .A2(_25384_),
    .ZN(_25385_)
  );
  INV_X1 _33517_ (
    .A(_25385_),
    .ZN(_25386_)
  );
  AND2_X1 _33518_ (
    .A1(_21744_),
    .A2(_00008_[2]),
    .ZN(_25387_)
  );
  INV_X1 _33519_ (
    .A(_25387_),
    .ZN(_25388_)
  );
  AND2_X1 _33520_ (
    .A1(_21524_),
    .A2(_22149_),
    .ZN(_25389_)
  );
  INV_X1 _33521_ (
    .A(_25389_),
    .ZN(_25390_)
  );
  AND2_X1 _33522_ (
    .A1(_00008_[0]),
    .A2(_25390_),
    .ZN(_25391_)
  );
  AND2_X1 _33523_ (
    .A1(_25388_),
    .A2(_25391_),
    .ZN(_25392_)
  );
  INV_X1 _33524_ (
    .A(_25392_),
    .ZN(_25393_)
  );
  AND2_X1 _33525_ (
    .A1(_21965_),
    .A2(_22149_),
    .ZN(_25394_)
  );
  INV_X1 _33526_ (
    .A(_25394_),
    .ZN(_25395_)
  );
  AND2_X1 _33527_ (
    .A1(_21681_),
    .A2(_00008_[2]),
    .ZN(_25396_)
  );
  INV_X1 _33528_ (
    .A(_25396_),
    .ZN(_25397_)
  );
  AND2_X1 _33529_ (
    .A1(_25395_),
    .A2(_25397_),
    .ZN(_25398_)
  );
  AND2_X1 _33530_ (
    .A1(_22147_),
    .A2(_25398_),
    .ZN(_25399_)
  );
  INV_X1 _33531_ (
    .A(_25399_),
    .ZN(_25400_)
  );
  AND2_X1 _33532_ (
    .A1(_25393_),
    .A2(_25400_),
    .ZN(_25401_)
  );
  AND2_X1 _33533_ (
    .A1(_22148_),
    .A2(_25401_),
    .ZN(_25402_)
  );
  INV_X1 _33534_ (
    .A(_25402_),
    .ZN(_25403_)
  );
  AND2_X1 _33535_ (
    .A1(_25386_),
    .A2(_25403_),
    .ZN(_25404_)
  );
  AND2_X1 _33536_ (
    .A1(_00008_[4]),
    .A2(_25369_),
    .ZN(_25405_)
  );
  AND2_X1 _33537_ (
    .A1(_25352_),
    .A2(_25405_),
    .ZN(_25406_)
  );
  INV_X1 _33538_ (
    .A(_25406_),
    .ZN(_25407_)
  );
  AND2_X1 _33539_ (
    .A1(_22151_),
    .A2(_25404_),
    .ZN(_25408_)
  );
  INV_X1 _33540_ (
    .A(_25408_),
    .ZN(_25409_)
  );
  AND2_X1 _33541_ (
    .A1(_25407_),
    .A2(_25409_),
    .ZN(_25410_)
  );
  AND2_X1 _33542_ (
    .A1(_22150_),
    .A2(_25410_),
    .ZN(_25411_)
  );
  INV_X1 _33543_ (
    .A(_25411_),
    .ZN(_25412_)
  );
  AND2_X1 _33544_ (
    .A1(_22546_),
    .A2(_25412_),
    .ZN(_25413_)
  );
  AND2_X1 _33545_ (
    .A1(_25335_),
    .A2(_25413_),
    .ZN(_25414_)
  );
  INV_X1 _33546_ (
    .A(_25414_),
    .ZN(_25415_)
  );
  AND2_X1 _33547_ (
    .A1(_25255_),
    .A2(_25415_),
    .ZN(_25416_)
  );
  INV_X1 _33548_ (
    .A(_25416_),
    .ZN(_25417_)
  );
  AND2_X1 _33549_ (
    .A1(_22271_),
    .A2(_25417_),
    .ZN(_25418_)
  );
  INV_X1 _33550_ (
    .A(_25418_),
    .ZN(_25419_)
  );
  AND2_X1 _33551_ (
    .A1(reg_op1[14]),
    .A2(_22285_),
    .ZN(_25420_)
  );
  INV_X1 _33552_ (
    .A(_25420_),
    .ZN(_25421_)
  );
  AND2_X1 _33553_ (
    .A1(_24814_),
    .A2(_25421_),
    .ZN(_25422_)
  );
  AND2_X1 _33554_ (
    .A1(reg_op1[19]),
    .A2(_22290_),
    .ZN(_25423_)
  );
  INV_X1 _33555_ (
    .A(_25423_),
    .ZN(_25424_)
  );
  AND2_X1 _33556_ (
    .A1(_24811_),
    .A2(_25424_),
    .ZN(_25425_)
  );
  AND2_X1 _33557_ (
    .A1(_22572_),
    .A2(_25422_),
    .ZN(_25426_)
  );
  INV_X1 _33558_ (
    .A(_25426_),
    .ZN(_25427_)
  );
  AND2_X1 _33559_ (
    .A1(_22573_),
    .A2(_25425_),
    .ZN(_25428_)
  );
  INV_X1 _33560_ (
    .A(_25428_),
    .ZN(_25429_)
  );
  AND2_X1 _33561_ (
    .A1(_22295_),
    .A2(_25429_),
    .ZN(_25430_)
  );
  AND2_X1 _33562_ (
    .A1(_25427_),
    .A2(_25430_),
    .ZN(_25431_)
  );
  INV_X1 _33563_ (
    .A(_25431_),
    .ZN(_25432_)
  );
  AND2_X1 _33564_ (
    .A1(_22333_),
    .A2(_25419_),
    .ZN(_25433_)
  );
  AND2_X1 _33565_ (
    .A1(_25432_),
    .A2(_25433_),
    .ZN(_25434_)
  );
  AND2_X1 _33566_ (
    .A1(reg_op1[15]),
    .A2(decoded_imm[15]),
    .ZN(_25435_)
  );
  INV_X1 _33567_ (
    .A(_25435_),
    .ZN(_25436_)
  );
  AND2_X1 _33568_ (
    .A1(_21182_),
    .A2(_21994_),
    .ZN(_25437_)
  );
  INV_X1 _33569_ (
    .A(_25437_),
    .ZN(_25438_)
  );
  AND2_X1 _33570_ (
    .A1(_25436_),
    .A2(_25438_),
    .ZN(_25439_)
  );
  INV_X1 _33571_ (
    .A(_25439_),
    .ZN(_25440_)
  );
  AND2_X1 _33572_ (
    .A1(_25238_),
    .A2(_25244_),
    .ZN(_25441_)
  );
  INV_X1 _33573_ (
    .A(_25441_),
    .ZN(_25442_)
  );
  AND2_X1 _33574_ (
    .A1(_25439_),
    .A2(_25442_),
    .ZN(_25443_)
  );
  INV_X1 _33575_ (
    .A(_25443_),
    .ZN(_25444_)
  );
  AND2_X1 _33576_ (
    .A1(_25440_),
    .A2(_25441_),
    .ZN(_25445_)
  );
  INV_X1 _33577_ (
    .A(_25445_),
    .ZN(_25446_)
  );
  AND2_X1 _33578_ (
    .A1(_22559_),
    .A2(_25446_),
    .ZN(_25447_)
  );
  AND2_X1 _33579_ (
    .A1(_25444_),
    .A2(_25447_),
    .ZN(_25448_)
  );
  INV_X1 _33580_ (
    .A(_25448_),
    .ZN(_25449_)
  );
  AND2_X1 _33581_ (
    .A1(_25434_),
    .A2(_25449_),
    .ZN(_25450_)
  );
  INV_X1 _33582_ (
    .A(_25450_),
    .ZN(_25451_)
  );
  AND2_X1 _33583_ (
    .A1(_25253_),
    .A2(_25451_),
    .ZN(_00072_)
  );
  AND2_X1 _33584_ (
    .A1(_21183_),
    .A2(_22334_),
    .ZN(_25452_)
  );
  INV_X1 _33585_ (
    .A(_25452_),
    .ZN(_25453_)
  );
  AND2_X1 _33586_ (
    .A1(reg_pc[16]),
    .A2(_22335_),
    .ZN(_25454_)
  );
  INV_X1 _33587_ (
    .A(_25454_),
    .ZN(_25455_)
  );
  AND2_X1 _33588_ (
    .A1(_21792_),
    .A2(_00008_[2]),
    .ZN(_25456_)
  );
  INV_X1 _33589_ (
    .A(_25456_),
    .ZN(_25457_)
  );
  AND2_X1 _33590_ (
    .A1(_21500_),
    .A2(_22149_),
    .ZN(_25458_)
  );
  INV_X1 _33591_ (
    .A(_25458_),
    .ZN(_25459_)
  );
  AND2_X1 _33592_ (
    .A1(_00008_[0]),
    .A2(_25459_),
    .ZN(_25460_)
  );
  AND2_X1 _33593_ (
    .A1(_25457_),
    .A2(_25460_),
    .ZN(_25461_)
  );
  INV_X1 _33594_ (
    .A(_25461_),
    .ZN(_25462_)
  );
  AND2_X1 _33595_ (
    .A1(_21553_),
    .A2(_22149_),
    .ZN(_25463_)
  );
  INV_X1 _33596_ (
    .A(_25463_),
    .ZN(_25464_)
  );
  AND2_X1 _33597_ (
    .A1(_21819_),
    .A2(_00008_[2]),
    .ZN(_25465_)
  );
  INV_X1 _33598_ (
    .A(_25465_),
    .ZN(_25466_)
  );
  AND2_X1 _33599_ (
    .A1(_25464_),
    .A2(_25466_),
    .ZN(_25467_)
  );
  AND2_X1 _33600_ (
    .A1(_22147_),
    .A2(_25467_),
    .ZN(_25468_)
  );
  INV_X1 _33601_ (
    .A(_25468_),
    .ZN(_25469_)
  );
  AND2_X1 _33602_ (
    .A1(_25462_),
    .A2(_25469_),
    .ZN(_25470_)
  );
  AND2_X1 _33603_ (
    .A1(_21745_),
    .A2(_00008_[2]),
    .ZN(_25471_)
  );
  INV_X1 _33604_ (
    .A(_25471_),
    .ZN(_25472_)
  );
  AND2_X1 _33605_ (
    .A1(_21525_),
    .A2(_22149_),
    .ZN(_25473_)
  );
  INV_X1 _33606_ (
    .A(_25473_),
    .ZN(_25474_)
  );
  AND2_X1 _33607_ (
    .A1(_00008_[0]),
    .A2(_25472_),
    .ZN(_25475_)
  );
  AND2_X1 _33608_ (
    .A1(_25474_),
    .A2(_25475_),
    .ZN(_25476_)
  );
  INV_X1 _33609_ (
    .A(_25476_),
    .ZN(_25477_)
  );
  AND2_X1 _33610_ (
    .A1(_21966_),
    .A2(_22149_),
    .ZN(_25478_)
  );
  INV_X1 _33611_ (
    .A(_25478_),
    .ZN(_25479_)
  );
  AND2_X1 _33612_ (
    .A1(_21682_),
    .A2(_00008_[2]),
    .ZN(_25480_)
  );
  INV_X1 _33613_ (
    .A(_25480_),
    .ZN(_25481_)
  );
  AND2_X1 _33614_ (
    .A1(_25479_),
    .A2(_25481_),
    .ZN(_25482_)
  );
  AND2_X1 _33615_ (
    .A1(_22147_),
    .A2(_25482_),
    .ZN(_25483_)
  );
  INV_X1 _33616_ (
    .A(_25483_),
    .ZN(_25484_)
  );
  AND2_X1 _33617_ (
    .A1(_25477_),
    .A2(_25484_),
    .ZN(_25485_)
  );
  AND2_X1 _33618_ (
    .A1(_00008_[1]),
    .A2(_25470_),
    .ZN(_25486_)
  );
  INV_X1 _33619_ (
    .A(_25486_),
    .ZN(_25487_)
  );
  AND2_X1 _33620_ (
    .A1(_22148_),
    .A2(_25485_),
    .ZN(_25488_)
  );
  INV_X1 _33621_ (
    .A(_25488_),
    .ZN(_25489_)
  );
  AND2_X1 _33622_ (
    .A1(_22150_),
    .A2(_25489_),
    .ZN(_25490_)
  );
  AND2_X1 _33623_ (
    .A1(_25487_),
    .A2(_25490_),
    .ZN(_25491_)
  );
  INV_X1 _33624_ (
    .A(_25491_),
    .ZN(_25492_)
  );
  AND2_X1 _33625_ (
    .A1(\cpuregs[13] [16]),
    .A2(_00008_[0]),
    .ZN(_25493_)
  );
  INV_X1 _33626_ (
    .A(_25493_),
    .ZN(_25494_)
  );
  AND2_X1 _33627_ (
    .A1(\cpuregs[12] [16]),
    .A2(_22147_),
    .ZN(_25495_)
  );
  INV_X1 _33628_ (
    .A(_25495_),
    .ZN(_25496_)
  );
  AND2_X1 _33629_ (
    .A1(_00008_[2]),
    .A2(_25496_),
    .ZN(_25497_)
  );
  AND2_X1 _33630_ (
    .A1(_25494_),
    .A2(_25497_),
    .ZN(_25498_)
  );
  INV_X1 _33631_ (
    .A(_25498_),
    .ZN(_25499_)
  );
  AND2_X1 _33632_ (
    .A1(\cpuregs[9] [16]),
    .A2(_00008_[0]),
    .ZN(_25500_)
  );
  INV_X1 _33633_ (
    .A(_25500_),
    .ZN(_25501_)
  );
  AND2_X1 _33634_ (
    .A1(\cpuregs[8] [16]),
    .A2(_22147_),
    .ZN(_25502_)
  );
  INV_X1 _33635_ (
    .A(_25502_),
    .ZN(_25503_)
  );
  AND2_X1 _33636_ (
    .A1(_22149_),
    .A2(_25503_),
    .ZN(_25504_)
  );
  AND2_X1 _33637_ (
    .A1(_25501_),
    .A2(_25504_),
    .ZN(_25505_)
  );
  INV_X1 _33638_ (
    .A(_25505_),
    .ZN(_25506_)
  );
  AND2_X1 _33639_ (
    .A1(_22148_),
    .A2(_25506_),
    .ZN(_25507_)
  );
  AND2_X1 _33640_ (
    .A1(_25499_),
    .A2(_25507_),
    .ZN(_25508_)
  );
  INV_X1 _33641_ (
    .A(_25508_),
    .ZN(_25509_)
  );
  AND2_X1 _33642_ (
    .A1(\cpuregs[15] [16]),
    .A2(_00008_[0]),
    .ZN(_25510_)
  );
  INV_X1 _33643_ (
    .A(_25510_),
    .ZN(_25511_)
  );
  AND2_X1 _33644_ (
    .A1(\cpuregs[14] [16]),
    .A2(_22147_),
    .ZN(_25512_)
  );
  INV_X1 _33645_ (
    .A(_25512_),
    .ZN(_25513_)
  );
  AND2_X1 _33646_ (
    .A1(_00008_[2]),
    .A2(_25513_),
    .ZN(_25514_)
  );
  AND2_X1 _33647_ (
    .A1(_25511_),
    .A2(_25514_),
    .ZN(_25515_)
  );
  INV_X1 _33648_ (
    .A(_25515_),
    .ZN(_25516_)
  );
  AND2_X1 _33649_ (
    .A1(\cpuregs[11] [16]),
    .A2(_00008_[0]),
    .ZN(_25517_)
  );
  INV_X1 _33650_ (
    .A(_25517_),
    .ZN(_25518_)
  );
  AND2_X1 _33651_ (
    .A1(\cpuregs[10] [16]),
    .A2(_22147_),
    .ZN(_25519_)
  );
  INV_X1 _33652_ (
    .A(_25519_),
    .ZN(_25520_)
  );
  AND2_X1 _33653_ (
    .A1(_22149_),
    .A2(_25520_),
    .ZN(_25521_)
  );
  AND2_X1 _33654_ (
    .A1(_25518_),
    .A2(_25521_),
    .ZN(_25522_)
  );
  INV_X1 _33655_ (
    .A(_25522_),
    .ZN(_25523_)
  );
  AND2_X1 _33656_ (
    .A1(_00008_[1]),
    .A2(_25523_),
    .ZN(_25524_)
  );
  AND2_X1 _33657_ (
    .A1(_25516_),
    .A2(_25524_),
    .ZN(_25525_)
  );
  INV_X1 _33658_ (
    .A(_25525_),
    .ZN(_25526_)
  );
  AND2_X1 _33659_ (
    .A1(_25509_),
    .A2(_25526_),
    .ZN(_25527_)
  );
  INV_X1 _33660_ (
    .A(_25527_),
    .ZN(_25528_)
  );
  AND2_X1 _33661_ (
    .A1(_00008_[3]),
    .A2(_25528_),
    .ZN(_25529_)
  );
  INV_X1 _33662_ (
    .A(_25529_),
    .ZN(_25530_)
  );
  AND2_X1 _33663_ (
    .A1(_22151_),
    .A2(_25492_),
    .ZN(_25531_)
  );
  AND2_X1 _33664_ (
    .A1(_25530_),
    .A2(_25531_),
    .ZN(_25532_)
  );
  INV_X1 _33665_ (
    .A(_25532_),
    .ZN(_25533_)
  );
  AND2_X1 _33666_ (
    .A1(_21878_),
    .A2(_22149_),
    .ZN(_25534_)
  );
  INV_X1 _33667_ (
    .A(_25534_),
    .ZN(_25535_)
  );
  AND2_X1 _33668_ (
    .A1(_21858_),
    .A2(_00008_[2]),
    .ZN(_25536_)
  );
  INV_X1 _33669_ (
    .A(_25536_),
    .ZN(_25537_)
  );
  AND2_X1 _33670_ (
    .A1(_25535_),
    .A2(_25537_),
    .ZN(_25538_)
  );
  AND2_X1 _33671_ (
    .A1(_22147_),
    .A2(_25538_),
    .ZN(_25539_)
  );
  INV_X1 _33672_ (
    .A(_25539_),
    .ZN(_25540_)
  );
  AND2_X1 _33673_ (
    .A1(_21946_),
    .A2(_00008_[2]),
    .ZN(_25541_)
  );
  INV_X1 _33674_ (
    .A(_25541_),
    .ZN(_25542_)
  );
  AND2_X1 _33675_ (
    .A1(_21930_),
    .A2(_22149_),
    .ZN(_25543_)
  );
  INV_X1 _33676_ (
    .A(_25543_),
    .ZN(_25544_)
  );
  AND2_X1 _33677_ (
    .A1(_00008_[0]),
    .A2(_25544_),
    .ZN(_25545_)
  );
  AND2_X1 _33678_ (
    .A1(_25542_),
    .A2(_25545_),
    .ZN(_25546_)
  );
  INV_X1 _33679_ (
    .A(_25546_),
    .ZN(_25547_)
  );
  AND2_X1 _33680_ (
    .A1(_25540_),
    .A2(_25547_),
    .ZN(_25548_)
  );
  AND2_X1 _33681_ (
    .A1(_00008_[3]),
    .A2(_25548_),
    .ZN(_25549_)
  );
  INV_X1 _33682_ (
    .A(_25549_),
    .ZN(_25550_)
  );
  AND2_X1 _33683_ (
    .A1(\cpuregs[18] [16]),
    .A2(_22149_),
    .ZN(_25551_)
  );
  INV_X1 _33684_ (
    .A(_25551_),
    .ZN(_25552_)
  );
  AND2_X1 _33685_ (
    .A1(\cpuregs[22] [16]),
    .A2(_00008_[2]),
    .ZN(_25553_)
  );
  INV_X1 _33686_ (
    .A(_25553_),
    .ZN(_25554_)
  );
  AND2_X1 _33687_ (
    .A1(_22147_),
    .A2(_25554_),
    .ZN(_25555_)
  );
  AND2_X1 _33688_ (
    .A1(_25552_),
    .A2(_25555_),
    .ZN(_25556_)
  );
  INV_X1 _33689_ (
    .A(_25556_),
    .ZN(_25557_)
  );
  AND2_X1 _33690_ (
    .A1(\cpuregs[19] [16]),
    .A2(_22149_),
    .ZN(_25558_)
  );
  INV_X1 _33691_ (
    .A(_25558_),
    .ZN(_25559_)
  );
  AND2_X1 _33692_ (
    .A1(\cpuregs[23] [16]),
    .A2(_00008_[2]),
    .ZN(_25560_)
  );
  INV_X1 _33693_ (
    .A(_25560_),
    .ZN(_25561_)
  );
  AND2_X1 _33694_ (
    .A1(_00008_[0]),
    .A2(_25561_),
    .ZN(_25562_)
  );
  AND2_X1 _33695_ (
    .A1(_25559_),
    .A2(_25562_),
    .ZN(_25563_)
  );
  INV_X1 _33696_ (
    .A(_25563_),
    .ZN(_25564_)
  );
  AND2_X1 _33697_ (
    .A1(_25557_),
    .A2(_25564_),
    .ZN(_25565_)
  );
  INV_X1 _33698_ (
    .A(_25565_),
    .ZN(_25566_)
  );
  AND2_X1 _33699_ (
    .A1(_22150_),
    .A2(_25566_),
    .ZN(_25567_)
  );
  INV_X1 _33700_ (
    .A(_25567_),
    .ZN(_25568_)
  );
  AND2_X1 _33701_ (
    .A1(_25550_),
    .A2(_25568_),
    .ZN(_25569_)
  );
  AND2_X1 _33702_ (
    .A1(\cpuregs[16] [16]),
    .A2(_22149_),
    .ZN(_25570_)
  );
  INV_X1 _33703_ (
    .A(_25570_),
    .ZN(_25571_)
  );
  AND2_X1 _33704_ (
    .A1(\cpuregs[20] [16]),
    .A2(_00008_[2]),
    .ZN(_25572_)
  );
  INV_X1 _33705_ (
    .A(_25572_),
    .ZN(_25573_)
  );
  AND2_X1 _33706_ (
    .A1(_22147_),
    .A2(_25573_),
    .ZN(_25574_)
  );
  AND2_X1 _33707_ (
    .A1(_25571_),
    .A2(_25574_),
    .ZN(_25575_)
  );
  INV_X1 _33708_ (
    .A(_25575_),
    .ZN(_25576_)
  );
  AND2_X1 _33709_ (
    .A1(\cpuregs[17] [16]),
    .A2(_22149_),
    .ZN(_25577_)
  );
  INV_X1 _33710_ (
    .A(_25577_),
    .ZN(_25578_)
  );
  AND2_X1 _33711_ (
    .A1(\cpuregs[21] [16]),
    .A2(_00008_[2]),
    .ZN(_25579_)
  );
  INV_X1 _33712_ (
    .A(_25579_),
    .ZN(_25580_)
  );
  AND2_X1 _33713_ (
    .A1(_00008_[0]),
    .A2(_25580_),
    .ZN(_25581_)
  );
  AND2_X1 _33714_ (
    .A1(_25578_),
    .A2(_25581_),
    .ZN(_25582_)
  );
  INV_X1 _33715_ (
    .A(_25582_),
    .ZN(_25583_)
  );
  AND2_X1 _33716_ (
    .A1(_25576_),
    .A2(_25583_),
    .ZN(_25584_)
  );
  INV_X1 _33717_ (
    .A(_25584_),
    .ZN(_25585_)
  );
  AND2_X1 _33718_ (
    .A1(_22150_),
    .A2(_25585_),
    .ZN(_25586_)
  );
  INV_X1 _33719_ (
    .A(_25586_),
    .ZN(_25587_)
  );
  AND2_X1 _33720_ (
    .A1(_21898_),
    .A2(_00008_[2]),
    .ZN(_25588_)
  );
  INV_X1 _33721_ (
    .A(_25588_),
    .ZN(_25589_)
  );
  AND2_X1 _33722_ (
    .A1(_21842_),
    .A2(_22149_),
    .ZN(_25590_)
  );
  INV_X1 _33723_ (
    .A(_25590_),
    .ZN(_25591_)
  );
  AND2_X1 _33724_ (
    .A1(_00008_[0]),
    .A2(_25591_),
    .ZN(_25592_)
  );
  AND2_X1 _33725_ (
    .A1(_25589_),
    .A2(_25592_),
    .ZN(_25593_)
  );
  INV_X1 _33726_ (
    .A(_25593_),
    .ZN(_25594_)
  );
  AND2_X1 _33727_ (
    .A1(_21576_),
    .A2(_22149_),
    .ZN(_25595_)
  );
  INV_X1 _33728_ (
    .A(_25595_),
    .ZN(_25596_)
  );
  AND2_X1 _33729_ (
    .A1(_21914_),
    .A2(_00008_[2]),
    .ZN(_25597_)
  );
  INV_X1 _33730_ (
    .A(_25597_),
    .ZN(_25598_)
  );
  AND2_X1 _33731_ (
    .A1(_25596_),
    .A2(_25598_),
    .ZN(_25599_)
  );
  AND2_X1 _33732_ (
    .A1(_22147_),
    .A2(_25599_),
    .ZN(_25600_)
  );
  INV_X1 _33733_ (
    .A(_25600_),
    .ZN(_25601_)
  );
  AND2_X1 _33734_ (
    .A1(_25594_),
    .A2(_25601_),
    .ZN(_25602_)
  );
  AND2_X1 _33735_ (
    .A1(_00008_[3]),
    .A2(_25602_),
    .ZN(_25603_)
  );
  INV_X1 _33736_ (
    .A(_25603_),
    .ZN(_25604_)
  );
  AND2_X1 _33737_ (
    .A1(_25587_),
    .A2(_25604_),
    .ZN(_25605_)
  );
  AND2_X1 _33738_ (
    .A1(_00008_[1]),
    .A2(_25569_),
    .ZN(_25606_)
  );
  INV_X1 _33739_ (
    .A(_25606_),
    .ZN(_25607_)
  );
  AND2_X1 _33740_ (
    .A1(_22148_),
    .A2(_25605_),
    .ZN(_25608_)
  );
  INV_X1 _33741_ (
    .A(_25608_),
    .ZN(_25609_)
  );
  AND2_X1 _33742_ (
    .A1(_00008_[4]),
    .A2(_25607_),
    .ZN(_25610_)
  );
  AND2_X1 _33743_ (
    .A1(_25609_),
    .A2(_25610_),
    .ZN(_25611_)
  );
  INV_X1 _33744_ (
    .A(_25611_),
    .ZN(_25612_)
  );
  AND2_X1 _33745_ (
    .A1(_22546_),
    .A2(_25612_),
    .ZN(_25613_)
  );
  AND2_X1 _33746_ (
    .A1(_25533_),
    .A2(_25613_),
    .ZN(_25614_)
  );
  INV_X1 _33747_ (
    .A(_25614_),
    .ZN(_25615_)
  );
  AND2_X1 _33748_ (
    .A1(_25455_),
    .A2(_25615_),
    .ZN(_25616_)
  );
  INV_X1 _33749_ (
    .A(_25616_),
    .ZN(_25617_)
  );
  AND2_X1 _33750_ (
    .A1(_22271_),
    .A2(_25617_),
    .ZN(_25618_)
  );
  INV_X1 _33751_ (
    .A(_25618_),
    .ZN(_25619_)
  );
  AND2_X1 _33752_ (
    .A1(reg_op1[15]),
    .A2(_22285_),
    .ZN(_25620_)
  );
  INV_X1 _33753_ (
    .A(_25620_),
    .ZN(_25621_)
  );
  AND2_X1 _33754_ (
    .A1(_25017_),
    .A2(_25621_),
    .ZN(_25622_)
  );
  AND2_X1 _33755_ (
    .A1(reg_op1[20]),
    .A2(_22290_),
    .ZN(_25623_)
  );
  INV_X1 _33756_ (
    .A(_25623_),
    .ZN(_25624_)
  );
  AND2_X1 _33757_ (
    .A1(_25014_),
    .A2(_25624_),
    .ZN(_25625_)
  );
  AND2_X1 _33758_ (
    .A1(_22572_),
    .A2(_25622_),
    .ZN(_25626_)
  );
  INV_X1 _33759_ (
    .A(_25626_),
    .ZN(_25627_)
  );
  AND2_X1 _33760_ (
    .A1(_22573_),
    .A2(_25625_),
    .ZN(_25628_)
  );
  INV_X1 _33761_ (
    .A(_25628_),
    .ZN(_25629_)
  );
  AND2_X1 _33762_ (
    .A1(_22295_),
    .A2(_25629_),
    .ZN(_25630_)
  );
  AND2_X1 _33763_ (
    .A1(_25627_),
    .A2(_25630_),
    .ZN(_25631_)
  );
  INV_X1 _33764_ (
    .A(_25631_),
    .ZN(_25632_)
  );
  AND2_X1 _33765_ (
    .A1(_22333_),
    .A2(_25632_),
    .ZN(_25633_)
  );
  AND2_X1 _33766_ (
    .A1(_25619_),
    .A2(_25633_),
    .ZN(_25634_)
  );
  AND2_X1 _33767_ (
    .A1(_25436_),
    .A2(_25444_),
    .ZN(_25635_)
  );
  INV_X1 _33768_ (
    .A(_25635_),
    .ZN(_25636_)
  );
  AND2_X1 _33769_ (
    .A1(reg_op1[16]),
    .A2(decoded_imm[16]),
    .ZN(_25637_)
  );
  INV_X1 _33770_ (
    .A(_25637_),
    .ZN(_25638_)
  );
  AND2_X1 _33771_ (
    .A1(_21183_),
    .A2(_21993_),
    .ZN(_25639_)
  );
  INV_X1 _33772_ (
    .A(_25639_),
    .ZN(_25640_)
  );
  AND2_X1 _33773_ (
    .A1(_25638_),
    .A2(_25640_),
    .ZN(_25641_)
  );
  INV_X1 _33774_ (
    .A(_25641_),
    .ZN(_25642_)
  );
  AND2_X1 _33775_ (
    .A1(_25636_),
    .A2(_25641_),
    .ZN(_25643_)
  );
  INV_X1 _33776_ (
    .A(_25643_),
    .ZN(_25644_)
  );
  AND2_X1 _33777_ (
    .A1(_25635_),
    .A2(_25642_),
    .ZN(_25645_)
  );
  INV_X1 _33778_ (
    .A(_25645_),
    .ZN(_25646_)
  );
  AND2_X1 _33779_ (
    .A1(_22559_),
    .A2(_25646_),
    .ZN(_25647_)
  );
  AND2_X1 _33780_ (
    .A1(_25644_),
    .A2(_25647_),
    .ZN(_25648_)
  );
  INV_X1 _33781_ (
    .A(_25648_),
    .ZN(_25649_)
  );
  AND2_X1 _33782_ (
    .A1(_25634_),
    .A2(_25649_),
    .ZN(_25650_)
  );
  INV_X1 _33783_ (
    .A(_25650_),
    .ZN(_25651_)
  );
  AND2_X1 _33784_ (
    .A1(_25453_),
    .A2(_25651_),
    .ZN(_00073_)
  );
  AND2_X1 _33785_ (
    .A1(_21184_),
    .A2(_22334_),
    .ZN(_25652_)
  );
  INV_X1 _33786_ (
    .A(_25652_),
    .ZN(_25653_)
  );
  AND2_X1 _33787_ (
    .A1(reg_op1[17]),
    .A2(decoded_imm[17]),
    .ZN(_25654_)
  );
  INV_X1 _33788_ (
    .A(_25654_),
    .ZN(_25655_)
  );
  AND2_X1 _33789_ (
    .A1(_21184_),
    .A2(_21992_),
    .ZN(_25656_)
  );
  INV_X1 _33790_ (
    .A(_25656_),
    .ZN(_25657_)
  );
  AND2_X1 _33791_ (
    .A1(_25655_),
    .A2(_25657_),
    .ZN(_25658_)
  );
  INV_X1 _33792_ (
    .A(_25658_),
    .ZN(_25659_)
  );
  AND2_X1 _33793_ (
    .A1(_25638_),
    .A2(_25659_),
    .ZN(_25660_)
  );
  AND2_X1 _33794_ (
    .A1(_25644_),
    .A2(_25660_),
    .ZN(_25661_)
  );
  INV_X1 _33795_ (
    .A(_25661_),
    .ZN(_25662_)
  );
  AND2_X1 _33796_ (
    .A1(_25643_),
    .A2(_25658_),
    .ZN(_25663_)
  );
  INV_X1 _33797_ (
    .A(_25663_),
    .ZN(_25664_)
  );
  AND2_X1 _33798_ (
    .A1(_25637_),
    .A2(_25658_),
    .ZN(_25665_)
  );
  INV_X1 _33799_ (
    .A(_25665_),
    .ZN(_25666_)
  );
  AND2_X1 _33800_ (
    .A1(_22559_),
    .A2(_25666_),
    .ZN(_25667_)
  );
  AND2_X1 _33801_ (
    .A1(_25664_),
    .A2(_25667_),
    .ZN(_25668_)
  );
  AND2_X1 _33802_ (
    .A1(_25662_),
    .A2(_25668_),
    .ZN(_25669_)
  );
  INV_X1 _33803_ (
    .A(_25669_),
    .ZN(_25670_)
  );
  AND2_X1 _33804_ (
    .A1(reg_pc[17]),
    .A2(_22335_),
    .ZN(_25671_)
  );
  INV_X1 _33805_ (
    .A(_25671_),
    .ZN(_25672_)
  );
  AND2_X1 _33806_ (
    .A1(\cpuregs[12] [17]),
    .A2(_00008_[2]),
    .ZN(_25673_)
  );
  INV_X1 _33807_ (
    .A(_25673_),
    .ZN(_25674_)
  );
  AND2_X1 _33808_ (
    .A1(\cpuregs[8] [17]),
    .A2(_22149_),
    .ZN(_25675_)
  );
  INV_X1 _33809_ (
    .A(_25675_),
    .ZN(_25676_)
  );
  AND2_X1 _33810_ (
    .A1(_25674_),
    .A2(_25676_),
    .ZN(_25677_)
  );
  INV_X1 _33811_ (
    .A(_25677_),
    .ZN(_25678_)
  );
  AND2_X1 _33812_ (
    .A1(_22147_),
    .A2(_25678_),
    .ZN(_25679_)
  );
  INV_X1 _33813_ (
    .A(_25679_),
    .ZN(_25680_)
  );
  AND2_X1 _33814_ (
    .A1(_21643_),
    .A2(_00008_[2]),
    .ZN(_25681_)
  );
  INV_X1 _33815_ (
    .A(_25681_),
    .ZN(_25682_)
  );
  AND2_X1 _33816_ (
    .A1(_21721_),
    .A2(_22149_),
    .ZN(_25683_)
  );
  INV_X1 _33817_ (
    .A(_25683_),
    .ZN(_25684_)
  );
  AND2_X1 _33818_ (
    .A1(_00008_[0]),
    .A2(_25682_),
    .ZN(_25685_)
  );
  AND2_X1 _33819_ (
    .A1(_25684_),
    .A2(_25685_),
    .ZN(_25686_)
  );
  INV_X1 _33820_ (
    .A(_25686_),
    .ZN(_25687_)
  );
  AND2_X1 _33821_ (
    .A1(_22148_),
    .A2(_25687_),
    .ZN(_25688_)
  );
  AND2_X1 _33822_ (
    .A1(_25680_),
    .A2(_25688_),
    .ZN(_25689_)
  );
  INV_X1 _33823_ (
    .A(_25689_),
    .ZN(_25690_)
  );
  AND2_X1 _33824_ (
    .A1(_21707_),
    .A2(_22149_),
    .ZN(_25691_)
  );
  INV_X1 _33825_ (
    .A(_25691_),
    .ZN(_25692_)
  );
  AND2_X1 _33826_ (
    .A1(_21397_),
    .A2(_00008_[2]),
    .ZN(_25693_)
  );
  INV_X1 _33827_ (
    .A(_25693_),
    .ZN(_25694_)
  );
  AND2_X1 _33828_ (
    .A1(_25692_),
    .A2(_25694_),
    .ZN(_25695_)
  );
  AND2_X1 _33829_ (
    .A1(_22147_),
    .A2(_25695_),
    .ZN(_25696_)
  );
  INV_X1 _33830_ (
    .A(_25696_),
    .ZN(_25697_)
  );
  AND2_X1 _33831_ (
    .A1(_21404_),
    .A2(_00008_[2]),
    .ZN(_25698_)
  );
  INV_X1 _33832_ (
    .A(_25698_),
    .ZN(_25699_)
  );
  AND2_X1 _33833_ (
    .A1(_21586_),
    .A2(_22149_),
    .ZN(_25700_)
  );
  INV_X1 _33834_ (
    .A(_25700_),
    .ZN(_25701_)
  );
  AND2_X1 _33835_ (
    .A1(_00008_[0]),
    .A2(_25699_),
    .ZN(_25702_)
  );
  AND2_X1 _33836_ (
    .A1(_25701_),
    .A2(_25702_),
    .ZN(_25703_)
  );
  INV_X1 _33837_ (
    .A(_25703_),
    .ZN(_25704_)
  );
  AND2_X1 _33838_ (
    .A1(_25697_),
    .A2(_25704_),
    .ZN(_25705_)
  );
  AND2_X1 _33839_ (
    .A1(_00008_[1]),
    .A2(_25705_),
    .ZN(_25706_)
  );
  INV_X1 _33840_ (
    .A(_25706_),
    .ZN(_25707_)
  );
  AND2_X1 _33841_ (
    .A1(_25690_),
    .A2(_25707_),
    .ZN(_25708_)
  );
  AND2_X1 _33842_ (
    .A1(\cpuregs[27] [17]),
    .A2(_00008_[0]),
    .ZN(_25709_)
  );
  INV_X1 _33843_ (
    .A(_25709_),
    .ZN(_25710_)
  );
  AND2_X1 _33844_ (
    .A1(\cpuregs[26] [17]),
    .A2(_22147_),
    .ZN(_25711_)
  );
  INV_X1 _33845_ (
    .A(_25711_),
    .ZN(_25712_)
  );
  AND2_X1 _33846_ (
    .A1(_22149_),
    .A2(_25712_),
    .ZN(_25713_)
  );
  AND2_X1 _33847_ (
    .A1(_25710_),
    .A2(_25713_),
    .ZN(_25714_)
  );
  INV_X1 _33848_ (
    .A(_25714_),
    .ZN(_25715_)
  );
  AND2_X1 _33849_ (
    .A1(\cpuregs[31] [17]),
    .A2(_00008_[0]),
    .ZN(_25716_)
  );
  INV_X1 _33850_ (
    .A(_25716_),
    .ZN(_25717_)
  );
  AND2_X1 _33851_ (
    .A1(\cpuregs[30] [17]),
    .A2(_22147_),
    .ZN(_25718_)
  );
  INV_X1 _33852_ (
    .A(_25718_),
    .ZN(_25719_)
  );
  AND2_X1 _33853_ (
    .A1(_00008_[2]),
    .A2(_25719_),
    .ZN(_25720_)
  );
  AND2_X1 _33854_ (
    .A1(_25717_),
    .A2(_25720_),
    .ZN(_25721_)
  );
  INV_X1 _33855_ (
    .A(_25721_),
    .ZN(_25722_)
  );
  AND2_X1 _33856_ (
    .A1(_25715_),
    .A2(_25722_),
    .ZN(_25723_)
  );
  INV_X1 _33857_ (
    .A(_25723_),
    .ZN(_25724_)
  );
  AND2_X1 _33858_ (
    .A1(_00008_[1]),
    .A2(_25724_),
    .ZN(_25725_)
  );
  INV_X1 _33859_ (
    .A(_25725_),
    .ZN(_25726_)
  );
  AND2_X1 _33860_ (
    .A1(\cpuregs[25] [17]),
    .A2(_00008_[0]),
    .ZN(_25727_)
  );
  INV_X1 _33861_ (
    .A(_25727_),
    .ZN(_25728_)
  );
  AND2_X1 _33862_ (
    .A1(\cpuregs[24] [17]),
    .A2(_22147_),
    .ZN(_25729_)
  );
  INV_X1 _33863_ (
    .A(_25729_),
    .ZN(_25730_)
  );
  AND2_X1 _33864_ (
    .A1(_22149_),
    .A2(_25730_),
    .ZN(_25731_)
  );
  AND2_X1 _33865_ (
    .A1(_25728_),
    .A2(_25731_),
    .ZN(_25732_)
  );
  INV_X1 _33866_ (
    .A(_25732_),
    .ZN(_25733_)
  );
  AND2_X1 _33867_ (
    .A1(\cpuregs[29] [17]),
    .A2(_00008_[0]),
    .ZN(_25734_)
  );
  INV_X1 _33868_ (
    .A(_25734_),
    .ZN(_25735_)
  );
  AND2_X1 _33869_ (
    .A1(\cpuregs[28] [17]),
    .A2(_22147_),
    .ZN(_25736_)
  );
  INV_X1 _33870_ (
    .A(_25736_),
    .ZN(_25737_)
  );
  AND2_X1 _33871_ (
    .A1(_00008_[2]),
    .A2(_25737_),
    .ZN(_25738_)
  );
  AND2_X1 _33872_ (
    .A1(_25735_),
    .A2(_25738_),
    .ZN(_25739_)
  );
  INV_X1 _33873_ (
    .A(_25739_),
    .ZN(_25740_)
  );
  AND2_X1 _33874_ (
    .A1(_25733_),
    .A2(_25740_),
    .ZN(_25741_)
  );
  INV_X1 _33875_ (
    .A(_25741_),
    .ZN(_25742_)
  );
  AND2_X1 _33876_ (
    .A1(_22148_),
    .A2(_25742_),
    .ZN(_25743_)
  );
  INV_X1 _33877_ (
    .A(_25743_),
    .ZN(_25744_)
  );
  AND2_X1 _33878_ (
    .A1(_00008_[4]),
    .A2(_25726_),
    .ZN(_25745_)
  );
  AND2_X1 _33879_ (
    .A1(_25744_),
    .A2(_25745_),
    .ZN(_25746_)
  );
  INV_X1 _33880_ (
    .A(_25746_),
    .ZN(_25747_)
  );
  AND2_X1 _33881_ (
    .A1(_22151_),
    .A2(_25708_),
    .ZN(_25748_)
  );
  INV_X1 _33882_ (
    .A(_25748_),
    .ZN(_25749_)
  );
  AND2_X1 _33883_ (
    .A1(_25747_),
    .A2(_25749_),
    .ZN(_25750_)
  );
  AND2_X1 _33884_ (
    .A1(_00008_[3]),
    .A2(_25750_),
    .ZN(_25751_)
  );
  INV_X1 _33885_ (
    .A(_25751_),
    .ZN(_25752_)
  );
  AND2_X1 _33886_ (
    .A1(_21793_),
    .A2(_00008_[2]),
    .ZN(_25753_)
  );
  INV_X1 _33887_ (
    .A(_25753_),
    .ZN(_25754_)
  );
  AND2_X1 _33888_ (
    .A1(_21501_),
    .A2(_22149_),
    .ZN(_25755_)
  );
  INV_X1 _33889_ (
    .A(_25755_),
    .ZN(_25756_)
  );
  AND2_X1 _33890_ (
    .A1(_21554_),
    .A2(_22149_),
    .ZN(_25757_)
  );
  INV_X1 _33891_ (
    .A(_25757_),
    .ZN(_25758_)
  );
  AND2_X1 _33892_ (
    .A1(_21820_),
    .A2(_00008_[2]),
    .ZN(_25759_)
  );
  INV_X1 _33893_ (
    .A(_25759_),
    .ZN(_25760_)
  );
  AND2_X1 _33894_ (
    .A1(_25758_),
    .A2(_25760_),
    .ZN(_25761_)
  );
  AND2_X1 _33895_ (
    .A1(_00008_[0]),
    .A2(_25756_),
    .ZN(_25762_)
  );
  AND2_X1 _33896_ (
    .A1(_25754_),
    .A2(_25762_),
    .ZN(_25763_)
  );
  INV_X1 _33897_ (
    .A(_25763_),
    .ZN(_25764_)
  );
  AND2_X1 _33898_ (
    .A1(_22147_),
    .A2(_25761_),
    .ZN(_25765_)
  );
  INV_X1 _33899_ (
    .A(_25765_),
    .ZN(_25766_)
  );
  AND2_X1 _33900_ (
    .A1(_25764_),
    .A2(_25766_),
    .ZN(_25767_)
  );
  AND2_X1 _33901_ (
    .A1(_00008_[1]),
    .A2(_25767_),
    .ZN(_25768_)
  );
  INV_X1 _33902_ (
    .A(_25768_),
    .ZN(_25769_)
  );
  AND2_X1 _33903_ (
    .A1(_21526_),
    .A2(_22149_),
    .ZN(_25770_)
  );
  INV_X1 _33904_ (
    .A(_25770_),
    .ZN(_25771_)
  );
  AND2_X1 _33905_ (
    .A1(_21746_),
    .A2(_00008_[2]),
    .ZN(_25772_)
  );
  INV_X1 _33906_ (
    .A(_25772_),
    .ZN(_25773_)
  );
  AND2_X1 _33907_ (
    .A1(_21967_),
    .A2(_22149_),
    .ZN(_25774_)
  );
  INV_X1 _33908_ (
    .A(_25774_),
    .ZN(_25775_)
  );
  AND2_X1 _33909_ (
    .A1(_21683_),
    .A2(_00008_[2]),
    .ZN(_25776_)
  );
  INV_X1 _33910_ (
    .A(_25776_),
    .ZN(_25777_)
  );
  AND2_X1 _33911_ (
    .A1(_25775_),
    .A2(_25777_),
    .ZN(_25778_)
  );
  AND2_X1 _33912_ (
    .A1(_00008_[0]),
    .A2(_25771_),
    .ZN(_25779_)
  );
  AND2_X1 _33913_ (
    .A1(_25773_),
    .A2(_25779_),
    .ZN(_25780_)
  );
  INV_X1 _33914_ (
    .A(_25780_),
    .ZN(_25781_)
  );
  AND2_X1 _33915_ (
    .A1(_22147_),
    .A2(_25778_),
    .ZN(_25782_)
  );
  INV_X1 _33916_ (
    .A(_25782_),
    .ZN(_25783_)
  );
  AND2_X1 _33917_ (
    .A1(_25781_),
    .A2(_25783_),
    .ZN(_25784_)
  );
  AND2_X1 _33918_ (
    .A1(_22148_),
    .A2(_25784_),
    .ZN(_25785_)
  );
  INV_X1 _33919_ (
    .A(_25785_),
    .ZN(_25786_)
  );
  AND2_X1 _33920_ (
    .A1(_25769_),
    .A2(_25786_),
    .ZN(_25787_)
  );
  INV_X1 _33921_ (
    .A(_25787_),
    .ZN(_25788_)
  );
  AND2_X1 _33922_ (
    .A1(_22151_),
    .A2(_25788_),
    .ZN(_25789_)
  );
  INV_X1 _33923_ (
    .A(_25789_),
    .ZN(_25790_)
  );
  AND2_X1 _33924_ (
    .A1(\cpuregs[17] [17]),
    .A2(_22148_),
    .ZN(_25791_)
  );
  INV_X1 _33925_ (
    .A(_25791_),
    .ZN(_25792_)
  );
  AND2_X1 _33926_ (
    .A1(\cpuregs[19] [17]),
    .A2(_00008_[1]),
    .ZN(_25793_)
  );
  INV_X1 _33927_ (
    .A(_25793_),
    .ZN(_25794_)
  );
  AND2_X1 _33928_ (
    .A1(_22149_),
    .A2(_25794_),
    .ZN(_25795_)
  );
  AND2_X1 _33929_ (
    .A1(_25792_),
    .A2(_25795_),
    .ZN(_25796_)
  );
  INV_X1 _33930_ (
    .A(_25796_),
    .ZN(_25797_)
  );
  AND2_X1 _33931_ (
    .A1(\cpuregs[21] [17]),
    .A2(_22148_),
    .ZN(_25798_)
  );
  INV_X1 _33932_ (
    .A(_25798_),
    .ZN(_25799_)
  );
  AND2_X1 _33933_ (
    .A1(\cpuregs[23] [17]),
    .A2(_00008_[1]),
    .ZN(_25800_)
  );
  INV_X1 _33934_ (
    .A(_25800_),
    .ZN(_25801_)
  );
  AND2_X1 _33935_ (
    .A1(_00008_[2]),
    .A2(_25801_),
    .ZN(_25802_)
  );
  AND2_X1 _33936_ (
    .A1(_25799_),
    .A2(_25802_),
    .ZN(_25803_)
  );
  INV_X1 _33937_ (
    .A(_25803_),
    .ZN(_25804_)
  );
  AND2_X1 _33938_ (
    .A1(_25797_),
    .A2(_25804_),
    .ZN(_25805_)
  );
  INV_X1 _33939_ (
    .A(_25805_),
    .ZN(_25806_)
  );
  AND2_X1 _33940_ (
    .A1(_00008_[0]),
    .A2(_25806_),
    .ZN(_25807_)
  );
  INV_X1 _33941_ (
    .A(_25807_),
    .ZN(_25808_)
  );
  AND2_X1 _33942_ (
    .A1(\cpuregs[16] [17]),
    .A2(_22148_),
    .ZN(_25809_)
  );
  INV_X1 _33943_ (
    .A(_25809_),
    .ZN(_25810_)
  );
  AND2_X1 _33944_ (
    .A1(\cpuregs[18] [17]),
    .A2(_00008_[1]),
    .ZN(_25811_)
  );
  INV_X1 _33945_ (
    .A(_25811_),
    .ZN(_25812_)
  );
  AND2_X1 _33946_ (
    .A1(_22149_),
    .A2(_25812_),
    .ZN(_25813_)
  );
  AND2_X1 _33947_ (
    .A1(_25810_),
    .A2(_25813_),
    .ZN(_25814_)
  );
  INV_X1 _33948_ (
    .A(_25814_),
    .ZN(_25815_)
  );
  AND2_X1 _33949_ (
    .A1(\cpuregs[20] [17]),
    .A2(_22148_),
    .ZN(_25816_)
  );
  INV_X1 _33950_ (
    .A(_25816_),
    .ZN(_25817_)
  );
  AND2_X1 _33951_ (
    .A1(\cpuregs[22] [17]),
    .A2(_00008_[1]),
    .ZN(_25818_)
  );
  INV_X1 _33952_ (
    .A(_25818_),
    .ZN(_25819_)
  );
  AND2_X1 _33953_ (
    .A1(_00008_[2]),
    .A2(_25819_),
    .ZN(_25820_)
  );
  AND2_X1 _33954_ (
    .A1(_25817_),
    .A2(_25820_),
    .ZN(_25821_)
  );
  INV_X1 _33955_ (
    .A(_25821_),
    .ZN(_25822_)
  );
  AND2_X1 _33956_ (
    .A1(_25815_),
    .A2(_25822_),
    .ZN(_25823_)
  );
  INV_X1 _33957_ (
    .A(_25823_),
    .ZN(_25824_)
  );
  AND2_X1 _33958_ (
    .A1(_22147_),
    .A2(_25824_),
    .ZN(_25825_)
  );
  INV_X1 _33959_ (
    .A(_25825_),
    .ZN(_25826_)
  );
  AND2_X1 _33960_ (
    .A1(_25808_),
    .A2(_25826_),
    .ZN(_25827_)
  );
  INV_X1 _33961_ (
    .A(_25827_),
    .ZN(_25828_)
  );
  AND2_X1 _33962_ (
    .A1(_00008_[4]),
    .A2(_25828_),
    .ZN(_25829_)
  );
  INV_X1 _33963_ (
    .A(_25829_),
    .ZN(_25830_)
  );
  AND2_X1 _33964_ (
    .A1(_25790_),
    .A2(_25830_),
    .ZN(_25831_)
  );
  INV_X1 _33965_ (
    .A(_25831_),
    .ZN(_25832_)
  );
  AND2_X1 _33966_ (
    .A1(_22150_),
    .A2(_25832_),
    .ZN(_25833_)
  );
  INV_X1 _33967_ (
    .A(_25833_),
    .ZN(_25834_)
  );
  AND2_X1 _33968_ (
    .A1(_22546_),
    .A2(_25752_),
    .ZN(_25835_)
  );
  AND2_X1 _33969_ (
    .A1(_25834_),
    .A2(_25835_),
    .ZN(_25836_)
  );
  INV_X1 _33970_ (
    .A(_25836_),
    .ZN(_25837_)
  );
  AND2_X1 _33971_ (
    .A1(_25672_),
    .A2(_25837_),
    .ZN(_25838_)
  );
  INV_X1 _33972_ (
    .A(_25838_),
    .ZN(_25839_)
  );
  AND2_X1 _33973_ (
    .A1(_22271_),
    .A2(_25839_),
    .ZN(_25840_)
  );
  INV_X1 _33974_ (
    .A(_25840_),
    .ZN(_25841_)
  );
  AND2_X1 _33975_ (
    .A1(reg_op1[16]),
    .A2(_22285_),
    .ZN(_25842_)
  );
  INV_X1 _33976_ (
    .A(_25842_),
    .ZN(_25843_)
  );
  AND2_X1 _33977_ (
    .A1(_25224_),
    .A2(_25843_),
    .ZN(_25844_)
  );
  AND2_X1 _33978_ (
    .A1(reg_op1[21]),
    .A2(_22290_),
    .ZN(_25845_)
  );
  INV_X1 _33979_ (
    .A(_25845_),
    .ZN(_25846_)
  );
  AND2_X1 _33980_ (
    .A1(_25221_),
    .A2(_25846_),
    .ZN(_25847_)
  );
  AND2_X1 _33981_ (
    .A1(_22573_),
    .A2(_25847_),
    .ZN(_25848_)
  );
  INV_X1 _33982_ (
    .A(_25848_),
    .ZN(_25849_)
  );
  AND2_X1 _33983_ (
    .A1(_22572_),
    .A2(_25844_),
    .ZN(_25850_)
  );
  INV_X1 _33984_ (
    .A(_25850_),
    .ZN(_25851_)
  );
  AND2_X1 _33985_ (
    .A1(_22295_),
    .A2(_25851_),
    .ZN(_25852_)
  );
  AND2_X1 _33986_ (
    .A1(_25849_),
    .A2(_25852_),
    .ZN(_25853_)
  );
  INV_X1 _33987_ (
    .A(_25853_),
    .ZN(_25854_)
  );
  AND2_X1 _33988_ (
    .A1(_25841_),
    .A2(_25854_),
    .ZN(_25855_)
  );
  AND2_X1 _33989_ (
    .A1(_25670_),
    .A2(_25855_),
    .ZN(_25856_)
  );
  AND2_X1 _33990_ (
    .A1(_22333_),
    .A2(_25856_),
    .ZN(_25857_)
  );
  INV_X1 _33991_ (
    .A(_25857_),
    .ZN(_25858_)
  );
  AND2_X1 _33992_ (
    .A1(_25653_),
    .A2(_25858_),
    .ZN(_00074_)
  );
  AND2_X1 _33993_ (
    .A1(_21185_),
    .A2(_22334_),
    .ZN(_25859_)
  );
  INV_X1 _33994_ (
    .A(_25859_),
    .ZN(_25860_)
  );
  AND2_X1 _33995_ (
    .A1(reg_pc[18]),
    .A2(_22335_),
    .ZN(_25861_)
  );
  INV_X1 _33996_ (
    .A(_25861_),
    .ZN(_25862_)
  );
  AND2_X1 _33997_ (
    .A1(\cpuregs[22] [18]),
    .A2(_00008_[2]),
    .ZN(_25863_)
  );
  INV_X1 _33998_ (
    .A(_25863_),
    .ZN(_25864_)
  );
  AND2_X1 _33999_ (
    .A1(\cpuregs[18] [18]),
    .A2(_22149_),
    .ZN(_25865_)
  );
  INV_X1 _34000_ (
    .A(_25865_),
    .ZN(_25866_)
  );
  AND2_X1 _34001_ (
    .A1(_25864_),
    .A2(_25866_),
    .ZN(_25867_)
  );
  INV_X1 _34002_ (
    .A(_25867_),
    .ZN(_25868_)
  );
  AND2_X1 _34003_ (
    .A1(_22147_),
    .A2(_25868_),
    .ZN(_25869_)
  );
  INV_X1 _34004_ (
    .A(_25869_),
    .ZN(_25870_)
  );
  AND2_X1 _34005_ (
    .A1(\cpuregs[23] [18]),
    .A2(_00008_[2]),
    .ZN(_25871_)
  );
  INV_X1 _34006_ (
    .A(_25871_),
    .ZN(_25872_)
  );
  AND2_X1 _34007_ (
    .A1(\cpuregs[19] [18]),
    .A2(_22149_),
    .ZN(_25873_)
  );
  INV_X1 _34008_ (
    .A(_25873_),
    .ZN(_25874_)
  );
  AND2_X1 _34009_ (
    .A1(_25872_),
    .A2(_25874_),
    .ZN(_25875_)
  );
  INV_X1 _34010_ (
    .A(_25875_),
    .ZN(_25876_)
  );
  AND2_X1 _34011_ (
    .A1(_00008_[0]),
    .A2(_25876_),
    .ZN(_25877_)
  );
  INV_X1 _34012_ (
    .A(_25877_),
    .ZN(_25878_)
  );
  AND2_X1 _34013_ (
    .A1(_25870_),
    .A2(_25878_),
    .ZN(_25879_)
  );
  AND2_X1 _34014_ (
    .A1(_00008_[1]),
    .A2(_25879_),
    .ZN(_25880_)
  );
  INV_X1 _34015_ (
    .A(_25880_),
    .ZN(_25881_)
  );
  AND2_X1 _34016_ (
    .A1(\cpuregs[20] [18]),
    .A2(_00008_[2]),
    .ZN(_25882_)
  );
  INV_X1 _34017_ (
    .A(_25882_),
    .ZN(_25883_)
  );
  AND2_X1 _34018_ (
    .A1(\cpuregs[16] [18]),
    .A2(_22149_),
    .ZN(_25884_)
  );
  INV_X1 _34019_ (
    .A(_25884_),
    .ZN(_25885_)
  );
  AND2_X1 _34020_ (
    .A1(_25883_),
    .A2(_25885_),
    .ZN(_25886_)
  );
  INV_X1 _34021_ (
    .A(_25886_),
    .ZN(_25887_)
  );
  AND2_X1 _34022_ (
    .A1(_22147_),
    .A2(_25887_),
    .ZN(_25888_)
  );
  INV_X1 _34023_ (
    .A(_25888_),
    .ZN(_25889_)
  );
  AND2_X1 _34024_ (
    .A1(\cpuregs[21] [18]),
    .A2(_00008_[2]),
    .ZN(_25890_)
  );
  INV_X1 _34025_ (
    .A(_25890_),
    .ZN(_25891_)
  );
  AND2_X1 _34026_ (
    .A1(\cpuregs[17] [18]),
    .A2(_22149_),
    .ZN(_25892_)
  );
  INV_X1 _34027_ (
    .A(_25892_),
    .ZN(_25893_)
  );
  AND2_X1 _34028_ (
    .A1(_25891_),
    .A2(_25893_),
    .ZN(_25894_)
  );
  INV_X1 _34029_ (
    .A(_25894_),
    .ZN(_25895_)
  );
  AND2_X1 _34030_ (
    .A1(_00008_[0]),
    .A2(_25895_),
    .ZN(_25896_)
  );
  INV_X1 _34031_ (
    .A(_25896_),
    .ZN(_25897_)
  );
  AND2_X1 _34032_ (
    .A1(_25889_),
    .A2(_25897_),
    .ZN(_25898_)
  );
  AND2_X1 _34033_ (
    .A1(_22148_),
    .A2(_25898_),
    .ZN(_25899_)
  );
  INV_X1 _34034_ (
    .A(_25899_),
    .ZN(_25900_)
  );
  AND2_X1 _34035_ (
    .A1(\cpuregs[27] [18]),
    .A2(_00008_[0]),
    .ZN(_25901_)
  );
  INV_X1 _34036_ (
    .A(_25901_),
    .ZN(_25902_)
  );
  AND2_X1 _34037_ (
    .A1(\cpuregs[26] [18]),
    .A2(_22147_),
    .ZN(_25903_)
  );
  INV_X1 _34038_ (
    .A(_25903_),
    .ZN(_25904_)
  );
  AND2_X1 _34039_ (
    .A1(_22149_),
    .A2(_25904_),
    .ZN(_25905_)
  );
  AND2_X1 _34040_ (
    .A1(_25902_),
    .A2(_25905_),
    .ZN(_25906_)
  );
  INV_X1 _34041_ (
    .A(_25906_),
    .ZN(_25907_)
  );
  AND2_X1 _34042_ (
    .A1(\cpuregs[31] [18]),
    .A2(_00008_[0]),
    .ZN(_25908_)
  );
  INV_X1 _34043_ (
    .A(_25908_),
    .ZN(_25909_)
  );
  AND2_X1 _34044_ (
    .A1(\cpuregs[30] [18]),
    .A2(_22147_),
    .ZN(_25910_)
  );
  INV_X1 _34045_ (
    .A(_25910_),
    .ZN(_25911_)
  );
  AND2_X1 _34046_ (
    .A1(_00008_[2]),
    .A2(_25911_),
    .ZN(_25912_)
  );
  AND2_X1 _34047_ (
    .A1(_25909_),
    .A2(_25912_),
    .ZN(_25913_)
  );
  INV_X1 _34048_ (
    .A(_25913_),
    .ZN(_25914_)
  );
  AND2_X1 _34049_ (
    .A1(_25907_),
    .A2(_25914_),
    .ZN(_25915_)
  );
  INV_X1 _34050_ (
    .A(_25915_),
    .ZN(_25916_)
  );
  AND2_X1 _34051_ (
    .A1(_00008_[1]),
    .A2(_25916_),
    .ZN(_25917_)
  );
  INV_X1 _34052_ (
    .A(_25917_),
    .ZN(_25918_)
  );
  AND2_X1 _34053_ (
    .A1(\cpuregs[25] [18]),
    .A2(_00008_[0]),
    .ZN(_25919_)
  );
  INV_X1 _34054_ (
    .A(_25919_),
    .ZN(_25920_)
  );
  AND2_X1 _34055_ (
    .A1(\cpuregs[24] [18]),
    .A2(_22147_),
    .ZN(_25921_)
  );
  INV_X1 _34056_ (
    .A(_25921_),
    .ZN(_25922_)
  );
  AND2_X1 _34057_ (
    .A1(_22149_),
    .A2(_25922_),
    .ZN(_25923_)
  );
  AND2_X1 _34058_ (
    .A1(_25920_),
    .A2(_25923_),
    .ZN(_25924_)
  );
  INV_X1 _34059_ (
    .A(_25924_),
    .ZN(_25925_)
  );
  AND2_X1 _34060_ (
    .A1(\cpuregs[29] [18]),
    .A2(_00008_[0]),
    .ZN(_25926_)
  );
  INV_X1 _34061_ (
    .A(_25926_),
    .ZN(_25927_)
  );
  AND2_X1 _34062_ (
    .A1(\cpuregs[28] [18]),
    .A2(_22147_),
    .ZN(_25928_)
  );
  INV_X1 _34063_ (
    .A(_25928_),
    .ZN(_25929_)
  );
  AND2_X1 _34064_ (
    .A1(_00008_[2]),
    .A2(_25929_),
    .ZN(_25930_)
  );
  AND2_X1 _34065_ (
    .A1(_25927_),
    .A2(_25930_),
    .ZN(_25931_)
  );
  INV_X1 _34066_ (
    .A(_25931_),
    .ZN(_25932_)
  );
  AND2_X1 _34067_ (
    .A1(_25925_),
    .A2(_25932_),
    .ZN(_25933_)
  );
  INV_X1 _34068_ (
    .A(_25933_),
    .ZN(_25934_)
  );
  AND2_X1 _34069_ (
    .A1(_22148_),
    .A2(_25934_),
    .ZN(_25935_)
  );
  INV_X1 _34070_ (
    .A(_25935_),
    .ZN(_25936_)
  );
  AND2_X1 _34071_ (
    .A1(_00008_[3]),
    .A2(_25918_),
    .ZN(_25937_)
  );
  AND2_X1 _34072_ (
    .A1(_25936_),
    .A2(_25937_),
    .ZN(_25938_)
  );
  INV_X1 _34073_ (
    .A(_25938_),
    .ZN(_25939_)
  );
  AND2_X1 _34074_ (
    .A1(_22150_),
    .A2(_25900_),
    .ZN(_25940_)
  );
  AND2_X1 _34075_ (
    .A1(_25881_),
    .A2(_25940_),
    .ZN(_25941_)
  );
  INV_X1 _34076_ (
    .A(_25941_),
    .ZN(_25942_)
  );
  AND2_X1 _34077_ (
    .A1(_00008_[4]),
    .A2(_25942_),
    .ZN(_25943_)
  );
  AND2_X1 _34078_ (
    .A1(_25939_),
    .A2(_25943_),
    .ZN(_25944_)
  );
  INV_X1 _34079_ (
    .A(_25944_),
    .ZN(_25945_)
  );
  AND2_X1 _34080_ (
    .A1(\cpuregs[9] [18]),
    .A2(_22149_),
    .ZN(_25946_)
  );
  INV_X1 _34081_ (
    .A(_25946_),
    .ZN(_25947_)
  );
  AND2_X1 _34082_ (
    .A1(\cpuregs[13] [18]),
    .A2(_00008_[2]),
    .ZN(_25948_)
  );
  INV_X1 _34083_ (
    .A(_25948_),
    .ZN(_25949_)
  );
  AND2_X1 _34084_ (
    .A1(_22148_),
    .A2(_25949_),
    .ZN(_25950_)
  );
  AND2_X1 _34085_ (
    .A1(_25947_),
    .A2(_25950_),
    .ZN(_25951_)
  );
  INV_X1 _34086_ (
    .A(_25951_),
    .ZN(_25952_)
  );
  AND2_X1 _34087_ (
    .A1(\cpuregs[15] [18]),
    .A2(_00008_[2]),
    .ZN(_25953_)
  );
  INV_X1 _34088_ (
    .A(_25953_),
    .ZN(_25954_)
  );
  AND2_X1 _34089_ (
    .A1(\cpuregs[11] [18]),
    .A2(_22149_),
    .ZN(_25955_)
  );
  INV_X1 _34090_ (
    .A(_25955_),
    .ZN(_25956_)
  );
  AND2_X1 _34091_ (
    .A1(_00008_[1]),
    .A2(_25956_),
    .ZN(_25957_)
  );
  AND2_X1 _34092_ (
    .A1(_25954_),
    .A2(_25957_),
    .ZN(_25958_)
  );
  INV_X1 _34093_ (
    .A(_25958_),
    .ZN(_25959_)
  );
  AND2_X1 _34094_ (
    .A1(_25952_),
    .A2(_25959_),
    .ZN(_25960_)
  );
  INV_X1 _34095_ (
    .A(_25960_),
    .ZN(_25961_)
  );
  AND2_X1 _34096_ (
    .A1(_00008_[0]),
    .A2(_25961_),
    .ZN(_25962_)
  );
  INV_X1 _34097_ (
    .A(_25962_),
    .ZN(_25963_)
  );
  AND2_X1 _34098_ (
    .A1(\cpuregs[8] [18]),
    .A2(_22149_),
    .ZN(_25964_)
  );
  INV_X1 _34099_ (
    .A(_25964_),
    .ZN(_25965_)
  );
  AND2_X1 _34100_ (
    .A1(\cpuregs[12] [18]),
    .A2(_00008_[2]),
    .ZN(_25966_)
  );
  INV_X1 _34101_ (
    .A(_25966_),
    .ZN(_25967_)
  );
  AND2_X1 _34102_ (
    .A1(_22148_),
    .A2(_25967_),
    .ZN(_25968_)
  );
  AND2_X1 _34103_ (
    .A1(_25965_),
    .A2(_25968_),
    .ZN(_25969_)
  );
  INV_X1 _34104_ (
    .A(_25969_),
    .ZN(_25970_)
  );
  AND2_X1 _34105_ (
    .A1(\cpuregs[10] [18]),
    .A2(_22149_),
    .ZN(_25971_)
  );
  INV_X1 _34106_ (
    .A(_25971_),
    .ZN(_25972_)
  );
  AND2_X1 _34107_ (
    .A1(\cpuregs[14] [18]),
    .A2(_00008_[2]),
    .ZN(_25973_)
  );
  INV_X1 _34108_ (
    .A(_25973_),
    .ZN(_25974_)
  );
  AND2_X1 _34109_ (
    .A1(_00008_[1]),
    .A2(_25974_),
    .ZN(_25975_)
  );
  AND2_X1 _34110_ (
    .A1(_25972_),
    .A2(_25975_),
    .ZN(_25976_)
  );
  INV_X1 _34111_ (
    .A(_25976_),
    .ZN(_25977_)
  );
  AND2_X1 _34112_ (
    .A1(_25970_),
    .A2(_25977_),
    .ZN(_25978_)
  );
  INV_X1 _34113_ (
    .A(_25978_),
    .ZN(_25979_)
  );
  AND2_X1 _34114_ (
    .A1(_22147_),
    .A2(_25979_),
    .ZN(_25980_)
  );
  INV_X1 _34115_ (
    .A(_25980_),
    .ZN(_25981_)
  );
  AND2_X1 _34116_ (
    .A1(_25963_),
    .A2(_25981_),
    .ZN(_25982_)
  );
  INV_X1 _34117_ (
    .A(_25982_),
    .ZN(_25983_)
  );
  AND2_X1 _34118_ (
    .A1(_00008_[3]),
    .A2(_25983_),
    .ZN(_25984_)
  );
  INV_X1 _34119_ (
    .A(_25984_),
    .ZN(_25985_)
  );
  AND2_X1 _34120_ (
    .A1(_21747_),
    .A2(_00008_[2]),
    .ZN(_25986_)
  );
  INV_X1 _34121_ (
    .A(_25986_),
    .ZN(_25987_)
  );
  AND2_X1 _34122_ (
    .A1(_21527_),
    .A2(_22149_),
    .ZN(_25988_)
  );
  INV_X1 _34123_ (
    .A(_25988_),
    .ZN(_25989_)
  );
  AND2_X1 _34124_ (
    .A1(_00008_[0]),
    .A2(_25989_),
    .ZN(_25990_)
  );
  AND2_X1 _34125_ (
    .A1(_25987_),
    .A2(_25990_),
    .ZN(_25991_)
  );
  INV_X1 _34126_ (
    .A(_25991_),
    .ZN(_25992_)
  );
  AND2_X1 _34127_ (
    .A1(_21968_),
    .A2(_22149_),
    .ZN(_25993_)
  );
  INV_X1 _34128_ (
    .A(_25993_),
    .ZN(_25994_)
  );
  AND2_X1 _34129_ (
    .A1(_21684_),
    .A2(_00008_[2]),
    .ZN(_25995_)
  );
  INV_X1 _34130_ (
    .A(_25995_),
    .ZN(_25996_)
  );
  AND2_X1 _34131_ (
    .A1(_25994_),
    .A2(_25996_),
    .ZN(_25997_)
  );
  AND2_X1 _34132_ (
    .A1(_22147_),
    .A2(_25997_),
    .ZN(_25998_)
  );
  INV_X1 _34133_ (
    .A(_25998_),
    .ZN(_25999_)
  );
  AND2_X1 _34134_ (
    .A1(_25992_),
    .A2(_25999_),
    .ZN(_26000_)
  );
  AND2_X1 _34135_ (
    .A1(_22148_),
    .A2(_26000_),
    .ZN(_26001_)
  );
  INV_X1 _34136_ (
    .A(_26001_),
    .ZN(_26002_)
  );
  AND2_X1 _34137_ (
    .A1(_21794_),
    .A2(_00008_[2]),
    .ZN(_26003_)
  );
  INV_X1 _34138_ (
    .A(_26003_),
    .ZN(_26004_)
  );
  AND2_X1 _34139_ (
    .A1(_21502_),
    .A2(_22149_),
    .ZN(_26005_)
  );
  INV_X1 _34140_ (
    .A(_26005_),
    .ZN(_26006_)
  );
  AND2_X1 _34141_ (
    .A1(_00008_[0]),
    .A2(_26006_),
    .ZN(_26007_)
  );
  AND2_X1 _34142_ (
    .A1(_26004_),
    .A2(_26007_),
    .ZN(_26008_)
  );
  INV_X1 _34143_ (
    .A(_26008_),
    .ZN(_26009_)
  );
  AND2_X1 _34144_ (
    .A1(_21555_),
    .A2(_22149_),
    .ZN(_26010_)
  );
  INV_X1 _34145_ (
    .A(_26010_),
    .ZN(_26011_)
  );
  AND2_X1 _34146_ (
    .A1(_21821_),
    .A2(_00008_[2]),
    .ZN(_26012_)
  );
  INV_X1 _34147_ (
    .A(_26012_),
    .ZN(_26013_)
  );
  AND2_X1 _34148_ (
    .A1(_26011_),
    .A2(_26013_),
    .ZN(_26014_)
  );
  AND2_X1 _34149_ (
    .A1(_22147_),
    .A2(_26014_),
    .ZN(_26015_)
  );
  INV_X1 _34150_ (
    .A(_26015_),
    .ZN(_26016_)
  );
  AND2_X1 _34151_ (
    .A1(_26009_),
    .A2(_26016_),
    .ZN(_26017_)
  );
  AND2_X1 _34152_ (
    .A1(_00008_[1]),
    .A2(_26017_),
    .ZN(_26018_)
  );
  INV_X1 _34153_ (
    .A(_26018_),
    .ZN(_26019_)
  );
  AND2_X1 _34154_ (
    .A1(_26002_),
    .A2(_26019_),
    .ZN(_26020_)
  );
  INV_X1 _34155_ (
    .A(_26020_),
    .ZN(_26021_)
  );
  AND2_X1 _34156_ (
    .A1(_22150_),
    .A2(_26021_),
    .ZN(_26022_)
  );
  INV_X1 _34157_ (
    .A(_26022_),
    .ZN(_26023_)
  );
  AND2_X1 _34158_ (
    .A1(_25985_),
    .A2(_26023_),
    .ZN(_26024_)
  );
  INV_X1 _34159_ (
    .A(_26024_),
    .ZN(_26025_)
  );
  AND2_X1 _34160_ (
    .A1(_22151_),
    .A2(_26025_),
    .ZN(_26026_)
  );
  INV_X1 _34161_ (
    .A(_26026_),
    .ZN(_26027_)
  );
  AND2_X1 _34162_ (
    .A1(_22546_),
    .A2(_25945_),
    .ZN(_26028_)
  );
  AND2_X1 _34163_ (
    .A1(_26027_),
    .A2(_26028_),
    .ZN(_26029_)
  );
  INV_X1 _34164_ (
    .A(_26029_),
    .ZN(_26030_)
  );
  AND2_X1 _34165_ (
    .A1(_25862_),
    .A2(_26030_),
    .ZN(_26031_)
  );
  INV_X1 _34166_ (
    .A(_26031_),
    .ZN(_26032_)
  );
  AND2_X1 _34167_ (
    .A1(_22271_),
    .A2(_26032_),
    .ZN(_26033_)
  );
  INV_X1 _34168_ (
    .A(_26033_),
    .ZN(_26034_)
  );
  AND2_X1 _34169_ (
    .A1(reg_op1[17]),
    .A2(_22285_),
    .ZN(_26035_)
  );
  INV_X1 _34170_ (
    .A(_26035_),
    .ZN(_26036_)
  );
  AND2_X1 _34171_ (
    .A1(_25424_),
    .A2(_26036_),
    .ZN(_26037_)
  );
  AND2_X1 _34172_ (
    .A1(reg_op1[22]),
    .A2(_22290_),
    .ZN(_26038_)
  );
  INV_X1 _34173_ (
    .A(_26038_),
    .ZN(_26039_)
  );
  AND2_X1 _34174_ (
    .A1(_25421_),
    .A2(_26039_),
    .ZN(_26040_)
  );
  AND2_X1 _34175_ (
    .A1(_22572_),
    .A2(_26037_),
    .ZN(_26041_)
  );
  INV_X1 _34176_ (
    .A(_26041_),
    .ZN(_26042_)
  );
  AND2_X1 _34177_ (
    .A1(_22573_),
    .A2(_26040_),
    .ZN(_26043_)
  );
  INV_X1 _34178_ (
    .A(_26043_),
    .ZN(_26044_)
  );
  AND2_X1 _34179_ (
    .A1(_22295_),
    .A2(_26044_),
    .ZN(_26045_)
  );
  AND2_X1 _34180_ (
    .A1(_26042_),
    .A2(_26045_),
    .ZN(_26046_)
  );
  INV_X1 _34181_ (
    .A(_26046_),
    .ZN(_26047_)
  );
  AND2_X1 _34182_ (
    .A1(_22333_),
    .A2(_26047_),
    .ZN(_26048_)
  );
  AND2_X1 _34183_ (
    .A1(_26034_),
    .A2(_26048_),
    .ZN(_26049_)
  );
  AND2_X1 _34184_ (
    .A1(_25655_),
    .A2(_25666_),
    .ZN(_26050_)
  );
  AND2_X1 _34185_ (
    .A1(_25664_),
    .A2(_26050_),
    .ZN(_26051_)
  );
  INV_X1 _34186_ (
    .A(_26051_),
    .ZN(_26052_)
  );
  AND2_X1 _34187_ (
    .A1(reg_op1[18]),
    .A2(decoded_imm[18]),
    .ZN(_26053_)
  );
  INV_X1 _34188_ (
    .A(_26053_),
    .ZN(_26054_)
  );
  AND2_X1 _34189_ (
    .A1(_21185_),
    .A2(_21991_),
    .ZN(_26055_)
  );
  INV_X1 _34190_ (
    .A(_26055_),
    .ZN(_26056_)
  );
  AND2_X1 _34191_ (
    .A1(_26054_),
    .A2(_26056_),
    .ZN(_26057_)
  );
  INV_X1 _34192_ (
    .A(_26057_),
    .ZN(_26058_)
  );
  AND2_X1 _34193_ (
    .A1(_26052_),
    .A2(_26057_),
    .ZN(_26059_)
  );
  INV_X1 _34194_ (
    .A(_26059_),
    .ZN(_26060_)
  );
  AND2_X1 _34195_ (
    .A1(_26051_),
    .A2(_26058_),
    .ZN(_26061_)
  );
  INV_X1 _34196_ (
    .A(_26061_),
    .ZN(_26062_)
  );
  AND2_X1 _34197_ (
    .A1(_22559_),
    .A2(_26062_),
    .ZN(_26063_)
  );
  AND2_X1 _34198_ (
    .A1(_26060_),
    .A2(_26063_),
    .ZN(_26064_)
  );
  INV_X1 _34199_ (
    .A(_26064_),
    .ZN(_26065_)
  );
  AND2_X1 _34200_ (
    .A1(_26049_),
    .A2(_26065_),
    .ZN(_26066_)
  );
  INV_X1 _34201_ (
    .A(_26066_),
    .ZN(_26067_)
  );
  AND2_X1 _34202_ (
    .A1(_25860_),
    .A2(_26067_),
    .ZN(_00075_)
  );
  AND2_X1 _34203_ (
    .A1(_21186_),
    .A2(_22334_),
    .ZN(_26068_)
  );
  INV_X1 _34204_ (
    .A(_26068_),
    .ZN(_26069_)
  );
  AND2_X1 _34205_ (
    .A1(reg_pc[19]),
    .A2(_22335_),
    .ZN(_26070_)
  );
  INV_X1 _34206_ (
    .A(_26070_),
    .ZN(_26071_)
  );
  AND2_X1 _34207_ (
    .A1(_21450_),
    .A2(_22149_),
    .ZN(_26072_)
  );
  INV_X1 _34208_ (
    .A(_26072_),
    .ZN(_26073_)
  );
  AND2_X1 _34209_ (
    .A1(_21661_),
    .A2(_00008_[2]),
    .ZN(_26074_)
  );
  INV_X1 _34210_ (
    .A(_26074_),
    .ZN(_26075_)
  );
  AND2_X1 _34211_ (
    .A1(_26073_),
    .A2(_26075_),
    .ZN(_26076_)
  );
  AND2_X1 _34212_ (
    .A1(_22147_),
    .A2(_26076_),
    .ZN(_26077_)
  );
  INV_X1 _34213_ (
    .A(_26077_),
    .ZN(_26078_)
  );
  AND2_X1 _34214_ (
    .A1(_21771_),
    .A2(_00008_[2]),
    .ZN(_26079_)
  );
  INV_X1 _34215_ (
    .A(_26079_),
    .ZN(_26080_)
  );
  AND2_X1 _34216_ (
    .A1(_21472_),
    .A2(_22149_),
    .ZN(_26081_)
  );
  INV_X1 _34217_ (
    .A(_26081_),
    .ZN(_26082_)
  );
  AND2_X1 _34218_ (
    .A1(_00008_[0]),
    .A2(_26080_),
    .ZN(_26083_)
  );
  AND2_X1 _34219_ (
    .A1(_26082_),
    .A2(_26083_),
    .ZN(_26084_)
  );
  INV_X1 _34220_ (
    .A(_26084_),
    .ZN(_26085_)
  );
  AND2_X1 _34221_ (
    .A1(_26078_),
    .A2(_26085_),
    .ZN(_26086_)
  );
  AND2_X1 _34222_ (
    .A1(_22148_),
    .A2(_26086_),
    .ZN(_26087_)
  );
  INV_X1 _34223_ (
    .A(_26087_),
    .ZN(_26088_)
  );
  AND2_X1 _34224_ (
    .A1(_21605_),
    .A2(_22149_),
    .ZN(_26089_)
  );
  INV_X1 _34225_ (
    .A(_26089_),
    .ZN(_26090_)
  );
  AND2_X1 _34226_ (
    .A1(_21425_),
    .A2(_00008_[2]),
    .ZN(_26091_)
  );
  INV_X1 _34227_ (
    .A(_26091_),
    .ZN(_26092_)
  );
  AND2_X1 _34228_ (
    .A1(_26090_),
    .A2(_26092_),
    .ZN(_26093_)
  );
  AND2_X1 _34229_ (
    .A1(_22147_),
    .A2(_26093_),
    .ZN(_26094_)
  );
  INV_X1 _34230_ (
    .A(_26094_),
    .ZN(_26095_)
  );
  AND2_X1 _34231_ (
    .A1(_21384_),
    .A2(_00008_[2]),
    .ZN(_26096_)
  );
  INV_X1 _34232_ (
    .A(_26096_),
    .ZN(_26097_)
  );
  AND2_X1 _34233_ (
    .A1(_21630_),
    .A2(_22149_),
    .ZN(_26098_)
  );
  INV_X1 _34234_ (
    .A(_26098_),
    .ZN(_26099_)
  );
  AND2_X1 _34235_ (
    .A1(_00008_[0]),
    .A2(_26099_),
    .ZN(_26100_)
  );
  AND2_X1 _34236_ (
    .A1(_26097_),
    .A2(_26100_),
    .ZN(_26101_)
  );
  INV_X1 _34237_ (
    .A(_26101_),
    .ZN(_26102_)
  );
  AND2_X1 _34238_ (
    .A1(_26095_),
    .A2(_26102_),
    .ZN(_26103_)
  );
  AND2_X1 _34239_ (
    .A1(_00008_[1]),
    .A2(_26103_),
    .ZN(_26104_)
  );
  INV_X1 _34240_ (
    .A(_26104_),
    .ZN(_26105_)
  );
  AND2_X1 _34241_ (
    .A1(_26088_),
    .A2(_26105_),
    .ZN(_26106_)
  );
  AND2_X1 _34242_ (
    .A1(_21880_),
    .A2(_22149_),
    .ZN(_26107_)
  );
  INV_X1 _34243_ (
    .A(_26107_),
    .ZN(_26108_)
  );
  AND2_X1 _34244_ (
    .A1(_21859_),
    .A2(_00008_[2]),
    .ZN(_26109_)
  );
  INV_X1 _34245_ (
    .A(_26109_),
    .ZN(_26110_)
  );
  AND2_X1 _34246_ (
    .A1(_26108_),
    .A2(_26110_),
    .ZN(_26111_)
  );
  AND2_X1 _34247_ (
    .A1(_22147_),
    .A2(_26111_),
    .ZN(_26112_)
  );
  INV_X1 _34248_ (
    .A(_26112_),
    .ZN(_26113_)
  );
  AND2_X1 _34249_ (
    .A1(_21947_),
    .A2(_00008_[2]),
    .ZN(_26114_)
  );
  INV_X1 _34250_ (
    .A(_26114_),
    .ZN(_26115_)
  );
  AND2_X1 _34251_ (
    .A1(_21931_),
    .A2(_22149_),
    .ZN(_26116_)
  );
  INV_X1 _34252_ (
    .A(_26116_),
    .ZN(_26117_)
  );
  AND2_X1 _34253_ (
    .A1(_00008_[0]),
    .A2(_26117_),
    .ZN(_26118_)
  );
  AND2_X1 _34254_ (
    .A1(_26115_),
    .A2(_26118_),
    .ZN(_26119_)
  );
  INV_X1 _34255_ (
    .A(_26119_),
    .ZN(_26120_)
  );
  AND2_X1 _34256_ (
    .A1(_26113_),
    .A2(_26120_),
    .ZN(_26121_)
  );
  AND2_X1 _34257_ (
    .A1(_00008_[1]),
    .A2(_26121_),
    .ZN(_26122_)
  );
  INV_X1 _34258_ (
    .A(_26122_),
    .ZN(_26123_)
  );
  AND2_X1 _34259_ (
    .A1(_21899_),
    .A2(_00008_[2]),
    .ZN(_26124_)
  );
  INV_X1 _34260_ (
    .A(_26124_),
    .ZN(_26125_)
  );
  AND2_X1 _34261_ (
    .A1(_21843_),
    .A2(_22149_),
    .ZN(_26126_)
  );
  INV_X1 _34262_ (
    .A(_26126_),
    .ZN(_26127_)
  );
  AND2_X1 _34263_ (
    .A1(_00008_[0]),
    .A2(_26127_),
    .ZN(_26128_)
  );
  AND2_X1 _34264_ (
    .A1(_26125_),
    .A2(_26128_),
    .ZN(_26129_)
  );
  INV_X1 _34265_ (
    .A(_26129_),
    .ZN(_26130_)
  );
  AND2_X1 _34266_ (
    .A1(_21577_),
    .A2(_22149_),
    .ZN(_26131_)
  );
  INV_X1 _34267_ (
    .A(_26131_),
    .ZN(_26132_)
  );
  AND2_X1 _34268_ (
    .A1(_21915_),
    .A2(_00008_[2]),
    .ZN(_26133_)
  );
  INV_X1 _34269_ (
    .A(_26133_),
    .ZN(_26134_)
  );
  AND2_X1 _34270_ (
    .A1(_26132_),
    .A2(_26134_),
    .ZN(_26135_)
  );
  AND2_X1 _34271_ (
    .A1(_22147_),
    .A2(_26135_),
    .ZN(_26136_)
  );
  INV_X1 _34272_ (
    .A(_26136_),
    .ZN(_26137_)
  );
  AND2_X1 _34273_ (
    .A1(_26130_),
    .A2(_26137_),
    .ZN(_26138_)
  );
  AND2_X1 _34274_ (
    .A1(_22148_),
    .A2(_26138_),
    .ZN(_26139_)
  );
  INV_X1 _34275_ (
    .A(_26139_),
    .ZN(_26140_)
  );
  AND2_X1 _34276_ (
    .A1(_00008_[3]),
    .A2(_26123_),
    .ZN(_26141_)
  );
  AND2_X1 _34277_ (
    .A1(_26140_),
    .A2(_26141_),
    .ZN(_26142_)
  );
  INV_X1 _34278_ (
    .A(_26142_),
    .ZN(_26143_)
  );
  AND2_X1 _34279_ (
    .A1(_22150_),
    .A2(_26106_),
    .ZN(_26144_)
  );
  INV_X1 _34280_ (
    .A(_26144_),
    .ZN(_26145_)
  );
  AND2_X1 _34281_ (
    .A1(_00008_[4]),
    .A2(_26145_),
    .ZN(_26146_)
  );
  AND2_X1 _34282_ (
    .A1(_26143_),
    .A2(_26146_),
    .ZN(_26147_)
  );
  INV_X1 _34283_ (
    .A(_26147_),
    .ZN(_26148_)
  );
  AND2_X1 _34284_ (
    .A1(\cpuregs[10] [19]),
    .A2(_22149_),
    .ZN(_26149_)
  );
  INV_X1 _34285_ (
    .A(_26149_),
    .ZN(_26150_)
  );
  AND2_X1 _34286_ (
    .A1(\cpuregs[14] [19]),
    .A2(_00008_[2]),
    .ZN(_26151_)
  );
  INV_X1 _34287_ (
    .A(_26151_),
    .ZN(_26152_)
  );
  AND2_X1 _34288_ (
    .A1(_22147_),
    .A2(_26152_),
    .ZN(_26153_)
  );
  AND2_X1 _34289_ (
    .A1(_26150_),
    .A2(_26153_),
    .ZN(_26154_)
  );
  INV_X1 _34290_ (
    .A(_26154_),
    .ZN(_26155_)
  );
  AND2_X1 _34291_ (
    .A1(\cpuregs[15] [19]),
    .A2(_00008_[2]),
    .ZN(_26156_)
  );
  INV_X1 _34292_ (
    .A(_26156_),
    .ZN(_26157_)
  );
  AND2_X1 _34293_ (
    .A1(\cpuregs[11] [19]),
    .A2(_22149_),
    .ZN(_26158_)
  );
  INV_X1 _34294_ (
    .A(_26158_),
    .ZN(_26159_)
  );
  AND2_X1 _34295_ (
    .A1(_00008_[0]),
    .A2(_26159_),
    .ZN(_26160_)
  );
  AND2_X1 _34296_ (
    .A1(_26157_),
    .A2(_26160_),
    .ZN(_26161_)
  );
  INV_X1 _34297_ (
    .A(_26161_),
    .ZN(_26162_)
  );
  AND2_X1 _34298_ (
    .A1(_26155_),
    .A2(_26162_),
    .ZN(_26163_)
  );
  INV_X1 _34299_ (
    .A(_26163_),
    .ZN(_26164_)
  );
  AND2_X1 _34300_ (
    .A1(_00008_[3]),
    .A2(_26164_),
    .ZN(_26165_)
  );
  INV_X1 _34301_ (
    .A(_26165_),
    .ZN(_26166_)
  );
  AND2_X1 _34302_ (
    .A1(\cpuregs[2] [19]),
    .A2(_22149_),
    .ZN(_26167_)
  );
  INV_X1 _34303_ (
    .A(_26167_),
    .ZN(_26168_)
  );
  AND2_X1 _34304_ (
    .A1(\cpuregs[6] [19]),
    .A2(_00008_[2]),
    .ZN(_26169_)
  );
  INV_X1 _34305_ (
    .A(_26169_),
    .ZN(_26170_)
  );
  AND2_X1 _34306_ (
    .A1(_22147_),
    .A2(_26170_),
    .ZN(_26171_)
  );
  AND2_X1 _34307_ (
    .A1(_26168_),
    .A2(_26171_),
    .ZN(_26172_)
  );
  INV_X1 _34308_ (
    .A(_26172_),
    .ZN(_26173_)
  );
  AND2_X1 _34309_ (
    .A1(\cpuregs[3] [19]),
    .A2(_22149_),
    .ZN(_26174_)
  );
  INV_X1 _34310_ (
    .A(_26174_),
    .ZN(_26175_)
  );
  AND2_X1 _34311_ (
    .A1(\cpuregs[7] [19]),
    .A2(_00008_[2]),
    .ZN(_26176_)
  );
  INV_X1 _34312_ (
    .A(_26176_),
    .ZN(_26177_)
  );
  AND2_X1 _34313_ (
    .A1(_00008_[0]),
    .A2(_26177_),
    .ZN(_26178_)
  );
  AND2_X1 _34314_ (
    .A1(_26175_),
    .A2(_26178_),
    .ZN(_26179_)
  );
  INV_X1 _34315_ (
    .A(_26179_),
    .ZN(_26180_)
  );
  AND2_X1 _34316_ (
    .A1(_26173_),
    .A2(_26180_),
    .ZN(_26181_)
  );
  INV_X1 _34317_ (
    .A(_26181_),
    .ZN(_26182_)
  );
  AND2_X1 _34318_ (
    .A1(_22150_),
    .A2(_26182_),
    .ZN(_26183_)
  );
  INV_X1 _34319_ (
    .A(_26183_),
    .ZN(_26184_)
  );
  AND2_X1 _34320_ (
    .A1(\cpuregs[8] [19]),
    .A2(_22149_),
    .ZN(_26185_)
  );
  INV_X1 _34321_ (
    .A(_26185_),
    .ZN(_26186_)
  );
  AND2_X1 _34322_ (
    .A1(\cpuregs[12] [19]),
    .A2(_00008_[2]),
    .ZN(_26187_)
  );
  INV_X1 _34323_ (
    .A(_26187_),
    .ZN(_26188_)
  );
  AND2_X1 _34324_ (
    .A1(_22147_),
    .A2(_26188_),
    .ZN(_26189_)
  );
  AND2_X1 _34325_ (
    .A1(_26186_),
    .A2(_26189_),
    .ZN(_26190_)
  );
  INV_X1 _34326_ (
    .A(_26190_),
    .ZN(_26191_)
  );
  AND2_X1 _34327_ (
    .A1(\cpuregs[13] [19]),
    .A2(_00008_[2]),
    .ZN(_26192_)
  );
  INV_X1 _34328_ (
    .A(_26192_),
    .ZN(_26193_)
  );
  AND2_X1 _34329_ (
    .A1(\cpuregs[9] [19]),
    .A2(_22149_),
    .ZN(_26194_)
  );
  INV_X1 _34330_ (
    .A(_26194_),
    .ZN(_26195_)
  );
  AND2_X1 _34331_ (
    .A1(_00008_[0]),
    .A2(_26195_),
    .ZN(_26196_)
  );
  AND2_X1 _34332_ (
    .A1(_26193_),
    .A2(_26196_),
    .ZN(_26197_)
  );
  INV_X1 _34333_ (
    .A(_26197_),
    .ZN(_26198_)
  );
  AND2_X1 _34334_ (
    .A1(_26191_),
    .A2(_26198_),
    .ZN(_26199_)
  );
  AND2_X1 _34335_ (
    .A1(\cpuregs[0] [19]),
    .A2(_22149_),
    .ZN(_26200_)
  );
  INV_X1 _34336_ (
    .A(_26200_),
    .ZN(_26201_)
  );
  AND2_X1 _34337_ (
    .A1(\cpuregs[4] [19]),
    .A2(_00008_[2]),
    .ZN(_26202_)
  );
  INV_X1 _34338_ (
    .A(_26202_),
    .ZN(_26203_)
  );
  AND2_X1 _34339_ (
    .A1(_22147_),
    .A2(_26203_),
    .ZN(_26204_)
  );
  AND2_X1 _34340_ (
    .A1(_26201_),
    .A2(_26204_),
    .ZN(_26205_)
  );
  INV_X1 _34341_ (
    .A(_26205_),
    .ZN(_26206_)
  );
  AND2_X1 _34342_ (
    .A1(\cpuregs[1] [19]),
    .A2(_22149_),
    .ZN(_26207_)
  );
  INV_X1 _34343_ (
    .A(_26207_),
    .ZN(_26208_)
  );
  AND2_X1 _34344_ (
    .A1(\cpuregs[5] [19]),
    .A2(_00008_[2]),
    .ZN(_26209_)
  );
  INV_X1 _34345_ (
    .A(_26209_),
    .ZN(_26210_)
  );
  AND2_X1 _34346_ (
    .A1(_00008_[0]),
    .A2(_26210_),
    .ZN(_26211_)
  );
  AND2_X1 _34347_ (
    .A1(_26208_),
    .A2(_26211_),
    .ZN(_26212_)
  );
  INV_X1 _34348_ (
    .A(_26212_),
    .ZN(_26213_)
  );
  AND2_X1 _34349_ (
    .A1(_00008_[3]),
    .A2(_26199_),
    .ZN(_26214_)
  );
  INV_X1 _34350_ (
    .A(_26214_),
    .ZN(_26215_)
  );
  AND2_X1 _34351_ (
    .A1(_22150_),
    .A2(_26213_),
    .ZN(_26216_)
  );
  AND2_X1 _34352_ (
    .A1(_26206_),
    .A2(_26216_),
    .ZN(_26217_)
  );
  INV_X1 _34353_ (
    .A(_26217_),
    .ZN(_26218_)
  );
  AND2_X1 _34354_ (
    .A1(_26215_),
    .A2(_26218_),
    .ZN(_26219_)
  );
  INV_X1 _34355_ (
    .A(_26219_),
    .ZN(_26220_)
  );
  AND2_X1 _34356_ (
    .A1(_22148_),
    .A2(_26220_),
    .ZN(_26221_)
  );
  INV_X1 _34357_ (
    .A(_26221_),
    .ZN(_26222_)
  );
  AND2_X1 _34358_ (
    .A1(_00008_[1]),
    .A2(_26184_),
    .ZN(_26223_)
  );
  AND2_X1 _34359_ (
    .A1(_26166_),
    .A2(_26223_),
    .ZN(_26224_)
  );
  INV_X1 _34360_ (
    .A(_26224_),
    .ZN(_26225_)
  );
  AND2_X1 _34361_ (
    .A1(_22151_),
    .A2(_26225_),
    .ZN(_26226_)
  );
  AND2_X1 _34362_ (
    .A1(_26222_),
    .A2(_26226_),
    .ZN(_26227_)
  );
  INV_X1 _34363_ (
    .A(_26227_),
    .ZN(_26228_)
  );
  AND2_X1 _34364_ (
    .A1(_22546_),
    .A2(_26148_),
    .ZN(_26229_)
  );
  AND2_X1 _34365_ (
    .A1(_26228_),
    .A2(_26229_),
    .ZN(_26230_)
  );
  INV_X1 _34366_ (
    .A(_26230_),
    .ZN(_26231_)
  );
  AND2_X1 _34367_ (
    .A1(_26071_),
    .A2(_26231_),
    .ZN(_26232_)
  );
  INV_X1 _34368_ (
    .A(_26232_),
    .ZN(_26233_)
  );
  AND2_X1 _34369_ (
    .A1(_22271_),
    .A2(_26233_),
    .ZN(_26234_)
  );
  INV_X1 _34370_ (
    .A(_26234_),
    .ZN(_26235_)
  );
  AND2_X1 _34371_ (
    .A1(reg_op1[18]),
    .A2(_22285_),
    .ZN(_26236_)
  );
  INV_X1 _34372_ (
    .A(_26236_),
    .ZN(_26237_)
  );
  AND2_X1 _34373_ (
    .A1(_25624_),
    .A2(_26237_),
    .ZN(_26238_)
  );
  AND2_X1 _34374_ (
    .A1(reg_op1[23]),
    .A2(_22290_),
    .ZN(_26239_)
  );
  INV_X1 _34375_ (
    .A(_26239_),
    .ZN(_26240_)
  );
  AND2_X1 _34376_ (
    .A1(_25621_),
    .A2(_26240_),
    .ZN(_26241_)
  );
  AND2_X1 _34377_ (
    .A1(_22573_),
    .A2(_26241_),
    .ZN(_26242_)
  );
  INV_X1 _34378_ (
    .A(_26242_),
    .ZN(_26243_)
  );
  AND2_X1 _34379_ (
    .A1(_22572_),
    .A2(_26238_),
    .ZN(_26244_)
  );
  INV_X1 _34380_ (
    .A(_26244_),
    .ZN(_26245_)
  );
  AND2_X1 _34381_ (
    .A1(_22295_),
    .A2(_26245_),
    .ZN(_26246_)
  );
  AND2_X1 _34382_ (
    .A1(_26243_),
    .A2(_26246_),
    .ZN(_26247_)
  );
  INV_X1 _34383_ (
    .A(_26247_),
    .ZN(_26248_)
  );
  AND2_X1 _34384_ (
    .A1(reg_op1[19]),
    .A2(decoded_imm[19]),
    .ZN(_26249_)
  );
  INV_X1 _34385_ (
    .A(_26249_),
    .ZN(_26250_)
  );
  AND2_X1 _34386_ (
    .A1(_21186_),
    .A2(_21990_),
    .ZN(_26251_)
  );
  INV_X1 _34387_ (
    .A(_26251_),
    .ZN(_26252_)
  );
  AND2_X1 _34388_ (
    .A1(_26250_),
    .A2(_26252_),
    .ZN(_26253_)
  );
  INV_X1 _34389_ (
    .A(_26253_),
    .ZN(_26254_)
  );
  AND2_X1 _34390_ (
    .A1(_26054_),
    .A2(_26254_),
    .ZN(_26255_)
  );
  AND2_X1 _34391_ (
    .A1(_26060_),
    .A2(_26255_),
    .ZN(_26256_)
  );
  INV_X1 _34392_ (
    .A(_26256_),
    .ZN(_26257_)
  );
  AND2_X1 _34393_ (
    .A1(_26059_),
    .A2(_26253_),
    .ZN(_26258_)
  );
  INV_X1 _34394_ (
    .A(_26258_),
    .ZN(_26259_)
  );
  AND2_X1 _34395_ (
    .A1(_26053_),
    .A2(_26253_),
    .ZN(_26260_)
  );
  INV_X1 _34396_ (
    .A(_26260_),
    .ZN(_26261_)
  );
  AND2_X1 _34397_ (
    .A1(_22559_),
    .A2(_26261_),
    .ZN(_26262_)
  );
  AND2_X1 _34398_ (
    .A1(_26259_),
    .A2(_26262_),
    .ZN(_26263_)
  );
  AND2_X1 _34399_ (
    .A1(_26257_),
    .A2(_26263_),
    .ZN(_26264_)
  );
  INV_X1 _34400_ (
    .A(_26264_),
    .ZN(_26265_)
  );
  AND2_X1 _34401_ (
    .A1(_26235_),
    .A2(_26248_),
    .ZN(_26266_)
  );
  AND2_X1 _34402_ (
    .A1(_26265_),
    .A2(_26266_),
    .ZN(_26267_)
  );
  AND2_X1 _34403_ (
    .A1(_22333_),
    .A2(_26267_),
    .ZN(_26268_)
  );
  INV_X1 _34404_ (
    .A(_26268_),
    .ZN(_26269_)
  );
  AND2_X1 _34405_ (
    .A1(_26069_),
    .A2(_26269_),
    .ZN(_00076_)
  );
  AND2_X1 _34406_ (
    .A1(_21187_),
    .A2(_22334_),
    .ZN(_26270_)
  );
  INV_X1 _34407_ (
    .A(_26270_),
    .ZN(_26271_)
  );
  AND2_X1 _34408_ (
    .A1(reg_pc[20]),
    .A2(_22335_),
    .ZN(_26272_)
  );
  INV_X1 _34409_ (
    .A(_26272_),
    .ZN(_26273_)
  );
  AND2_X1 _34410_ (
    .A1(_21451_),
    .A2(_22149_),
    .ZN(_26274_)
  );
  INV_X1 _34411_ (
    .A(_26274_),
    .ZN(_26275_)
  );
  AND2_X1 _34412_ (
    .A1(_21662_),
    .A2(_00008_[2]),
    .ZN(_26276_)
  );
  INV_X1 _34413_ (
    .A(_26276_),
    .ZN(_26277_)
  );
  AND2_X1 _34414_ (
    .A1(_26275_),
    .A2(_26277_),
    .ZN(_26278_)
  );
  AND2_X1 _34415_ (
    .A1(_22147_),
    .A2(_26278_),
    .ZN(_26279_)
  );
  INV_X1 _34416_ (
    .A(_26279_),
    .ZN(_26280_)
  );
  AND2_X1 _34417_ (
    .A1(_21772_),
    .A2(_00008_[2]),
    .ZN(_26281_)
  );
  INV_X1 _34418_ (
    .A(_26281_),
    .ZN(_26282_)
  );
  AND2_X1 _34419_ (
    .A1(_21473_),
    .A2(_22149_),
    .ZN(_26283_)
  );
  INV_X1 _34420_ (
    .A(_26283_),
    .ZN(_26284_)
  );
  AND2_X1 _34421_ (
    .A1(_00008_[0]),
    .A2(_26282_),
    .ZN(_26285_)
  );
  AND2_X1 _34422_ (
    .A1(_26284_),
    .A2(_26285_),
    .ZN(_26286_)
  );
  INV_X1 _34423_ (
    .A(_26286_),
    .ZN(_26287_)
  );
  AND2_X1 _34424_ (
    .A1(_26280_),
    .A2(_26287_),
    .ZN(_26288_)
  );
  AND2_X1 _34425_ (
    .A1(_22148_),
    .A2(_26288_),
    .ZN(_26289_)
  );
  INV_X1 _34426_ (
    .A(_26289_),
    .ZN(_26290_)
  );
  AND2_X1 _34427_ (
    .A1(_21606_),
    .A2(_22149_),
    .ZN(_26291_)
  );
  INV_X1 _34428_ (
    .A(_26291_),
    .ZN(_26292_)
  );
  AND2_X1 _34429_ (
    .A1(_21426_),
    .A2(_00008_[2]),
    .ZN(_26293_)
  );
  INV_X1 _34430_ (
    .A(_26293_),
    .ZN(_26294_)
  );
  AND2_X1 _34431_ (
    .A1(_26292_),
    .A2(_26294_),
    .ZN(_26295_)
  );
  AND2_X1 _34432_ (
    .A1(_22147_),
    .A2(_26295_),
    .ZN(_26296_)
  );
  INV_X1 _34433_ (
    .A(_26296_),
    .ZN(_26297_)
  );
  AND2_X1 _34434_ (
    .A1(_21385_),
    .A2(_00008_[2]),
    .ZN(_26298_)
  );
  INV_X1 _34435_ (
    .A(_26298_),
    .ZN(_26299_)
  );
  AND2_X1 _34436_ (
    .A1(_21631_),
    .A2(_22149_),
    .ZN(_26300_)
  );
  INV_X1 _34437_ (
    .A(_26300_),
    .ZN(_26301_)
  );
  AND2_X1 _34438_ (
    .A1(_00008_[0]),
    .A2(_26301_),
    .ZN(_26302_)
  );
  AND2_X1 _34439_ (
    .A1(_26299_),
    .A2(_26302_),
    .ZN(_26303_)
  );
  INV_X1 _34440_ (
    .A(_26303_),
    .ZN(_26304_)
  );
  AND2_X1 _34441_ (
    .A1(_26297_),
    .A2(_26304_),
    .ZN(_26305_)
  );
  AND2_X1 _34442_ (
    .A1(_00008_[1]),
    .A2(_26305_),
    .ZN(_26306_)
  );
  INV_X1 _34443_ (
    .A(_26306_),
    .ZN(_26307_)
  );
  AND2_X1 _34444_ (
    .A1(_26290_),
    .A2(_26307_),
    .ZN(_26308_)
  );
  AND2_X1 _34445_ (
    .A1(\cpuregs[27] [20]),
    .A2(_00008_[0]),
    .ZN(_26309_)
  );
  INV_X1 _34446_ (
    .A(_26309_),
    .ZN(_26310_)
  );
  AND2_X1 _34447_ (
    .A1(\cpuregs[26] [20]),
    .A2(_22147_),
    .ZN(_26311_)
  );
  INV_X1 _34448_ (
    .A(_26311_),
    .ZN(_26312_)
  );
  AND2_X1 _34449_ (
    .A1(_22149_),
    .A2(_26312_),
    .ZN(_26313_)
  );
  AND2_X1 _34450_ (
    .A1(_26310_),
    .A2(_26313_),
    .ZN(_26314_)
  );
  INV_X1 _34451_ (
    .A(_26314_),
    .ZN(_26315_)
  );
  AND2_X1 _34452_ (
    .A1(\cpuregs[31] [20]),
    .A2(_00008_[0]),
    .ZN(_26316_)
  );
  INV_X1 _34453_ (
    .A(_26316_),
    .ZN(_26317_)
  );
  AND2_X1 _34454_ (
    .A1(\cpuregs[30] [20]),
    .A2(_22147_),
    .ZN(_26318_)
  );
  INV_X1 _34455_ (
    .A(_26318_),
    .ZN(_26319_)
  );
  AND2_X1 _34456_ (
    .A1(_00008_[2]),
    .A2(_26319_),
    .ZN(_26320_)
  );
  AND2_X1 _34457_ (
    .A1(_26317_),
    .A2(_26320_),
    .ZN(_26321_)
  );
  INV_X1 _34458_ (
    .A(_26321_),
    .ZN(_26322_)
  );
  AND2_X1 _34459_ (
    .A1(_26315_),
    .A2(_26322_),
    .ZN(_26323_)
  );
  INV_X1 _34460_ (
    .A(_26323_),
    .ZN(_26324_)
  );
  AND2_X1 _34461_ (
    .A1(_00008_[1]),
    .A2(_26324_),
    .ZN(_26325_)
  );
  INV_X1 _34462_ (
    .A(_26325_),
    .ZN(_26326_)
  );
  AND2_X1 _34463_ (
    .A1(\cpuregs[25] [20]),
    .A2(_00008_[0]),
    .ZN(_26327_)
  );
  INV_X1 _34464_ (
    .A(_26327_),
    .ZN(_26328_)
  );
  AND2_X1 _34465_ (
    .A1(\cpuregs[24] [20]),
    .A2(_22147_),
    .ZN(_26329_)
  );
  INV_X1 _34466_ (
    .A(_26329_),
    .ZN(_26330_)
  );
  AND2_X1 _34467_ (
    .A1(_22149_),
    .A2(_26330_),
    .ZN(_26331_)
  );
  AND2_X1 _34468_ (
    .A1(_26328_),
    .A2(_26331_),
    .ZN(_26332_)
  );
  INV_X1 _34469_ (
    .A(_26332_),
    .ZN(_26333_)
  );
  AND2_X1 _34470_ (
    .A1(\cpuregs[29] [20]),
    .A2(_00008_[0]),
    .ZN(_26334_)
  );
  INV_X1 _34471_ (
    .A(_26334_),
    .ZN(_26335_)
  );
  AND2_X1 _34472_ (
    .A1(\cpuregs[28] [20]),
    .A2(_22147_),
    .ZN(_26336_)
  );
  INV_X1 _34473_ (
    .A(_26336_),
    .ZN(_26337_)
  );
  AND2_X1 _34474_ (
    .A1(_00008_[2]),
    .A2(_26337_),
    .ZN(_26338_)
  );
  AND2_X1 _34475_ (
    .A1(_26335_),
    .A2(_26338_),
    .ZN(_26339_)
  );
  INV_X1 _34476_ (
    .A(_26339_),
    .ZN(_26340_)
  );
  AND2_X1 _34477_ (
    .A1(_26333_),
    .A2(_26340_),
    .ZN(_26341_)
  );
  INV_X1 _34478_ (
    .A(_26341_),
    .ZN(_26342_)
  );
  AND2_X1 _34479_ (
    .A1(_22148_),
    .A2(_26342_),
    .ZN(_26343_)
  );
  INV_X1 _34480_ (
    .A(_26343_),
    .ZN(_26344_)
  );
  AND2_X1 _34481_ (
    .A1(_00008_[3]),
    .A2(_26326_),
    .ZN(_26345_)
  );
  AND2_X1 _34482_ (
    .A1(_26344_),
    .A2(_26345_),
    .ZN(_26346_)
  );
  INV_X1 _34483_ (
    .A(_26346_),
    .ZN(_26347_)
  );
  AND2_X1 _34484_ (
    .A1(_22150_),
    .A2(_26308_),
    .ZN(_26348_)
  );
  INV_X1 _34485_ (
    .A(_26348_),
    .ZN(_26349_)
  );
  AND2_X1 _34486_ (
    .A1(_00008_[4]),
    .A2(_26349_),
    .ZN(_26350_)
  );
  AND2_X1 _34487_ (
    .A1(_26347_),
    .A2(_26350_),
    .ZN(_26351_)
  );
  INV_X1 _34488_ (
    .A(_26351_),
    .ZN(_26352_)
  );
  AND2_X1 _34489_ (
    .A1(\cpuregs[10] [20]),
    .A2(_22149_),
    .ZN(_26353_)
  );
  INV_X1 _34490_ (
    .A(_26353_),
    .ZN(_26354_)
  );
  AND2_X1 _34491_ (
    .A1(\cpuregs[14] [20]),
    .A2(_00008_[2]),
    .ZN(_26355_)
  );
  INV_X1 _34492_ (
    .A(_26355_),
    .ZN(_26356_)
  );
  AND2_X1 _34493_ (
    .A1(_22147_),
    .A2(_26356_),
    .ZN(_26357_)
  );
  AND2_X1 _34494_ (
    .A1(_26354_),
    .A2(_26357_),
    .ZN(_26358_)
  );
  INV_X1 _34495_ (
    .A(_26358_),
    .ZN(_26359_)
  );
  AND2_X1 _34496_ (
    .A1(\cpuregs[15] [20]),
    .A2(_00008_[2]),
    .ZN(_26360_)
  );
  INV_X1 _34497_ (
    .A(_26360_),
    .ZN(_26361_)
  );
  AND2_X1 _34498_ (
    .A1(\cpuregs[11] [20]),
    .A2(_22149_),
    .ZN(_26362_)
  );
  INV_X1 _34499_ (
    .A(_26362_),
    .ZN(_26363_)
  );
  AND2_X1 _34500_ (
    .A1(_00008_[0]),
    .A2(_26363_),
    .ZN(_26364_)
  );
  AND2_X1 _34501_ (
    .A1(_26361_),
    .A2(_26364_),
    .ZN(_26365_)
  );
  INV_X1 _34502_ (
    .A(_26365_),
    .ZN(_26366_)
  );
  AND2_X1 _34503_ (
    .A1(_26359_),
    .A2(_26366_),
    .ZN(_26367_)
  );
  INV_X1 _34504_ (
    .A(_26367_),
    .ZN(_26368_)
  );
  AND2_X1 _34505_ (
    .A1(_00008_[3]),
    .A2(_26368_),
    .ZN(_26369_)
  );
  INV_X1 _34506_ (
    .A(_26369_),
    .ZN(_26370_)
  );
  AND2_X1 _34507_ (
    .A1(\cpuregs[2] [20]),
    .A2(_22149_),
    .ZN(_26371_)
  );
  INV_X1 _34508_ (
    .A(_26371_),
    .ZN(_26372_)
  );
  AND2_X1 _34509_ (
    .A1(\cpuregs[6] [20]),
    .A2(_00008_[2]),
    .ZN(_26373_)
  );
  INV_X1 _34510_ (
    .A(_26373_),
    .ZN(_26374_)
  );
  AND2_X1 _34511_ (
    .A1(_22147_),
    .A2(_26374_),
    .ZN(_26375_)
  );
  AND2_X1 _34512_ (
    .A1(_26372_),
    .A2(_26375_),
    .ZN(_26376_)
  );
  INV_X1 _34513_ (
    .A(_26376_),
    .ZN(_26377_)
  );
  AND2_X1 _34514_ (
    .A1(\cpuregs[3] [20]),
    .A2(_22149_),
    .ZN(_26378_)
  );
  INV_X1 _34515_ (
    .A(_26378_),
    .ZN(_26379_)
  );
  AND2_X1 _34516_ (
    .A1(\cpuregs[7] [20]),
    .A2(_00008_[2]),
    .ZN(_26380_)
  );
  INV_X1 _34517_ (
    .A(_26380_),
    .ZN(_26381_)
  );
  AND2_X1 _34518_ (
    .A1(_00008_[0]),
    .A2(_26381_),
    .ZN(_26382_)
  );
  AND2_X1 _34519_ (
    .A1(_26379_),
    .A2(_26382_),
    .ZN(_26383_)
  );
  INV_X1 _34520_ (
    .A(_26383_),
    .ZN(_26384_)
  );
  AND2_X1 _34521_ (
    .A1(_26377_),
    .A2(_26384_),
    .ZN(_26385_)
  );
  INV_X1 _34522_ (
    .A(_26385_),
    .ZN(_26386_)
  );
  AND2_X1 _34523_ (
    .A1(_22150_),
    .A2(_26386_),
    .ZN(_26387_)
  );
  INV_X1 _34524_ (
    .A(_26387_),
    .ZN(_26388_)
  );
  AND2_X1 _34525_ (
    .A1(\cpuregs[8] [20]),
    .A2(_22149_),
    .ZN(_26389_)
  );
  INV_X1 _34526_ (
    .A(_26389_),
    .ZN(_26390_)
  );
  AND2_X1 _34527_ (
    .A1(\cpuregs[12] [20]),
    .A2(_00008_[2]),
    .ZN(_26391_)
  );
  INV_X1 _34528_ (
    .A(_26391_),
    .ZN(_26392_)
  );
  AND2_X1 _34529_ (
    .A1(_22147_),
    .A2(_26392_),
    .ZN(_26393_)
  );
  AND2_X1 _34530_ (
    .A1(_26390_),
    .A2(_26393_),
    .ZN(_26394_)
  );
  INV_X1 _34531_ (
    .A(_26394_),
    .ZN(_26395_)
  );
  AND2_X1 _34532_ (
    .A1(\cpuregs[13] [20]),
    .A2(_00008_[2]),
    .ZN(_26396_)
  );
  INV_X1 _34533_ (
    .A(_26396_),
    .ZN(_26397_)
  );
  AND2_X1 _34534_ (
    .A1(\cpuregs[9] [20]),
    .A2(_22149_),
    .ZN(_26398_)
  );
  INV_X1 _34535_ (
    .A(_26398_),
    .ZN(_26399_)
  );
  AND2_X1 _34536_ (
    .A1(_00008_[0]),
    .A2(_26399_),
    .ZN(_26400_)
  );
  AND2_X1 _34537_ (
    .A1(_26397_),
    .A2(_26400_),
    .ZN(_26401_)
  );
  INV_X1 _34538_ (
    .A(_26401_),
    .ZN(_26402_)
  );
  AND2_X1 _34539_ (
    .A1(_26395_),
    .A2(_26402_),
    .ZN(_26403_)
  );
  AND2_X1 _34540_ (
    .A1(\cpuregs[0] [20]),
    .A2(_22149_),
    .ZN(_26404_)
  );
  INV_X1 _34541_ (
    .A(_26404_),
    .ZN(_26405_)
  );
  AND2_X1 _34542_ (
    .A1(\cpuregs[4] [20]),
    .A2(_00008_[2]),
    .ZN(_26406_)
  );
  INV_X1 _34543_ (
    .A(_26406_),
    .ZN(_26407_)
  );
  AND2_X1 _34544_ (
    .A1(_22147_),
    .A2(_26407_),
    .ZN(_26408_)
  );
  AND2_X1 _34545_ (
    .A1(_26405_),
    .A2(_26408_),
    .ZN(_26409_)
  );
  INV_X1 _34546_ (
    .A(_26409_),
    .ZN(_26410_)
  );
  AND2_X1 _34547_ (
    .A1(\cpuregs[1] [20]),
    .A2(_22149_),
    .ZN(_26411_)
  );
  INV_X1 _34548_ (
    .A(_26411_),
    .ZN(_26412_)
  );
  AND2_X1 _34549_ (
    .A1(\cpuregs[5] [20]),
    .A2(_00008_[2]),
    .ZN(_26413_)
  );
  INV_X1 _34550_ (
    .A(_26413_),
    .ZN(_26414_)
  );
  AND2_X1 _34551_ (
    .A1(_00008_[0]),
    .A2(_26414_),
    .ZN(_26415_)
  );
  AND2_X1 _34552_ (
    .A1(_26412_),
    .A2(_26415_),
    .ZN(_26416_)
  );
  INV_X1 _34553_ (
    .A(_26416_),
    .ZN(_26417_)
  );
  AND2_X1 _34554_ (
    .A1(_00008_[3]),
    .A2(_26403_),
    .ZN(_26418_)
  );
  INV_X1 _34555_ (
    .A(_26418_),
    .ZN(_26419_)
  );
  AND2_X1 _34556_ (
    .A1(_22150_),
    .A2(_26417_),
    .ZN(_26420_)
  );
  AND2_X1 _34557_ (
    .A1(_26410_),
    .A2(_26420_),
    .ZN(_26421_)
  );
  INV_X1 _34558_ (
    .A(_26421_),
    .ZN(_26422_)
  );
  AND2_X1 _34559_ (
    .A1(_26419_),
    .A2(_26422_),
    .ZN(_26423_)
  );
  INV_X1 _34560_ (
    .A(_26423_),
    .ZN(_26424_)
  );
  AND2_X1 _34561_ (
    .A1(_22148_),
    .A2(_26424_),
    .ZN(_26425_)
  );
  INV_X1 _34562_ (
    .A(_26425_),
    .ZN(_26426_)
  );
  AND2_X1 _34563_ (
    .A1(_00008_[1]),
    .A2(_26388_),
    .ZN(_26427_)
  );
  AND2_X1 _34564_ (
    .A1(_26370_),
    .A2(_26427_),
    .ZN(_26428_)
  );
  INV_X1 _34565_ (
    .A(_26428_),
    .ZN(_26429_)
  );
  AND2_X1 _34566_ (
    .A1(_22151_),
    .A2(_26429_),
    .ZN(_26430_)
  );
  AND2_X1 _34567_ (
    .A1(_26426_),
    .A2(_26430_),
    .ZN(_26431_)
  );
  INV_X1 _34568_ (
    .A(_26431_),
    .ZN(_26432_)
  );
  AND2_X1 _34569_ (
    .A1(_22546_),
    .A2(_26352_),
    .ZN(_26433_)
  );
  AND2_X1 _34570_ (
    .A1(_26432_),
    .A2(_26433_),
    .ZN(_26434_)
  );
  INV_X1 _34571_ (
    .A(_26434_),
    .ZN(_26435_)
  );
  AND2_X1 _34572_ (
    .A1(_26273_),
    .A2(_26435_),
    .ZN(_26436_)
  );
  INV_X1 _34573_ (
    .A(_26436_),
    .ZN(_26437_)
  );
  AND2_X1 _34574_ (
    .A1(_22271_),
    .A2(_26437_),
    .ZN(_26438_)
  );
  INV_X1 _34575_ (
    .A(_26438_),
    .ZN(_26439_)
  );
  AND2_X1 _34576_ (
    .A1(reg_op1[19]),
    .A2(_22285_),
    .ZN(_26440_)
  );
  INV_X1 _34577_ (
    .A(_26440_),
    .ZN(_26441_)
  );
  AND2_X1 _34578_ (
    .A1(_25846_),
    .A2(_26441_),
    .ZN(_26442_)
  );
  AND2_X1 _34579_ (
    .A1(reg_op1[24]),
    .A2(_22290_),
    .ZN(_26443_)
  );
  INV_X1 _34580_ (
    .A(_26443_),
    .ZN(_26444_)
  );
  AND2_X1 _34581_ (
    .A1(_25843_),
    .A2(_26444_),
    .ZN(_26445_)
  );
  AND2_X1 _34582_ (
    .A1(_22572_),
    .A2(_26442_),
    .ZN(_26446_)
  );
  INV_X1 _34583_ (
    .A(_26446_),
    .ZN(_26447_)
  );
  AND2_X1 _34584_ (
    .A1(_22573_),
    .A2(_26445_),
    .ZN(_26448_)
  );
  INV_X1 _34585_ (
    .A(_26448_),
    .ZN(_26449_)
  );
  AND2_X1 _34586_ (
    .A1(_22295_),
    .A2(_26449_),
    .ZN(_26450_)
  );
  AND2_X1 _34587_ (
    .A1(_26447_),
    .A2(_26450_),
    .ZN(_26451_)
  );
  INV_X1 _34588_ (
    .A(_26451_),
    .ZN(_26452_)
  );
  AND2_X1 _34589_ (
    .A1(_22333_),
    .A2(_26452_),
    .ZN(_26453_)
  );
  AND2_X1 _34590_ (
    .A1(_26439_),
    .A2(_26453_),
    .ZN(_26454_)
  );
  AND2_X1 _34591_ (
    .A1(reg_op1[20]),
    .A2(decoded_imm[20]),
    .ZN(_26455_)
  );
  INV_X1 _34592_ (
    .A(_26455_),
    .ZN(_26456_)
  );
  AND2_X1 _34593_ (
    .A1(_21187_),
    .A2(_21989_),
    .ZN(_26457_)
  );
  INV_X1 _34594_ (
    .A(_26457_),
    .ZN(_26458_)
  );
  AND2_X1 _34595_ (
    .A1(_26456_),
    .A2(_26458_),
    .ZN(_26459_)
  );
  INV_X1 _34596_ (
    .A(_26459_),
    .ZN(_26460_)
  );
  AND2_X1 _34597_ (
    .A1(_26250_),
    .A2(_26261_),
    .ZN(_26461_)
  );
  AND2_X1 _34598_ (
    .A1(_26259_),
    .A2(_26461_),
    .ZN(_26462_)
  );
  INV_X1 _34599_ (
    .A(_26462_),
    .ZN(_26463_)
  );
  AND2_X1 _34600_ (
    .A1(_26459_),
    .A2(_26463_),
    .ZN(_26464_)
  );
  INV_X1 _34601_ (
    .A(_26464_),
    .ZN(_26465_)
  );
  AND2_X1 _34602_ (
    .A1(_26460_),
    .A2(_26462_),
    .ZN(_26466_)
  );
  INV_X1 _34603_ (
    .A(_26466_),
    .ZN(_26467_)
  );
  AND2_X1 _34604_ (
    .A1(_22559_),
    .A2(_26467_),
    .ZN(_26468_)
  );
  AND2_X1 _34605_ (
    .A1(_26465_),
    .A2(_26468_),
    .ZN(_26469_)
  );
  INV_X1 _34606_ (
    .A(_26469_),
    .ZN(_26470_)
  );
  AND2_X1 _34607_ (
    .A1(_26454_),
    .A2(_26470_),
    .ZN(_26471_)
  );
  INV_X1 _34608_ (
    .A(_26471_),
    .ZN(_26472_)
  );
  AND2_X1 _34609_ (
    .A1(_26271_),
    .A2(_26472_),
    .ZN(_00077_)
  );
  AND2_X1 _34610_ (
    .A1(_21188_),
    .A2(_22334_),
    .ZN(_26473_)
  );
  INV_X1 _34611_ (
    .A(_26473_),
    .ZN(_26474_)
  );
  AND2_X1 _34612_ (
    .A1(reg_op1[21]),
    .A2(decoded_imm[21]),
    .ZN(_26475_)
  );
  INV_X1 _34613_ (
    .A(_26475_),
    .ZN(_26476_)
  );
  AND2_X1 _34614_ (
    .A1(_21188_),
    .A2(_21988_),
    .ZN(_26477_)
  );
  INV_X1 _34615_ (
    .A(_26477_),
    .ZN(_26478_)
  );
  AND2_X1 _34616_ (
    .A1(_26476_),
    .A2(_26478_),
    .ZN(_26479_)
  );
  INV_X1 _34617_ (
    .A(_26479_),
    .ZN(_26480_)
  );
  AND2_X1 _34618_ (
    .A1(_26456_),
    .A2(_26465_),
    .ZN(_26481_)
  );
  AND2_X1 _34619_ (
    .A1(_26480_),
    .A2(_26481_),
    .ZN(_26482_)
  );
  INV_X1 _34620_ (
    .A(_26482_),
    .ZN(_26483_)
  );
  AND2_X1 _34621_ (
    .A1(reg_pc[21]),
    .A2(_22335_),
    .ZN(_26484_)
  );
  INV_X1 _34622_ (
    .A(_26484_),
    .ZN(_26485_)
  );
  AND2_X1 _34623_ (
    .A1(\cpuregs[20] [21]),
    .A2(_00008_[2]),
    .ZN(_26486_)
  );
  INV_X1 _34624_ (
    .A(_26486_),
    .ZN(_26487_)
  );
  AND2_X1 _34625_ (
    .A1(\cpuregs[16] [21]),
    .A2(_22149_),
    .ZN(_26488_)
  );
  INV_X1 _34626_ (
    .A(_26488_),
    .ZN(_26489_)
  );
  AND2_X1 _34627_ (
    .A1(_26487_),
    .A2(_26489_),
    .ZN(_26490_)
  );
  AND2_X1 _34628_ (
    .A1(\cpuregs[21] [21]),
    .A2(_00008_[2]),
    .ZN(_26491_)
  );
  INV_X1 _34629_ (
    .A(_26491_),
    .ZN(_26492_)
  );
  AND2_X1 _34630_ (
    .A1(\cpuregs[17] [21]),
    .A2(_22149_),
    .ZN(_26493_)
  );
  INV_X1 _34631_ (
    .A(_26493_),
    .ZN(_26494_)
  );
  AND2_X1 _34632_ (
    .A1(_22147_),
    .A2(_26490_),
    .ZN(_26495_)
  );
  INV_X1 _34633_ (
    .A(_26495_),
    .ZN(_26496_)
  );
  AND2_X1 _34634_ (
    .A1(_00008_[0]),
    .A2(_26492_),
    .ZN(_26497_)
  );
  AND2_X1 _34635_ (
    .A1(_26494_),
    .A2(_26497_),
    .ZN(_26498_)
  );
  INV_X1 _34636_ (
    .A(_26498_),
    .ZN(_26499_)
  );
  AND2_X1 _34637_ (
    .A1(_26496_),
    .A2(_26499_),
    .ZN(_26500_)
  );
  INV_X1 _34638_ (
    .A(_26500_),
    .ZN(_26501_)
  );
  AND2_X1 _34639_ (
    .A1(_22150_),
    .A2(_26501_),
    .ZN(_26502_)
  );
  INV_X1 _34640_ (
    .A(_26502_),
    .ZN(_26503_)
  );
  AND2_X1 _34641_ (
    .A1(\cpuregs[28] [21]),
    .A2(_00008_[2]),
    .ZN(_26504_)
  );
  INV_X1 _34642_ (
    .A(_26504_),
    .ZN(_26505_)
  );
  AND2_X1 _34643_ (
    .A1(\cpuregs[24] [21]),
    .A2(_22149_),
    .ZN(_26506_)
  );
  INV_X1 _34644_ (
    .A(_26506_),
    .ZN(_26507_)
  );
  AND2_X1 _34645_ (
    .A1(_26505_),
    .A2(_26507_),
    .ZN(_26508_)
  );
  INV_X1 _34646_ (
    .A(_26508_),
    .ZN(_26509_)
  );
  AND2_X1 _34647_ (
    .A1(_22147_),
    .A2(_26509_),
    .ZN(_26510_)
  );
  INV_X1 _34648_ (
    .A(_26510_),
    .ZN(_26511_)
  );
  AND2_X1 _34649_ (
    .A1(\cpuregs[29] [21]),
    .A2(_00008_[2]),
    .ZN(_26512_)
  );
  INV_X1 _34650_ (
    .A(_26512_),
    .ZN(_26513_)
  );
  AND2_X1 _34651_ (
    .A1(\cpuregs[25] [21]),
    .A2(_22149_),
    .ZN(_26514_)
  );
  INV_X1 _34652_ (
    .A(_26514_),
    .ZN(_26515_)
  );
  AND2_X1 _34653_ (
    .A1(_26513_),
    .A2(_26515_),
    .ZN(_26516_)
  );
  INV_X1 _34654_ (
    .A(_26516_),
    .ZN(_26517_)
  );
  AND2_X1 _34655_ (
    .A1(_00008_[0]),
    .A2(_26517_),
    .ZN(_26518_)
  );
  INV_X1 _34656_ (
    .A(_26518_),
    .ZN(_26519_)
  );
  AND2_X1 _34657_ (
    .A1(_26511_),
    .A2(_26519_),
    .ZN(_26520_)
  );
  AND2_X1 _34658_ (
    .A1(_00008_[3]),
    .A2(_26520_),
    .ZN(_26521_)
  );
  INV_X1 _34659_ (
    .A(_26521_),
    .ZN(_26522_)
  );
  AND2_X1 _34660_ (
    .A1(\cpuregs[27] [21]),
    .A2(_00008_[0]),
    .ZN(_26523_)
  );
  INV_X1 _34661_ (
    .A(_26523_),
    .ZN(_26524_)
  );
  AND2_X1 _34662_ (
    .A1(\cpuregs[26] [21]),
    .A2(_22147_),
    .ZN(_26525_)
  );
  INV_X1 _34663_ (
    .A(_26525_),
    .ZN(_26526_)
  );
  AND2_X1 _34664_ (
    .A1(_22149_),
    .A2(_26526_),
    .ZN(_26527_)
  );
  AND2_X1 _34665_ (
    .A1(_26524_),
    .A2(_26527_),
    .ZN(_26528_)
  );
  INV_X1 _34666_ (
    .A(_26528_),
    .ZN(_26529_)
  );
  AND2_X1 _34667_ (
    .A1(\cpuregs[31] [21]),
    .A2(_00008_[0]),
    .ZN(_26530_)
  );
  INV_X1 _34668_ (
    .A(_26530_),
    .ZN(_26531_)
  );
  AND2_X1 _34669_ (
    .A1(\cpuregs[30] [21]),
    .A2(_22147_),
    .ZN(_26532_)
  );
  INV_X1 _34670_ (
    .A(_26532_),
    .ZN(_26533_)
  );
  AND2_X1 _34671_ (
    .A1(_00008_[2]),
    .A2(_26533_),
    .ZN(_26534_)
  );
  AND2_X1 _34672_ (
    .A1(_26531_),
    .A2(_26534_),
    .ZN(_26535_)
  );
  INV_X1 _34673_ (
    .A(_26535_),
    .ZN(_26536_)
  );
  AND2_X1 _34674_ (
    .A1(_26529_),
    .A2(_26536_),
    .ZN(_26537_)
  );
  INV_X1 _34675_ (
    .A(_26537_),
    .ZN(_26538_)
  );
  AND2_X1 _34676_ (
    .A1(_00008_[3]),
    .A2(_26538_),
    .ZN(_26539_)
  );
  INV_X1 _34677_ (
    .A(_26539_),
    .ZN(_26540_)
  );
  AND2_X1 _34678_ (
    .A1(\cpuregs[22] [21]),
    .A2(_00008_[2]),
    .ZN(_26541_)
  );
  INV_X1 _34679_ (
    .A(_26541_),
    .ZN(_26542_)
  );
  AND2_X1 _34680_ (
    .A1(\cpuregs[18] [21]),
    .A2(_22149_),
    .ZN(_26543_)
  );
  INV_X1 _34681_ (
    .A(_26543_),
    .ZN(_26544_)
  );
  AND2_X1 _34682_ (
    .A1(_22147_),
    .A2(_26544_),
    .ZN(_26545_)
  );
  AND2_X1 _34683_ (
    .A1(_26542_),
    .A2(_26545_),
    .ZN(_26546_)
  );
  INV_X1 _34684_ (
    .A(_26546_),
    .ZN(_26547_)
  );
  AND2_X1 _34685_ (
    .A1(\cpuregs[19] [21]),
    .A2(_22149_),
    .ZN(_26548_)
  );
  INV_X1 _34686_ (
    .A(_26548_),
    .ZN(_26549_)
  );
  AND2_X1 _34687_ (
    .A1(\cpuregs[23] [21]),
    .A2(_00008_[2]),
    .ZN(_26550_)
  );
  INV_X1 _34688_ (
    .A(_26550_),
    .ZN(_26551_)
  );
  AND2_X1 _34689_ (
    .A1(_00008_[0]),
    .A2(_26551_),
    .ZN(_26552_)
  );
  AND2_X1 _34690_ (
    .A1(_26549_),
    .A2(_26552_),
    .ZN(_26553_)
  );
  INV_X1 _34691_ (
    .A(_26553_),
    .ZN(_26554_)
  );
  AND2_X1 _34692_ (
    .A1(_26547_),
    .A2(_26554_),
    .ZN(_26555_)
  );
  INV_X1 _34693_ (
    .A(_26555_),
    .ZN(_26556_)
  );
  AND2_X1 _34694_ (
    .A1(_22150_),
    .A2(_26556_),
    .ZN(_26557_)
  );
  INV_X1 _34695_ (
    .A(_26557_),
    .ZN(_26558_)
  );
  AND2_X1 _34696_ (
    .A1(_26540_),
    .A2(_26558_),
    .ZN(_26559_)
  );
  AND2_X1 _34697_ (
    .A1(_00008_[1]),
    .A2(_26559_),
    .ZN(_26560_)
  );
  INV_X1 _34698_ (
    .A(_26560_),
    .ZN(_26561_)
  );
  AND2_X1 _34699_ (
    .A1(_22148_),
    .A2(_26522_),
    .ZN(_26562_)
  );
  AND2_X1 _34700_ (
    .A1(_26503_),
    .A2(_26562_),
    .ZN(_26563_)
  );
  INV_X1 _34701_ (
    .A(_26563_),
    .ZN(_26564_)
  );
  AND2_X1 _34702_ (
    .A1(_00008_[4]),
    .A2(_26564_),
    .ZN(_26565_)
  );
  AND2_X1 _34703_ (
    .A1(_26561_),
    .A2(_26565_),
    .ZN(_26566_)
  );
  INV_X1 _34704_ (
    .A(_26566_),
    .ZN(_26567_)
  );
  AND2_X1 _34705_ (
    .A1(\cpuregs[9] [21]),
    .A2(_22149_),
    .ZN(_26568_)
  );
  INV_X1 _34706_ (
    .A(_26568_),
    .ZN(_26569_)
  );
  AND2_X1 _34707_ (
    .A1(\cpuregs[13] [21]),
    .A2(_00008_[2]),
    .ZN(_26570_)
  );
  INV_X1 _34708_ (
    .A(_26570_),
    .ZN(_26571_)
  );
  AND2_X1 _34709_ (
    .A1(_22148_),
    .A2(_26571_),
    .ZN(_26572_)
  );
  AND2_X1 _34710_ (
    .A1(_26569_),
    .A2(_26572_),
    .ZN(_26573_)
  );
  INV_X1 _34711_ (
    .A(_26573_),
    .ZN(_26574_)
  );
  AND2_X1 _34712_ (
    .A1(\cpuregs[15] [21]),
    .A2(_00008_[2]),
    .ZN(_26575_)
  );
  INV_X1 _34713_ (
    .A(_26575_),
    .ZN(_26576_)
  );
  AND2_X1 _34714_ (
    .A1(\cpuregs[11] [21]),
    .A2(_22149_),
    .ZN(_26577_)
  );
  INV_X1 _34715_ (
    .A(_26577_),
    .ZN(_26578_)
  );
  AND2_X1 _34716_ (
    .A1(_00008_[1]),
    .A2(_26578_),
    .ZN(_26579_)
  );
  AND2_X1 _34717_ (
    .A1(_26576_),
    .A2(_26579_),
    .ZN(_26580_)
  );
  INV_X1 _34718_ (
    .A(_26580_),
    .ZN(_26581_)
  );
  AND2_X1 _34719_ (
    .A1(_26574_),
    .A2(_26581_),
    .ZN(_26582_)
  );
  INV_X1 _34720_ (
    .A(_26582_),
    .ZN(_26583_)
  );
  AND2_X1 _34721_ (
    .A1(_00008_[0]),
    .A2(_26583_),
    .ZN(_26584_)
  );
  INV_X1 _34722_ (
    .A(_26584_),
    .ZN(_26585_)
  );
  AND2_X1 _34723_ (
    .A1(\cpuregs[8] [21]),
    .A2(_22149_),
    .ZN(_26586_)
  );
  INV_X1 _34724_ (
    .A(_26586_),
    .ZN(_26587_)
  );
  AND2_X1 _34725_ (
    .A1(\cpuregs[12] [21]),
    .A2(_00008_[2]),
    .ZN(_26588_)
  );
  INV_X1 _34726_ (
    .A(_26588_),
    .ZN(_26589_)
  );
  AND2_X1 _34727_ (
    .A1(_22148_),
    .A2(_26589_),
    .ZN(_26590_)
  );
  AND2_X1 _34728_ (
    .A1(_26587_),
    .A2(_26590_),
    .ZN(_26591_)
  );
  INV_X1 _34729_ (
    .A(_26591_),
    .ZN(_26592_)
  );
  AND2_X1 _34730_ (
    .A1(\cpuregs[10] [21]),
    .A2(_22149_),
    .ZN(_26593_)
  );
  INV_X1 _34731_ (
    .A(_26593_),
    .ZN(_26594_)
  );
  AND2_X1 _34732_ (
    .A1(\cpuregs[14] [21]),
    .A2(_00008_[2]),
    .ZN(_26595_)
  );
  INV_X1 _34733_ (
    .A(_26595_),
    .ZN(_26596_)
  );
  AND2_X1 _34734_ (
    .A1(_00008_[1]),
    .A2(_26596_),
    .ZN(_26597_)
  );
  AND2_X1 _34735_ (
    .A1(_26594_),
    .A2(_26597_),
    .ZN(_26598_)
  );
  INV_X1 _34736_ (
    .A(_26598_),
    .ZN(_26599_)
  );
  AND2_X1 _34737_ (
    .A1(_26592_),
    .A2(_26599_),
    .ZN(_26600_)
  );
  INV_X1 _34738_ (
    .A(_26600_),
    .ZN(_26601_)
  );
  AND2_X1 _34739_ (
    .A1(_22147_),
    .A2(_26601_),
    .ZN(_26602_)
  );
  INV_X1 _34740_ (
    .A(_26602_),
    .ZN(_26603_)
  );
  AND2_X1 _34741_ (
    .A1(_26585_),
    .A2(_26603_),
    .ZN(_26604_)
  );
  INV_X1 _34742_ (
    .A(_26604_),
    .ZN(_26605_)
  );
  AND2_X1 _34743_ (
    .A1(_00008_[3]),
    .A2(_26605_),
    .ZN(_26606_)
  );
  INV_X1 _34744_ (
    .A(_26606_),
    .ZN(_26607_)
  );
  AND2_X1 _34745_ (
    .A1(_21749_),
    .A2(_00008_[2]),
    .ZN(_26608_)
  );
  INV_X1 _34746_ (
    .A(_26608_),
    .ZN(_26609_)
  );
  AND2_X1 _34747_ (
    .A1(_21529_),
    .A2(_22149_),
    .ZN(_26610_)
  );
  INV_X1 _34748_ (
    .A(_26610_),
    .ZN(_26611_)
  );
  AND2_X1 _34749_ (
    .A1(_00008_[0]),
    .A2(_26611_),
    .ZN(_26612_)
  );
  AND2_X1 _34750_ (
    .A1(_26609_),
    .A2(_26612_),
    .ZN(_26613_)
  );
  INV_X1 _34751_ (
    .A(_26613_),
    .ZN(_26614_)
  );
  AND2_X1 _34752_ (
    .A1(_21970_),
    .A2(_22149_),
    .ZN(_26615_)
  );
  INV_X1 _34753_ (
    .A(_26615_),
    .ZN(_26616_)
  );
  AND2_X1 _34754_ (
    .A1(_21686_),
    .A2(_00008_[2]),
    .ZN(_26617_)
  );
  INV_X1 _34755_ (
    .A(_26617_),
    .ZN(_26618_)
  );
  AND2_X1 _34756_ (
    .A1(_26616_),
    .A2(_26618_),
    .ZN(_26619_)
  );
  AND2_X1 _34757_ (
    .A1(_22147_),
    .A2(_26619_),
    .ZN(_26620_)
  );
  INV_X1 _34758_ (
    .A(_26620_),
    .ZN(_26621_)
  );
  AND2_X1 _34759_ (
    .A1(_26614_),
    .A2(_26621_),
    .ZN(_26622_)
  );
  AND2_X1 _34760_ (
    .A1(_22148_),
    .A2(_26622_),
    .ZN(_26623_)
  );
  INV_X1 _34761_ (
    .A(_26623_),
    .ZN(_26624_)
  );
  AND2_X1 _34762_ (
    .A1(_21796_),
    .A2(_00008_[2]),
    .ZN(_26625_)
  );
  INV_X1 _34763_ (
    .A(_26625_),
    .ZN(_26626_)
  );
  AND2_X1 _34764_ (
    .A1(_21504_),
    .A2(_22149_),
    .ZN(_26627_)
  );
  INV_X1 _34765_ (
    .A(_26627_),
    .ZN(_26628_)
  );
  AND2_X1 _34766_ (
    .A1(_00008_[0]),
    .A2(_26628_),
    .ZN(_26629_)
  );
  AND2_X1 _34767_ (
    .A1(_26626_),
    .A2(_26629_),
    .ZN(_26630_)
  );
  INV_X1 _34768_ (
    .A(_26630_),
    .ZN(_26631_)
  );
  AND2_X1 _34769_ (
    .A1(_21557_),
    .A2(_22149_),
    .ZN(_26632_)
  );
  INV_X1 _34770_ (
    .A(_26632_),
    .ZN(_26633_)
  );
  AND2_X1 _34771_ (
    .A1(_21823_),
    .A2(_00008_[2]),
    .ZN(_26634_)
  );
  INV_X1 _34772_ (
    .A(_26634_),
    .ZN(_26635_)
  );
  AND2_X1 _34773_ (
    .A1(_26633_),
    .A2(_26635_),
    .ZN(_26636_)
  );
  AND2_X1 _34774_ (
    .A1(_22147_),
    .A2(_26636_),
    .ZN(_26637_)
  );
  INV_X1 _34775_ (
    .A(_26637_),
    .ZN(_26638_)
  );
  AND2_X1 _34776_ (
    .A1(_26631_),
    .A2(_26638_),
    .ZN(_26639_)
  );
  AND2_X1 _34777_ (
    .A1(_00008_[1]),
    .A2(_26639_),
    .ZN(_26640_)
  );
  INV_X1 _34778_ (
    .A(_26640_),
    .ZN(_26641_)
  );
  AND2_X1 _34779_ (
    .A1(_26624_),
    .A2(_26641_),
    .ZN(_26642_)
  );
  INV_X1 _34780_ (
    .A(_26642_),
    .ZN(_26643_)
  );
  AND2_X1 _34781_ (
    .A1(_22150_),
    .A2(_26643_),
    .ZN(_26644_)
  );
  INV_X1 _34782_ (
    .A(_26644_),
    .ZN(_26645_)
  );
  AND2_X1 _34783_ (
    .A1(_26607_),
    .A2(_26645_),
    .ZN(_26646_)
  );
  INV_X1 _34784_ (
    .A(_26646_),
    .ZN(_26647_)
  );
  AND2_X1 _34785_ (
    .A1(_22151_),
    .A2(_26647_),
    .ZN(_26648_)
  );
  INV_X1 _34786_ (
    .A(_26648_),
    .ZN(_26649_)
  );
  AND2_X1 _34787_ (
    .A1(_22546_),
    .A2(_26567_),
    .ZN(_26650_)
  );
  AND2_X1 _34788_ (
    .A1(_26649_),
    .A2(_26650_),
    .ZN(_26651_)
  );
  INV_X1 _34789_ (
    .A(_26651_),
    .ZN(_26652_)
  );
  AND2_X1 _34790_ (
    .A1(_26485_),
    .A2(_26652_),
    .ZN(_26653_)
  );
  INV_X1 _34791_ (
    .A(_26653_),
    .ZN(_26654_)
  );
  AND2_X1 _34792_ (
    .A1(_22271_),
    .A2(_26654_),
    .ZN(_26655_)
  );
  INV_X1 _34793_ (
    .A(_26655_),
    .ZN(_26656_)
  );
  AND2_X1 _34794_ (
    .A1(reg_op1[20]),
    .A2(_22285_),
    .ZN(_26657_)
  );
  INV_X1 _34795_ (
    .A(_26657_),
    .ZN(_26658_)
  );
  AND2_X1 _34796_ (
    .A1(_26039_),
    .A2(_26658_),
    .ZN(_26659_)
  );
  AND2_X1 _34797_ (
    .A1(reg_op1[25]),
    .A2(_22290_),
    .ZN(_26660_)
  );
  INV_X1 _34798_ (
    .A(_26660_),
    .ZN(_26661_)
  );
  AND2_X1 _34799_ (
    .A1(_26036_),
    .A2(_26661_),
    .ZN(_26662_)
  );
  AND2_X1 _34800_ (
    .A1(_26464_),
    .A2(_26479_),
    .ZN(_26663_)
  );
  INV_X1 _34801_ (
    .A(_26663_),
    .ZN(_26664_)
  );
  AND2_X1 _34802_ (
    .A1(_26455_),
    .A2(_26479_),
    .ZN(_26665_)
  );
  INV_X1 _34803_ (
    .A(_26665_),
    .ZN(_26666_)
  );
  AND2_X1 _34804_ (
    .A1(_22559_),
    .A2(_26666_),
    .ZN(_26667_)
  );
  AND2_X1 _34805_ (
    .A1(_26664_),
    .A2(_26667_),
    .ZN(_26668_)
  );
  AND2_X1 _34806_ (
    .A1(_26483_),
    .A2(_26668_),
    .ZN(_26669_)
  );
  INV_X1 _34807_ (
    .A(_26669_),
    .ZN(_26670_)
  );
  AND2_X1 _34808_ (
    .A1(_22573_),
    .A2(_26662_),
    .ZN(_26671_)
  );
  INV_X1 _34809_ (
    .A(_26671_),
    .ZN(_26672_)
  );
  AND2_X1 _34810_ (
    .A1(_22572_),
    .A2(_26659_),
    .ZN(_26673_)
  );
  INV_X1 _34811_ (
    .A(_26673_),
    .ZN(_26674_)
  );
  AND2_X1 _34812_ (
    .A1(_22295_),
    .A2(_26672_),
    .ZN(_26675_)
  );
  AND2_X1 _34813_ (
    .A1(_26674_),
    .A2(_26675_),
    .ZN(_26676_)
  );
  INV_X1 _34814_ (
    .A(_26676_),
    .ZN(_26677_)
  );
  AND2_X1 _34815_ (
    .A1(_26656_),
    .A2(_26677_),
    .ZN(_26678_)
  );
  AND2_X1 _34816_ (
    .A1(_26670_),
    .A2(_26678_),
    .ZN(_26679_)
  );
  AND2_X1 _34817_ (
    .A1(_22333_),
    .A2(_26679_),
    .ZN(_26680_)
  );
  INV_X1 _34818_ (
    .A(_26680_),
    .ZN(_26681_)
  );
  AND2_X1 _34819_ (
    .A1(_26474_),
    .A2(_26681_),
    .ZN(_00078_)
  );
  AND2_X1 _34820_ (
    .A1(_21189_),
    .A2(_22334_),
    .ZN(_26682_)
  );
  INV_X1 _34821_ (
    .A(_26682_),
    .ZN(_26683_)
  );
  AND2_X1 _34822_ (
    .A1(reg_pc[22]),
    .A2(_22335_),
    .ZN(_26684_)
  );
  INV_X1 _34823_ (
    .A(_26684_),
    .ZN(_26685_)
  );
  AND2_X1 _34824_ (
    .A1(\cpuregs[12] [22]),
    .A2(_00008_[2]),
    .ZN(_26686_)
  );
  INV_X1 _34825_ (
    .A(_26686_),
    .ZN(_26687_)
  );
  AND2_X1 _34826_ (
    .A1(\cpuregs[8] [22]),
    .A2(_22149_),
    .ZN(_26688_)
  );
  INV_X1 _34827_ (
    .A(_26688_),
    .ZN(_26689_)
  );
  AND2_X1 _34828_ (
    .A1(_26687_),
    .A2(_26689_),
    .ZN(_26690_)
  );
  INV_X1 _34829_ (
    .A(_26690_),
    .ZN(_26691_)
  );
  AND2_X1 _34830_ (
    .A1(_22147_),
    .A2(_26691_),
    .ZN(_26692_)
  );
  INV_X1 _34831_ (
    .A(_26692_),
    .ZN(_26693_)
  );
  AND2_X1 _34832_ (
    .A1(\cpuregs[9] [22]),
    .A2(_22149_),
    .ZN(_26694_)
  );
  INV_X1 _34833_ (
    .A(_26694_),
    .ZN(_26695_)
  );
  AND2_X1 _34834_ (
    .A1(\cpuregs[13] [22]),
    .A2(_00008_[2]),
    .ZN(_26696_)
  );
  INV_X1 _34835_ (
    .A(_26696_),
    .ZN(_26697_)
  );
  AND2_X1 _34836_ (
    .A1(_26695_),
    .A2(_26697_),
    .ZN(_26698_)
  );
  INV_X1 _34837_ (
    .A(_26698_),
    .ZN(_26699_)
  );
  AND2_X1 _34838_ (
    .A1(_00008_[0]),
    .A2(_26699_),
    .ZN(_26700_)
  );
  INV_X1 _34839_ (
    .A(_26700_),
    .ZN(_26701_)
  );
  AND2_X1 _34840_ (
    .A1(_26693_),
    .A2(_26701_),
    .ZN(_26702_)
  );
  AND2_X1 _34841_ (
    .A1(\cpuregs[5] [22]),
    .A2(_00008_[2]),
    .ZN(_26703_)
  );
  INV_X1 _34842_ (
    .A(_26703_),
    .ZN(_26704_)
  );
  AND2_X1 _34843_ (
    .A1(\cpuregs[1] [22]),
    .A2(_22149_),
    .ZN(_26705_)
  );
  INV_X1 _34844_ (
    .A(_26705_),
    .ZN(_26706_)
  );
  AND2_X1 _34845_ (
    .A1(_26704_),
    .A2(_26706_),
    .ZN(_26707_)
  );
  AND2_X1 _34846_ (
    .A1(\cpuregs[4] [22]),
    .A2(_00008_[2]),
    .ZN(_26708_)
  );
  INV_X1 _34847_ (
    .A(_26708_),
    .ZN(_26709_)
  );
  AND2_X1 _34848_ (
    .A1(\cpuregs[0] [22]),
    .A2(_22149_),
    .ZN(_26710_)
  );
  INV_X1 _34849_ (
    .A(_26710_),
    .ZN(_26711_)
  );
  AND2_X1 _34850_ (
    .A1(_26709_),
    .A2(_26711_),
    .ZN(_26712_)
  );
  AND2_X1 _34851_ (
    .A1(_00008_[0]),
    .A2(_26707_),
    .ZN(_26713_)
  );
  INV_X1 _34852_ (
    .A(_26713_),
    .ZN(_26714_)
  );
  AND2_X1 _34853_ (
    .A1(_22147_),
    .A2(_26712_),
    .ZN(_26715_)
  );
  INV_X1 _34854_ (
    .A(_26715_),
    .ZN(_26716_)
  );
  AND2_X1 _34855_ (
    .A1(_26714_),
    .A2(_26716_),
    .ZN(_26717_)
  );
  INV_X1 _34856_ (
    .A(_26717_),
    .ZN(_26718_)
  );
  AND2_X1 _34857_ (
    .A1(_00008_[3]),
    .A2(_26702_),
    .ZN(_26719_)
  );
  INV_X1 _34858_ (
    .A(_26719_),
    .ZN(_26720_)
  );
  AND2_X1 _34859_ (
    .A1(_22150_),
    .A2(_26718_),
    .ZN(_26721_)
  );
  INV_X1 _34860_ (
    .A(_26721_),
    .ZN(_26722_)
  );
  AND2_X1 _34861_ (
    .A1(_26720_),
    .A2(_26722_),
    .ZN(_26723_)
  );
  AND2_X1 _34862_ (
    .A1(_22148_),
    .A2(_26723_),
    .ZN(_26724_)
  );
  INV_X1 _34863_ (
    .A(_26724_),
    .ZN(_26725_)
  );
  AND2_X1 _34864_ (
    .A1(\cpuregs[11] [22]),
    .A2(_22149_),
    .ZN(_26726_)
  );
  INV_X1 _34865_ (
    .A(_26726_),
    .ZN(_26727_)
  );
  AND2_X1 _34866_ (
    .A1(\cpuregs[15] [22]),
    .A2(_00008_[2]),
    .ZN(_26728_)
  );
  INV_X1 _34867_ (
    .A(_26728_),
    .ZN(_26729_)
  );
  AND2_X1 _34868_ (
    .A1(_26727_),
    .A2(_26729_),
    .ZN(_26730_)
  );
  INV_X1 _34869_ (
    .A(_26730_),
    .ZN(_26731_)
  );
  AND2_X1 _34870_ (
    .A1(_00008_[0]),
    .A2(_26731_),
    .ZN(_26732_)
  );
  INV_X1 _34871_ (
    .A(_26732_),
    .ZN(_26733_)
  );
  AND2_X1 _34872_ (
    .A1(\cpuregs[14] [22]),
    .A2(_00008_[2]),
    .ZN(_26734_)
  );
  INV_X1 _34873_ (
    .A(_26734_),
    .ZN(_26735_)
  );
  AND2_X1 _34874_ (
    .A1(\cpuregs[10] [22]),
    .A2(_22149_),
    .ZN(_26736_)
  );
  INV_X1 _34875_ (
    .A(_26736_),
    .ZN(_26737_)
  );
  AND2_X1 _34876_ (
    .A1(_26735_),
    .A2(_26737_),
    .ZN(_26738_)
  );
  INV_X1 _34877_ (
    .A(_26738_),
    .ZN(_26739_)
  );
  AND2_X1 _34878_ (
    .A1(_22147_),
    .A2(_26739_),
    .ZN(_26740_)
  );
  INV_X1 _34879_ (
    .A(_26740_),
    .ZN(_26741_)
  );
  AND2_X1 _34880_ (
    .A1(_26733_),
    .A2(_26741_),
    .ZN(_26742_)
  );
  AND2_X1 _34881_ (
    .A1(\cpuregs[7] [22]),
    .A2(_00008_[2]),
    .ZN(_26743_)
  );
  INV_X1 _34882_ (
    .A(_26743_),
    .ZN(_26744_)
  );
  AND2_X1 _34883_ (
    .A1(\cpuregs[3] [22]),
    .A2(_22149_),
    .ZN(_26745_)
  );
  INV_X1 _34884_ (
    .A(_26745_),
    .ZN(_26746_)
  );
  AND2_X1 _34885_ (
    .A1(_26744_),
    .A2(_26746_),
    .ZN(_26747_)
  );
  AND2_X1 _34886_ (
    .A1(\cpuregs[6] [22]),
    .A2(_00008_[2]),
    .ZN(_26748_)
  );
  INV_X1 _34887_ (
    .A(_26748_),
    .ZN(_26749_)
  );
  AND2_X1 _34888_ (
    .A1(\cpuregs[2] [22]),
    .A2(_22149_),
    .ZN(_26750_)
  );
  INV_X1 _34889_ (
    .A(_26750_),
    .ZN(_26751_)
  );
  AND2_X1 _34890_ (
    .A1(_26749_),
    .A2(_26751_),
    .ZN(_26752_)
  );
  AND2_X1 _34891_ (
    .A1(_00008_[0]),
    .A2(_26747_),
    .ZN(_26753_)
  );
  INV_X1 _34892_ (
    .A(_26753_),
    .ZN(_26754_)
  );
  AND2_X1 _34893_ (
    .A1(_22147_),
    .A2(_26752_),
    .ZN(_26755_)
  );
  INV_X1 _34894_ (
    .A(_26755_),
    .ZN(_26756_)
  );
  AND2_X1 _34895_ (
    .A1(_26754_),
    .A2(_26756_),
    .ZN(_26757_)
  );
  INV_X1 _34896_ (
    .A(_26757_),
    .ZN(_26758_)
  );
  AND2_X1 _34897_ (
    .A1(_00008_[3]),
    .A2(_26742_),
    .ZN(_26759_)
  );
  INV_X1 _34898_ (
    .A(_26759_),
    .ZN(_26760_)
  );
  AND2_X1 _34899_ (
    .A1(_22150_),
    .A2(_26758_),
    .ZN(_26761_)
  );
  INV_X1 _34900_ (
    .A(_26761_),
    .ZN(_26762_)
  );
  AND2_X1 _34901_ (
    .A1(_00008_[1]),
    .A2(_26762_),
    .ZN(_26763_)
  );
  AND2_X1 _34902_ (
    .A1(_26760_),
    .A2(_26763_),
    .ZN(_26764_)
  );
  INV_X1 _34903_ (
    .A(_26764_),
    .ZN(_26765_)
  );
  AND2_X1 _34904_ (
    .A1(_26725_),
    .A2(_26765_),
    .ZN(_26766_)
  );
  AND2_X1 _34905_ (
    .A1(_22151_),
    .A2(_26766_),
    .ZN(_26767_)
  );
  INV_X1 _34906_ (
    .A(_26767_),
    .ZN(_26768_)
  );
  AND2_X1 _34907_ (
    .A1(\cpuregs[26] [22]),
    .A2(_22149_),
    .ZN(_26769_)
  );
  INV_X1 _34908_ (
    .A(_26769_),
    .ZN(_26770_)
  );
  AND2_X1 _34909_ (
    .A1(\cpuregs[30] [22]),
    .A2(_00008_[2]),
    .ZN(_26771_)
  );
  INV_X1 _34910_ (
    .A(_26771_),
    .ZN(_26772_)
  );
  AND2_X1 _34911_ (
    .A1(_22147_),
    .A2(_26772_),
    .ZN(_26773_)
  );
  AND2_X1 _34912_ (
    .A1(_26770_),
    .A2(_26773_),
    .ZN(_26774_)
  );
  INV_X1 _34913_ (
    .A(_26774_),
    .ZN(_26775_)
  );
  AND2_X1 _34914_ (
    .A1(\cpuregs[31] [22]),
    .A2(_00008_[2]),
    .ZN(_26776_)
  );
  INV_X1 _34915_ (
    .A(_26776_),
    .ZN(_26777_)
  );
  AND2_X1 _34916_ (
    .A1(\cpuregs[27] [22]),
    .A2(_22149_),
    .ZN(_26778_)
  );
  INV_X1 _34917_ (
    .A(_26778_),
    .ZN(_26779_)
  );
  AND2_X1 _34918_ (
    .A1(_00008_[0]),
    .A2(_26779_),
    .ZN(_26780_)
  );
  AND2_X1 _34919_ (
    .A1(_26777_),
    .A2(_26780_),
    .ZN(_26781_)
  );
  INV_X1 _34920_ (
    .A(_26781_),
    .ZN(_26782_)
  );
  AND2_X1 _34921_ (
    .A1(_26775_),
    .A2(_26782_),
    .ZN(_26783_)
  );
  INV_X1 _34922_ (
    .A(_26783_),
    .ZN(_26784_)
  );
  AND2_X1 _34923_ (
    .A1(_00008_[3]),
    .A2(_26784_),
    .ZN(_26785_)
  );
  INV_X1 _34924_ (
    .A(_26785_),
    .ZN(_26786_)
  );
  AND2_X1 _34925_ (
    .A1(\cpuregs[18] [22]),
    .A2(_22149_),
    .ZN(_26787_)
  );
  INV_X1 _34926_ (
    .A(_26787_),
    .ZN(_26788_)
  );
  AND2_X1 _34927_ (
    .A1(\cpuregs[22] [22]),
    .A2(_00008_[2]),
    .ZN(_26789_)
  );
  INV_X1 _34928_ (
    .A(_26789_),
    .ZN(_26790_)
  );
  AND2_X1 _34929_ (
    .A1(_22147_),
    .A2(_26790_),
    .ZN(_26791_)
  );
  AND2_X1 _34930_ (
    .A1(_26788_),
    .A2(_26791_),
    .ZN(_26792_)
  );
  INV_X1 _34931_ (
    .A(_26792_),
    .ZN(_26793_)
  );
  AND2_X1 _34932_ (
    .A1(\cpuregs[19] [22]),
    .A2(_22149_),
    .ZN(_26794_)
  );
  INV_X1 _34933_ (
    .A(_26794_),
    .ZN(_26795_)
  );
  AND2_X1 _34934_ (
    .A1(\cpuregs[23] [22]),
    .A2(_00008_[2]),
    .ZN(_26796_)
  );
  INV_X1 _34935_ (
    .A(_26796_),
    .ZN(_26797_)
  );
  AND2_X1 _34936_ (
    .A1(_00008_[0]),
    .A2(_26797_),
    .ZN(_26798_)
  );
  AND2_X1 _34937_ (
    .A1(_26795_),
    .A2(_26798_),
    .ZN(_26799_)
  );
  INV_X1 _34938_ (
    .A(_26799_),
    .ZN(_26800_)
  );
  AND2_X1 _34939_ (
    .A1(_26793_),
    .A2(_26800_),
    .ZN(_26801_)
  );
  INV_X1 _34940_ (
    .A(_26801_),
    .ZN(_26802_)
  );
  AND2_X1 _34941_ (
    .A1(_22150_),
    .A2(_26802_),
    .ZN(_26803_)
  );
  INV_X1 _34942_ (
    .A(_26803_),
    .ZN(_26804_)
  );
  AND2_X1 _34943_ (
    .A1(\cpuregs[16] [22]),
    .A2(_22149_),
    .ZN(_26805_)
  );
  INV_X1 _34944_ (
    .A(_26805_),
    .ZN(_26806_)
  );
  AND2_X1 _34945_ (
    .A1(\cpuregs[20] [22]),
    .A2(_00008_[2]),
    .ZN(_26807_)
  );
  INV_X1 _34946_ (
    .A(_26807_),
    .ZN(_26808_)
  );
  AND2_X1 _34947_ (
    .A1(_22147_),
    .A2(_26808_),
    .ZN(_26809_)
  );
  AND2_X1 _34948_ (
    .A1(_26806_),
    .A2(_26809_),
    .ZN(_26810_)
  );
  INV_X1 _34949_ (
    .A(_26810_),
    .ZN(_26811_)
  );
  AND2_X1 _34950_ (
    .A1(\cpuregs[17] [22]),
    .A2(_22149_),
    .ZN(_26812_)
  );
  INV_X1 _34951_ (
    .A(_26812_),
    .ZN(_26813_)
  );
  AND2_X1 _34952_ (
    .A1(\cpuregs[21] [22]),
    .A2(_00008_[2]),
    .ZN(_26814_)
  );
  INV_X1 _34953_ (
    .A(_26814_),
    .ZN(_26815_)
  );
  AND2_X1 _34954_ (
    .A1(_00008_[0]),
    .A2(_26815_),
    .ZN(_26816_)
  );
  AND2_X1 _34955_ (
    .A1(_26813_),
    .A2(_26816_),
    .ZN(_26817_)
  );
  INV_X1 _34956_ (
    .A(_26817_),
    .ZN(_26818_)
  );
  AND2_X1 _34957_ (
    .A1(_26811_),
    .A2(_26818_),
    .ZN(_26819_)
  );
  INV_X1 _34958_ (
    .A(_26819_),
    .ZN(_26820_)
  );
  AND2_X1 _34959_ (
    .A1(_22150_),
    .A2(_26820_),
    .ZN(_26821_)
  );
  INV_X1 _34960_ (
    .A(_26821_),
    .ZN(_26822_)
  );
  AND2_X1 _34961_ (
    .A1(\cpuregs[24] [22]),
    .A2(_22149_),
    .ZN(_26823_)
  );
  INV_X1 _34962_ (
    .A(_26823_),
    .ZN(_26824_)
  );
  AND2_X1 _34963_ (
    .A1(\cpuregs[28] [22]),
    .A2(_00008_[2]),
    .ZN(_26825_)
  );
  INV_X1 _34964_ (
    .A(_26825_),
    .ZN(_26826_)
  );
  AND2_X1 _34965_ (
    .A1(_22147_),
    .A2(_26826_),
    .ZN(_26827_)
  );
  AND2_X1 _34966_ (
    .A1(_26824_),
    .A2(_26827_),
    .ZN(_26828_)
  );
  INV_X1 _34967_ (
    .A(_26828_),
    .ZN(_26829_)
  );
  AND2_X1 _34968_ (
    .A1(\cpuregs[25] [22]),
    .A2(_22149_),
    .ZN(_26830_)
  );
  INV_X1 _34969_ (
    .A(_26830_),
    .ZN(_26831_)
  );
  AND2_X1 _34970_ (
    .A1(\cpuregs[29] [22]),
    .A2(_00008_[2]),
    .ZN(_26832_)
  );
  INV_X1 _34971_ (
    .A(_26832_),
    .ZN(_26833_)
  );
  AND2_X1 _34972_ (
    .A1(_00008_[0]),
    .A2(_26833_),
    .ZN(_26834_)
  );
  AND2_X1 _34973_ (
    .A1(_26831_),
    .A2(_26834_),
    .ZN(_26835_)
  );
  INV_X1 _34974_ (
    .A(_26835_),
    .ZN(_26836_)
  );
  AND2_X1 _34975_ (
    .A1(_26829_),
    .A2(_26836_),
    .ZN(_26837_)
  );
  INV_X1 _34976_ (
    .A(_26837_),
    .ZN(_26838_)
  );
  AND2_X1 _34977_ (
    .A1(_00008_[3]),
    .A2(_26838_),
    .ZN(_26839_)
  );
  INV_X1 _34978_ (
    .A(_26839_),
    .ZN(_26840_)
  );
  AND2_X1 _34979_ (
    .A1(_26822_),
    .A2(_26840_),
    .ZN(_26841_)
  );
  AND2_X1 _34980_ (
    .A1(_00008_[1]),
    .A2(_26804_),
    .ZN(_26842_)
  );
  AND2_X1 _34981_ (
    .A1(_26786_),
    .A2(_26842_),
    .ZN(_26843_)
  );
  INV_X1 _34982_ (
    .A(_26843_),
    .ZN(_26844_)
  );
  AND2_X1 _34983_ (
    .A1(_22148_),
    .A2(_26841_),
    .ZN(_26845_)
  );
  INV_X1 _34984_ (
    .A(_26845_),
    .ZN(_26846_)
  );
  AND2_X1 _34985_ (
    .A1(_00008_[4]),
    .A2(_26844_),
    .ZN(_26847_)
  );
  AND2_X1 _34986_ (
    .A1(_26846_),
    .A2(_26847_),
    .ZN(_26848_)
  );
  INV_X1 _34987_ (
    .A(_26848_),
    .ZN(_26849_)
  );
  AND2_X1 _34988_ (
    .A1(_22546_),
    .A2(_26849_),
    .ZN(_26850_)
  );
  AND2_X1 _34989_ (
    .A1(_26768_),
    .A2(_26850_),
    .ZN(_26851_)
  );
  INV_X1 _34990_ (
    .A(_26851_),
    .ZN(_26852_)
  );
  AND2_X1 _34991_ (
    .A1(_26685_),
    .A2(_26852_),
    .ZN(_26853_)
  );
  INV_X1 _34992_ (
    .A(_26853_),
    .ZN(_26854_)
  );
  AND2_X1 _34993_ (
    .A1(_22271_),
    .A2(_26854_),
    .ZN(_26855_)
  );
  INV_X1 _34994_ (
    .A(_26855_),
    .ZN(_26856_)
  );
  AND2_X1 _34995_ (
    .A1(reg_op1[21]),
    .A2(_22285_),
    .ZN(_26857_)
  );
  INV_X1 _34996_ (
    .A(_26857_),
    .ZN(_26858_)
  );
  AND2_X1 _34997_ (
    .A1(_26240_),
    .A2(_26858_),
    .ZN(_26859_)
  );
  AND2_X1 _34998_ (
    .A1(reg_op1[26]),
    .A2(_22290_),
    .ZN(_26860_)
  );
  INV_X1 _34999_ (
    .A(_26860_),
    .ZN(_26861_)
  );
  AND2_X1 _35000_ (
    .A1(_26237_),
    .A2(_26861_),
    .ZN(_26862_)
  );
  AND2_X1 _35001_ (
    .A1(_22572_),
    .A2(_26859_),
    .ZN(_26863_)
  );
  INV_X1 _35002_ (
    .A(_26863_),
    .ZN(_26864_)
  );
  AND2_X1 _35003_ (
    .A1(_22573_),
    .A2(_26862_),
    .ZN(_26865_)
  );
  INV_X1 _35004_ (
    .A(_26865_),
    .ZN(_26866_)
  );
  AND2_X1 _35005_ (
    .A1(_22295_),
    .A2(_26866_),
    .ZN(_26867_)
  );
  AND2_X1 _35006_ (
    .A1(_26864_),
    .A2(_26867_),
    .ZN(_26868_)
  );
  INV_X1 _35007_ (
    .A(_26868_),
    .ZN(_26869_)
  );
  AND2_X1 _35008_ (
    .A1(_22333_),
    .A2(_26869_),
    .ZN(_26870_)
  );
  AND2_X1 _35009_ (
    .A1(_26856_),
    .A2(_26870_),
    .ZN(_26871_)
  );
  AND2_X1 _35010_ (
    .A1(reg_op1[22]),
    .A2(decoded_imm[22]),
    .ZN(_26872_)
  );
  INV_X1 _35011_ (
    .A(_26872_),
    .ZN(_26873_)
  );
  AND2_X1 _35012_ (
    .A1(_21189_),
    .A2(_21987_),
    .ZN(_26874_)
  );
  INV_X1 _35013_ (
    .A(_26874_),
    .ZN(_26875_)
  );
  AND2_X1 _35014_ (
    .A1(_26873_),
    .A2(_26875_),
    .ZN(_26876_)
  );
  INV_X1 _35015_ (
    .A(_26876_),
    .ZN(_26877_)
  );
  AND2_X1 _35016_ (
    .A1(_26476_),
    .A2(_26666_),
    .ZN(_26878_)
  );
  AND2_X1 _35017_ (
    .A1(_26664_),
    .A2(_26878_),
    .ZN(_26879_)
  );
  INV_X1 _35018_ (
    .A(_26879_),
    .ZN(_26880_)
  );
  AND2_X1 _35019_ (
    .A1(_26876_),
    .A2(_26880_),
    .ZN(_26881_)
  );
  INV_X1 _35020_ (
    .A(_26881_),
    .ZN(_26882_)
  );
  AND2_X1 _35021_ (
    .A1(_26877_),
    .A2(_26879_),
    .ZN(_26883_)
  );
  INV_X1 _35022_ (
    .A(_26883_),
    .ZN(_26884_)
  );
  AND2_X1 _35023_ (
    .A1(_22559_),
    .A2(_26884_),
    .ZN(_26885_)
  );
  AND2_X1 _35024_ (
    .A1(_26882_),
    .A2(_26885_),
    .ZN(_26886_)
  );
  INV_X1 _35025_ (
    .A(_26886_),
    .ZN(_26887_)
  );
  AND2_X1 _35026_ (
    .A1(_26871_),
    .A2(_26887_),
    .ZN(_26888_)
  );
  INV_X1 _35027_ (
    .A(_26888_),
    .ZN(_26889_)
  );
  AND2_X1 _35028_ (
    .A1(_26683_),
    .A2(_26889_),
    .ZN(_00079_)
  );
  AND2_X1 _35029_ (
    .A1(_21190_),
    .A2(_22334_),
    .ZN(_26890_)
  );
  INV_X1 _35030_ (
    .A(_26890_),
    .ZN(_26891_)
  );
  AND2_X1 _35031_ (
    .A1(reg_op1[23]),
    .A2(decoded_imm[23]),
    .ZN(_26892_)
  );
  INV_X1 _35032_ (
    .A(_26892_),
    .ZN(_26893_)
  );
  AND2_X1 _35033_ (
    .A1(_21190_),
    .A2(_21986_),
    .ZN(_26894_)
  );
  INV_X1 _35034_ (
    .A(_26894_),
    .ZN(_26895_)
  );
  AND2_X1 _35035_ (
    .A1(_26893_),
    .A2(_26895_),
    .ZN(_26896_)
  );
  INV_X1 _35036_ (
    .A(_26896_),
    .ZN(_26897_)
  );
  AND2_X1 _35037_ (
    .A1(_26873_),
    .A2(_26882_),
    .ZN(_26898_)
  );
  INV_X1 _35038_ (
    .A(_26898_),
    .ZN(_26899_)
  );
  AND2_X1 _35039_ (
    .A1(_26897_),
    .A2(_26898_),
    .ZN(_26900_)
  );
  INV_X1 _35040_ (
    .A(_26900_),
    .ZN(_26901_)
  );
  AND2_X1 _35041_ (
    .A1(_26896_),
    .A2(_26899_),
    .ZN(_26902_)
  );
  INV_X1 _35042_ (
    .A(_26902_),
    .ZN(_26903_)
  );
  AND2_X1 _35043_ (
    .A1(_22559_),
    .A2(_26903_),
    .ZN(_26904_)
  );
  AND2_X1 _35044_ (
    .A1(_26901_),
    .A2(_26904_),
    .ZN(_26905_)
  );
  INV_X1 _35045_ (
    .A(_26905_),
    .ZN(_26906_)
  );
  AND2_X1 _35046_ (
    .A1(reg_pc[23]),
    .A2(_22335_),
    .ZN(_26907_)
  );
  INV_X1 _35047_ (
    .A(_26907_),
    .ZN(_26908_)
  );
  AND2_X1 _35048_ (
    .A1(_21710_),
    .A2(_22149_),
    .ZN(_26909_)
  );
  INV_X1 _35049_ (
    .A(_26909_),
    .ZN(_26910_)
  );
  AND2_X1 _35050_ (
    .A1(_21398_),
    .A2(_00008_[2]),
    .ZN(_26911_)
  );
  INV_X1 _35051_ (
    .A(_26911_),
    .ZN(_26912_)
  );
  AND2_X1 _35052_ (
    .A1(_26910_),
    .A2(_26912_),
    .ZN(_26913_)
  );
  AND2_X1 _35053_ (
    .A1(_22147_),
    .A2(_26913_),
    .ZN(_26914_)
  );
  INV_X1 _35054_ (
    .A(_26914_),
    .ZN(_26915_)
  );
  AND2_X1 _35055_ (
    .A1(_21405_),
    .A2(_00008_[2]),
    .ZN(_26916_)
  );
  INV_X1 _35056_ (
    .A(_26916_),
    .ZN(_26917_)
  );
  AND2_X1 _35057_ (
    .A1(_21587_),
    .A2(_22149_),
    .ZN(_26918_)
  );
  INV_X1 _35058_ (
    .A(_26918_),
    .ZN(_26919_)
  );
  AND2_X1 _35059_ (
    .A1(_00008_[0]),
    .A2(_26919_),
    .ZN(_26920_)
  );
  AND2_X1 _35060_ (
    .A1(_26917_),
    .A2(_26920_),
    .ZN(_26921_)
  );
  INV_X1 _35061_ (
    .A(_26921_),
    .ZN(_26922_)
  );
  AND2_X1 _35062_ (
    .A1(_26915_),
    .A2(_26922_),
    .ZN(_26923_)
  );
  AND2_X1 _35063_ (
    .A1(_00008_[1]),
    .A2(_26923_),
    .ZN(_26924_)
  );
  INV_X1 _35064_ (
    .A(_26924_),
    .ZN(_26925_)
  );
  AND2_X1 _35065_ (
    .A1(_21644_),
    .A2(_00008_[2]),
    .ZN(_26926_)
  );
  INV_X1 _35066_ (
    .A(_26926_),
    .ZN(_26927_)
  );
  AND2_X1 _35067_ (
    .A1(_21722_),
    .A2(_22149_),
    .ZN(_26928_)
  );
  INV_X1 _35068_ (
    .A(_26928_),
    .ZN(_26929_)
  );
  AND2_X1 _35069_ (
    .A1(_00008_[0]),
    .A2(_26929_),
    .ZN(_26930_)
  );
  AND2_X1 _35070_ (
    .A1(_26927_),
    .A2(_26930_),
    .ZN(_26931_)
  );
  INV_X1 _35071_ (
    .A(_26931_),
    .ZN(_26932_)
  );
  AND2_X1 _35072_ (
    .A1(_21729_),
    .A2(_22149_),
    .ZN(_26933_)
  );
  INV_X1 _35073_ (
    .A(_26933_),
    .ZN(_26934_)
  );
  AND2_X1 _35074_ (
    .A1(_21484_),
    .A2(_00008_[2]),
    .ZN(_26935_)
  );
  INV_X1 _35075_ (
    .A(_26935_),
    .ZN(_26936_)
  );
  AND2_X1 _35076_ (
    .A1(_26934_),
    .A2(_26936_),
    .ZN(_26937_)
  );
  AND2_X1 _35077_ (
    .A1(_22147_),
    .A2(_26937_),
    .ZN(_26938_)
  );
  INV_X1 _35078_ (
    .A(_26938_),
    .ZN(_26939_)
  );
  AND2_X1 _35079_ (
    .A1(_26932_),
    .A2(_26939_),
    .ZN(_26940_)
  );
  AND2_X1 _35080_ (
    .A1(_22148_),
    .A2(_26940_),
    .ZN(_26941_)
  );
  INV_X1 _35081_ (
    .A(_26941_),
    .ZN(_26942_)
  );
  AND2_X1 _35082_ (
    .A1(_26925_),
    .A2(_26942_),
    .ZN(_26943_)
  );
  AND2_X1 _35083_ (
    .A1(_22151_),
    .A2(_26943_),
    .ZN(_26944_)
  );
  INV_X1 _35084_ (
    .A(_26944_),
    .ZN(_26945_)
  );
  AND2_X1 _35085_ (
    .A1(_21578_),
    .A2(_22149_),
    .ZN(_26946_)
  );
  INV_X1 _35086_ (
    .A(_26946_),
    .ZN(_26947_)
  );
  AND2_X1 _35087_ (
    .A1(_21916_),
    .A2(_00008_[2]),
    .ZN(_26948_)
  );
  INV_X1 _35088_ (
    .A(_26948_),
    .ZN(_26949_)
  );
  AND2_X1 _35089_ (
    .A1(_26947_),
    .A2(_26949_),
    .ZN(_26950_)
  );
  AND2_X1 _35090_ (
    .A1(_22147_),
    .A2(_26950_),
    .ZN(_26951_)
  );
  INV_X1 _35091_ (
    .A(_26951_),
    .ZN(_26952_)
  );
  AND2_X1 _35092_ (
    .A1(_21900_),
    .A2(_00008_[2]),
    .ZN(_26953_)
  );
  INV_X1 _35093_ (
    .A(_26953_),
    .ZN(_26954_)
  );
  AND2_X1 _35094_ (
    .A1(_21844_),
    .A2(_22149_),
    .ZN(_26955_)
  );
  INV_X1 _35095_ (
    .A(_26955_),
    .ZN(_26956_)
  );
  AND2_X1 _35096_ (
    .A1(_00008_[0]),
    .A2(_26956_),
    .ZN(_26957_)
  );
  AND2_X1 _35097_ (
    .A1(_26954_),
    .A2(_26957_),
    .ZN(_26958_)
  );
  INV_X1 _35098_ (
    .A(_26958_),
    .ZN(_26959_)
  );
  AND2_X1 _35099_ (
    .A1(_26952_),
    .A2(_26959_),
    .ZN(_26960_)
  );
  AND2_X1 _35100_ (
    .A1(_22148_),
    .A2(_26960_),
    .ZN(_26961_)
  );
  INV_X1 _35101_ (
    .A(_26961_),
    .ZN(_26962_)
  );
  AND2_X1 _35102_ (
    .A1(_21948_),
    .A2(_00008_[2]),
    .ZN(_26963_)
  );
  INV_X1 _35103_ (
    .A(_26963_),
    .ZN(_26964_)
  );
  AND2_X1 _35104_ (
    .A1(_21932_),
    .A2(_22149_),
    .ZN(_26965_)
  );
  INV_X1 _35105_ (
    .A(_26965_),
    .ZN(_26966_)
  );
  AND2_X1 _35106_ (
    .A1(_00008_[0]),
    .A2(_26966_),
    .ZN(_26967_)
  );
  AND2_X1 _35107_ (
    .A1(_26964_),
    .A2(_26967_),
    .ZN(_26968_)
  );
  INV_X1 _35108_ (
    .A(_26968_),
    .ZN(_26969_)
  );
  AND2_X1 _35109_ (
    .A1(_21882_),
    .A2(_22149_),
    .ZN(_26970_)
  );
  INV_X1 _35110_ (
    .A(_26970_),
    .ZN(_26971_)
  );
  AND2_X1 _35111_ (
    .A1(_21860_),
    .A2(_00008_[2]),
    .ZN(_26972_)
  );
  INV_X1 _35112_ (
    .A(_26972_),
    .ZN(_26973_)
  );
  AND2_X1 _35113_ (
    .A1(_26971_),
    .A2(_26973_),
    .ZN(_26974_)
  );
  AND2_X1 _35114_ (
    .A1(_22147_),
    .A2(_26974_),
    .ZN(_26975_)
  );
  INV_X1 _35115_ (
    .A(_26975_),
    .ZN(_26976_)
  );
  AND2_X1 _35116_ (
    .A1(_26969_),
    .A2(_26976_),
    .ZN(_26977_)
  );
  AND2_X1 _35117_ (
    .A1(_00008_[1]),
    .A2(_26977_),
    .ZN(_26978_)
  );
  INV_X1 _35118_ (
    .A(_26978_),
    .ZN(_26979_)
  );
  AND2_X1 _35119_ (
    .A1(_00008_[4]),
    .A2(_26979_),
    .ZN(_26980_)
  );
  AND2_X1 _35120_ (
    .A1(_26962_),
    .A2(_26980_),
    .ZN(_26981_)
  );
  INV_X1 _35121_ (
    .A(_26981_),
    .ZN(_26982_)
  );
  AND2_X1 _35122_ (
    .A1(_26945_),
    .A2(_26982_),
    .ZN(_26983_)
  );
  AND2_X1 _35123_ (
    .A1(_00008_[3]),
    .A2(_26983_),
    .ZN(_26984_)
  );
  INV_X1 _35124_ (
    .A(_26984_),
    .ZN(_26985_)
  );
  AND2_X1 _35125_ (
    .A1(\cpuregs[16] [23]),
    .A2(_22147_),
    .ZN(_26986_)
  );
  INV_X1 _35126_ (
    .A(_26986_),
    .ZN(_26987_)
  );
  AND2_X1 _35127_ (
    .A1(\cpuregs[17] [23]),
    .A2(_00008_[0]),
    .ZN(_26988_)
  );
  INV_X1 _35128_ (
    .A(_26988_),
    .ZN(_26989_)
  );
  AND2_X1 _35129_ (
    .A1(_26987_),
    .A2(_26989_),
    .ZN(_26990_)
  );
  INV_X1 _35130_ (
    .A(_26990_),
    .ZN(_26991_)
  );
  AND2_X1 _35131_ (
    .A1(_22149_),
    .A2(_26991_),
    .ZN(_26992_)
  );
  INV_X1 _35132_ (
    .A(_26992_),
    .ZN(_26993_)
  );
  AND2_X1 _35133_ (
    .A1(\cpuregs[20] [23]),
    .A2(_22147_),
    .ZN(_26994_)
  );
  INV_X1 _35134_ (
    .A(_26994_),
    .ZN(_26995_)
  );
  AND2_X1 _35135_ (
    .A1(\cpuregs[21] [23]),
    .A2(_00008_[0]),
    .ZN(_26996_)
  );
  INV_X1 _35136_ (
    .A(_26996_),
    .ZN(_26997_)
  );
  AND2_X1 _35137_ (
    .A1(_26995_),
    .A2(_26997_),
    .ZN(_26998_)
  );
  INV_X1 _35138_ (
    .A(_26998_),
    .ZN(_26999_)
  );
  AND2_X1 _35139_ (
    .A1(_00008_[2]),
    .A2(_26999_),
    .ZN(_27000_)
  );
  INV_X1 _35140_ (
    .A(_27000_),
    .ZN(_27001_)
  );
  AND2_X1 _35141_ (
    .A1(_22148_),
    .A2(_27001_),
    .ZN(_27002_)
  );
  AND2_X1 _35142_ (
    .A1(_26993_),
    .A2(_27002_),
    .ZN(_27003_)
  );
  INV_X1 _35143_ (
    .A(_27003_),
    .ZN(_27004_)
  );
  AND2_X1 _35144_ (
    .A1(_21608_),
    .A2(_22149_),
    .ZN(_27005_)
  );
  INV_X1 _35145_ (
    .A(_27005_),
    .ZN(_27006_)
  );
  AND2_X1 _35146_ (
    .A1(_21428_),
    .A2(_00008_[2]),
    .ZN(_27007_)
  );
  INV_X1 _35147_ (
    .A(_27007_),
    .ZN(_27008_)
  );
  AND2_X1 _35148_ (
    .A1(_27006_),
    .A2(_27008_),
    .ZN(_27009_)
  );
  AND2_X1 _35149_ (
    .A1(_22147_),
    .A2(_27009_),
    .ZN(_27010_)
  );
  INV_X1 _35150_ (
    .A(_27010_),
    .ZN(_27011_)
  );
  AND2_X1 _35151_ (
    .A1(_21387_),
    .A2(_00008_[2]),
    .ZN(_27012_)
  );
  INV_X1 _35152_ (
    .A(_27012_),
    .ZN(_27013_)
  );
  AND2_X1 _35153_ (
    .A1(_21633_),
    .A2(_22149_),
    .ZN(_27014_)
  );
  INV_X1 _35154_ (
    .A(_27014_),
    .ZN(_27015_)
  );
  AND2_X1 _35155_ (
    .A1(_00008_[0]),
    .A2(_27015_),
    .ZN(_27016_)
  );
  AND2_X1 _35156_ (
    .A1(_27013_),
    .A2(_27016_),
    .ZN(_27017_)
  );
  INV_X1 _35157_ (
    .A(_27017_),
    .ZN(_27018_)
  );
  AND2_X1 _35158_ (
    .A1(_27011_),
    .A2(_27018_),
    .ZN(_27019_)
  );
  AND2_X1 _35159_ (
    .A1(_00008_[1]),
    .A2(_27019_),
    .ZN(_27020_)
  );
  INV_X1 _35160_ (
    .A(_27020_),
    .ZN(_27021_)
  );
  AND2_X1 _35161_ (
    .A1(_21797_),
    .A2(_00008_[2]),
    .ZN(_27022_)
  );
  INV_X1 _35162_ (
    .A(_27022_),
    .ZN(_27023_)
  );
  AND2_X1 _35163_ (
    .A1(_21505_),
    .A2(_22149_),
    .ZN(_27024_)
  );
  INV_X1 _35164_ (
    .A(_27024_),
    .ZN(_27025_)
  );
  AND2_X1 _35165_ (
    .A1(_00008_[0]),
    .A2(_27025_),
    .ZN(_27026_)
  );
  AND2_X1 _35166_ (
    .A1(_27023_),
    .A2(_27026_),
    .ZN(_27027_)
  );
  INV_X1 _35167_ (
    .A(_27027_),
    .ZN(_27028_)
  );
  AND2_X1 _35168_ (
    .A1(_21559_),
    .A2(_22149_),
    .ZN(_27029_)
  );
  INV_X1 _35169_ (
    .A(_27029_),
    .ZN(_27030_)
  );
  AND2_X1 _35170_ (
    .A1(_21825_),
    .A2(_00008_[2]),
    .ZN(_27031_)
  );
  INV_X1 _35171_ (
    .A(_27031_),
    .ZN(_27032_)
  );
  AND2_X1 _35172_ (
    .A1(_27030_),
    .A2(_27032_),
    .ZN(_27033_)
  );
  AND2_X1 _35173_ (
    .A1(_22147_),
    .A2(_27033_),
    .ZN(_27034_)
  );
  INV_X1 _35174_ (
    .A(_27034_),
    .ZN(_27035_)
  );
  AND2_X1 _35175_ (
    .A1(_27028_),
    .A2(_27035_),
    .ZN(_27036_)
  );
  AND2_X1 _35176_ (
    .A1(_00008_[1]),
    .A2(_27036_),
    .ZN(_27037_)
  );
  INV_X1 _35177_ (
    .A(_27037_),
    .ZN(_27038_)
  );
  AND2_X1 _35178_ (
    .A1(_21750_),
    .A2(_00008_[2]),
    .ZN(_27039_)
  );
  INV_X1 _35179_ (
    .A(_27039_),
    .ZN(_27040_)
  );
  AND2_X1 _35180_ (
    .A1(_21530_),
    .A2(_22149_),
    .ZN(_27041_)
  );
  INV_X1 _35181_ (
    .A(_27041_),
    .ZN(_27042_)
  );
  AND2_X1 _35182_ (
    .A1(_00008_[0]),
    .A2(_27042_),
    .ZN(_27043_)
  );
  AND2_X1 _35183_ (
    .A1(_27040_),
    .A2(_27043_),
    .ZN(_27044_)
  );
  INV_X1 _35184_ (
    .A(_27044_),
    .ZN(_27045_)
  );
  AND2_X1 _35185_ (
    .A1(_21971_),
    .A2(_22149_),
    .ZN(_27046_)
  );
  INV_X1 _35186_ (
    .A(_27046_),
    .ZN(_27047_)
  );
  AND2_X1 _35187_ (
    .A1(_21687_),
    .A2(_00008_[2]),
    .ZN(_27048_)
  );
  INV_X1 _35188_ (
    .A(_27048_),
    .ZN(_27049_)
  );
  AND2_X1 _35189_ (
    .A1(_27047_),
    .A2(_27049_),
    .ZN(_27050_)
  );
  AND2_X1 _35190_ (
    .A1(_22147_),
    .A2(_27050_),
    .ZN(_27051_)
  );
  INV_X1 _35191_ (
    .A(_27051_),
    .ZN(_27052_)
  );
  AND2_X1 _35192_ (
    .A1(_27045_),
    .A2(_27052_),
    .ZN(_27053_)
  );
  AND2_X1 _35193_ (
    .A1(_22148_),
    .A2(_27053_),
    .ZN(_27054_)
  );
  INV_X1 _35194_ (
    .A(_27054_),
    .ZN(_27055_)
  );
  AND2_X1 _35195_ (
    .A1(_27038_),
    .A2(_27055_),
    .ZN(_27056_)
  );
  AND2_X1 _35196_ (
    .A1(_00008_[4]),
    .A2(_27021_),
    .ZN(_27057_)
  );
  AND2_X1 _35197_ (
    .A1(_27004_),
    .A2(_27057_),
    .ZN(_27058_)
  );
  INV_X1 _35198_ (
    .A(_27058_),
    .ZN(_27059_)
  );
  AND2_X1 _35199_ (
    .A1(_22151_),
    .A2(_27056_),
    .ZN(_27060_)
  );
  INV_X1 _35200_ (
    .A(_27060_),
    .ZN(_27061_)
  );
  AND2_X1 _35201_ (
    .A1(_27059_),
    .A2(_27061_),
    .ZN(_27062_)
  );
  AND2_X1 _35202_ (
    .A1(_22150_),
    .A2(_27062_),
    .ZN(_27063_)
  );
  INV_X1 _35203_ (
    .A(_27063_),
    .ZN(_27064_)
  );
  AND2_X1 _35204_ (
    .A1(_22546_),
    .A2(_27064_),
    .ZN(_27065_)
  );
  AND2_X1 _35205_ (
    .A1(_26985_),
    .A2(_27065_),
    .ZN(_27066_)
  );
  INV_X1 _35206_ (
    .A(_27066_),
    .ZN(_27067_)
  );
  AND2_X1 _35207_ (
    .A1(_26908_),
    .A2(_27067_),
    .ZN(_27068_)
  );
  INV_X1 _35208_ (
    .A(_27068_),
    .ZN(_27069_)
  );
  AND2_X1 _35209_ (
    .A1(_22271_),
    .A2(_27069_),
    .ZN(_27070_)
  );
  INV_X1 _35210_ (
    .A(_27070_),
    .ZN(_27071_)
  );
  AND2_X1 _35211_ (
    .A1(reg_op1[22]),
    .A2(_22285_),
    .ZN(_27072_)
  );
  INV_X1 _35212_ (
    .A(_27072_),
    .ZN(_27073_)
  );
  AND2_X1 _35213_ (
    .A1(_26444_),
    .A2(_27073_),
    .ZN(_27074_)
  );
  INV_X1 _35214_ (
    .A(_27074_),
    .ZN(_27075_)
  );
  AND2_X1 _35215_ (
    .A1(_22572_),
    .A2(_27075_),
    .ZN(_27076_)
  );
  INV_X1 _35216_ (
    .A(_27076_),
    .ZN(_27077_)
  );
  AND2_X1 _35217_ (
    .A1(reg_op1[27]),
    .A2(_22290_),
    .ZN(_27078_)
  );
  INV_X1 _35218_ (
    .A(_27078_),
    .ZN(_27079_)
  );
  AND2_X1 _35219_ (
    .A1(_26441_),
    .A2(_27079_),
    .ZN(_27080_)
  );
  INV_X1 _35220_ (
    .A(_27080_),
    .ZN(_27081_)
  );
  AND2_X1 _35221_ (
    .A1(_22573_),
    .A2(_27081_),
    .ZN(_27082_)
  );
  INV_X1 _35222_ (
    .A(_27082_),
    .ZN(_27083_)
  );
  AND2_X1 _35223_ (
    .A1(_27077_),
    .A2(_27083_),
    .ZN(_27084_)
  );
  INV_X1 _35224_ (
    .A(_27084_),
    .ZN(_27085_)
  );
  AND2_X1 _35225_ (
    .A1(_22295_),
    .A2(_27085_),
    .ZN(_27086_)
  );
  INV_X1 _35226_ (
    .A(_27086_),
    .ZN(_27087_)
  );
  AND2_X1 _35227_ (
    .A1(_22333_),
    .A2(_27087_),
    .ZN(_27088_)
  );
  AND2_X1 _35228_ (
    .A1(_27071_),
    .A2(_27088_),
    .ZN(_27089_)
  );
  AND2_X1 _35229_ (
    .A1(_26906_),
    .A2(_27089_),
    .ZN(_27090_)
  );
  INV_X1 _35230_ (
    .A(_27090_),
    .ZN(_27091_)
  );
  AND2_X1 _35231_ (
    .A1(_26891_),
    .A2(_27091_),
    .ZN(_00080_)
  );
  AND2_X1 _35232_ (
    .A1(_21191_),
    .A2(_22334_),
    .ZN(_27092_)
  );
  INV_X1 _35233_ (
    .A(_27092_),
    .ZN(_27093_)
  );
  AND2_X1 _35234_ (
    .A1(reg_pc[24]),
    .A2(_22335_),
    .ZN(_27094_)
  );
  INV_X1 _35235_ (
    .A(_27094_),
    .ZN(_27095_)
  );
  AND2_X1 _35236_ (
    .A1(_21453_),
    .A2(_22149_),
    .ZN(_27096_)
  );
  INV_X1 _35237_ (
    .A(_27096_),
    .ZN(_27097_)
  );
  AND2_X1 _35238_ (
    .A1(_21664_),
    .A2(_00008_[2]),
    .ZN(_27098_)
  );
  INV_X1 _35239_ (
    .A(_27098_),
    .ZN(_27099_)
  );
  AND2_X1 _35240_ (
    .A1(_27097_),
    .A2(_27099_),
    .ZN(_27100_)
  );
  AND2_X1 _35241_ (
    .A1(_22147_),
    .A2(_27100_),
    .ZN(_27101_)
  );
  INV_X1 _35242_ (
    .A(_27101_),
    .ZN(_27102_)
  );
  AND2_X1 _35243_ (
    .A1(_21774_),
    .A2(_00008_[2]),
    .ZN(_27103_)
  );
  INV_X1 _35244_ (
    .A(_27103_),
    .ZN(_27104_)
  );
  AND2_X1 _35245_ (
    .A1(_21475_),
    .A2(_22149_),
    .ZN(_27105_)
  );
  INV_X1 _35246_ (
    .A(_27105_),
    .ZN(_27106_)
  );
  AND2_X1 _35247_ (
    .A1(_00008_[0]),
    .A2(_27104_),
    .ZN(_27107_)
  );
  AND2_X1 _35248_ (
    .A1(_27106_),
    .A2(_27107_),
    .ZN(_27108_)
  );
  INV_X1 _35249_ (
    .A(_27108_),
    .ZN(_27109_)
  );
  AND2_X1 _35250_ (
    .A1(_27102_),
    .A2(_27109_),
    .ZN(_27110_)
  );
  AND2_X1 _35251_ (
    .A1(_22148_),
    .A2(_27110_),
    .ZN(_27111_)
  );
  INV_X1 _35252_ (
    .A(_27111_),
    .ZN(_27112_)
  );
  AND2_X1 _35253_ (
    .A1(_21609_),
    .A2(_22149_),
    .ZN(_27113_)
  );
  INV_X1 _35254_ (
    .A(_27113_),
    .ZN(_27114_)
  );
  AND2_X1 _35255_ (
    .A1(_21429_),
    .A2(_00008_[2]),
    .ZN(_27115_)
  );
  INV_X1 _35256_ (
    .A(_27115_),
    .ZN(_27116_)
  );
  AND2_X1 _35257_ (
    .A1(_27114_),
    .A2(_27116_),
    .ZN(_27117_)
  );
  AND2_X1 _35258_ (
    .A1(_22147_),
    .A2(_27117_),
    .ZN(_27118_)
  );
  INV_X1 _35259_ (
    .A(_27118_),
    .ZN(_27119_)
  );
  AND2_X1 _35260_ (
    .A1(_21388_),
    .A2(_00008_[2]),
    .ZN(_27120_)
  );
  INV_X1 _35261_ (
    .A(_27120_),
    .ZN(_27121_)
  );
  AND2_X1 _35262_ (
    .A1(_21634_),
    .A2(_22149_),
    .ZN(_27122_)
  );
  INV_X1 _35263_ (
    .A(_27122_),
    .ZN(_27123_)
  );
  AND2_X1 _35264_ (
    .A1(_00008_[0]),
    .A2(_27123_),
    .ZN(_27124_)
  );
  AND2_X1 _35265_ (
    .A1(_27121_),
    .A2(_27124_),
    .ZN(_27125_)
  );
  INV_X1 _35266_ (
    .A(_27125_),
    .ZN(_27126_)
  );
  AND2_X1 _35267_ (
    .A1(_27119_),
    .A2(_27126_),
    .ZN(_27127_)
  );
  AND2_X1 _35268_ (
    .A1(_00008_[1]),
    .A2(_27127_),
    .ZN(_27128_)
  );
  INV_X1 _35269_ (
    .A(_27128_),
    .ZN(_27129_)
  );
  AND2_X1 _35270_ (
    .A1(_27112_),
    .A2(_27129_),
    .ZN(_27130_)
  );
  AND2_X1 _35271_ (
    .A1(\cpuregs[27] [24]),
    .A2(_00008_[0]),
    .ZN(_27131_)
  );
  INV_X1 _35272_ (
    .A(_27131_),
    .ZN(_27132_)
  );
  AND2_X1 _35273_ (
    .A1(\cpuregs[26] [24]),
    .A2(_22147_),
    .ZN(_27133_)
  );
  INV_X1 _35274_ (
    .A(_27133_),
    .ZN(_27134_)
  );
  AND2_X1 _35275_ (
    .A1(_22149_),
    .A2(_27134_),
    .ZN(_27135_)
  );
  AND2_X1 _35276_ (
    .A1(_27132_),
    .A2(_27135_),
    .ZN(_27136_)
  );
  INV_X1 _35277_ (
    .A(_27136_),
    .ZN(_27137_)
  );
  AND2_X1 _35278_ (
    .A1(\cpuregs[31] [24]),
    .A2(_00008_[0]),
    .ZN(_27138_)
  );
  INV_X1 _35279_ (
    .A(_27138_),
    .ZN(_27139_)
  );
  AND2_X1 _35280_ (
    .A1(\cpuregs[30] [24]),
    .A2(_22147_),
    .ZN(_27140_)
  );
  INV_X1 _35281_ (
    .A(_27140_),
    .ZN(_27141_)
  );
  AND2_X1 _35282_ (
    .A1(_00008_[2]),
    .A2(_27141_),
    .ZN(_27142_)
  );
  AND2_X1 _35283_ (
    .A1(_27139_),
    .A2(_27142_),
    .ZN(_27143_)
  );
  INV_X1 _35284_ (
    .A(_27143_),
    .ZN(_27144_)
  );
  AND2_X1 _35285_ (
    .A1(_27137_),
    .A2(_27144_),
    .ZN(_27145_)
  );
  INV_X1 _35286_ (
    .A(_27145_),
    .ZN(_27146_)
  );
  AND2_X1 _35287_ (
    .A1(_00008_[1]),
    .A2(_27146_),
    .ZN(_27147_)
  );
  INV_X1 _35288_ (
    .A(_27147_),
    .ZN(_27148_)
  );
  AND2_X1 _35289_ (
    .A1(\cpuregs[25] [24]),
    .A2(_00008_[0]),
    .ZN(_27149_)
  );
  INV_X1 _35290_ (
    .A(_27149_),
    .ZN(_27150_)
  );
  AND2_X1 _35291_ (
    .A1(\cpuregs[24] [24]),
    .A2(_22147_),
    .ZN(_27151_)
  );
  INV_X1 _35292_ (
    .A(_27151_),
    .ZN(_27152_)
  );
  AND2_X1 _35293_ (
    .A1(_22149_),
    .A2(_27152_),
    .ZN(_27153_)
  );
  AND2_X1 _35294_ (
    .A1(_27150_),
    .A2(_27153_),
    .ZN(_27154_)
  );
  INV_X1 _35295_ (
    .A(_27154_),
    .ZN(_27155_)
  );
  AND2_X1 _35296_ (
    .A1(\cpuregs[29] [24]),
    .A2(_00008_[0]),
    .ZN(_27156_)
  );
  INV_X1 _35297_ (
    .A(_27156_),
    .ZN(_27157_)
  );
  AND2_X1 _35298_ (
    .A1(\cpuregs[28] [24]),
    .A2(_22147_),
    .ZN(_27158_)
  );
  INV_X1 _35299_ (
    .A(_27158_),
    .ZN(_27159_)
  );
  AND2_X1 _35300_ (
    .A1(_00008_[2]),
    .A2(_27159_),
    .ZN(_27160_)
  );
  AND2_X1 _35301_ (
    .A1(_27157_),
    .A2(_27160_),
    .ZN(_27161_)
  );
  INV_X1 _35302_ (
    .A(_27161_),
    .ZN(_27162_)
  );
  AND2_X1 _35303_ (
    .A1(_27155_),
    .A2(_27162_),
    .ZN(_27163_)
  );
  INV_X1 _35304_ (
    .A(_27163_),
    .ZN(_27164_)
  );
  AND2_X1 _35305_ (
    .A1(_22148_),
    .A2(_27164_),
    .ZN(_27165_)
  );
  INV_X1 _35306_ (
    .A(_27165_),
    .ZN(_27166_)
  );
  AND2_X1 _35307_ (
    .A1(_00008_[3]),
    .A2(_27148_),
    .ZN(_27167_)
  );
  AND2_X1 _35308_ (
    .A1(_27166_),
    .A2(_27167_),
    .ZN(_27168_)
  );
  INV_X1 _35309_ (
    .A(_27168_),
    .ZN(_27169_)
  );
  AND2_X1 _35310_ (
    .A1(_22150_),
    .A2(_27130_),
    .ZN(_27170_)
  );
  INV_X1 _35311_ (
    .A(_27170_),
    .ZN(_27171_)
  );
  AND2_X1 _35312_ (
    .A1(_00008_[4]),
    .A2(_27171_),
    .ZN(_27172_)
  );
  AND2_X1 _35313_ (
    .A1(_27169_),
    .A2(_27172_),
    .ZN(_27173_)
  );
  INV_X1 _35314_ (
    .A(_27173_),
    .ZN(_27174_)
  );
  AND2_X1 _35315_ (
    .A1(\cpuregs[10] [24]),
    .A2(_22149_),
    .ZN(_27175_)
  );
  INV_X1 _35316_ (
    .A(_27175_),
    .ZN(_27176_)
  );
  AND2_X1 _35317_ (
    .A1(\cpuregs[14] [24]),
    .A2(_00008_[2]),
    .ZN(_27177_)
  );
  INV_X1 _35318_ (
    .A(_27177_),
    .ZN(_27178_)
  );
  AND2_X1 _35319_ (
    .A1(_22147_),
    .A2(_27178_),
    .ZN(_27179_)
  );
  AND2_X1 _35320_ (
    .A1(_27176_),
    .A2(_27179_),
    .ZN(_27180_)
  );
  INV_X1 _35321_ (
    .A(_27180_),
    .ZN(_27181_)
  );
  AND2_X1 _35322_ (
    .A1(\cpuregs[15] [24]),
    .A2(_00008_[2]),
    .ZN(_27182_)
  );
  INV_X1 _35323_ (
    .A(_27182_),
    .ZN(_27183_)
  );
  AND2_X1 _35324_ (
    .A1(\cpuregs[11] [24]),
    .A2(_22149_),
    .ZN(_27184_)
  );
  INV_X1 _35325_ (
    .A(_27184_),
    .ZN(_27185_)
  );
  AND2_X1 _35326_ (
    .A1(_00008_[0]),
    .A2(_27185_),
    .ZN(_27186_)
  );
  AND2_X1 _35327_ (
    .A1(_27183_),
    .A2(_27186_),
    .ZN(_27187_)
  );
  INV_X1 _35328_ (
    .A(_27187_),
    .ZN(_27188_)
  );
  AND2_X1 _35329_ (
    .A1(_27181_),
    .A2(_27188_),
    .ZN(_27189_)
  );
  AND2_X1 _35330_ (
    .A1(\cpuregs[2] [24]),
    .A2(_22149_),
    .ZN(_27190_)
  );
  INV_X1 _35331_ (
    .A(_27190_),
    .ZN(_27191_)
  );
  AND2_X1 _35332_ (
    .A1(\cpuregs[6] [24]),
    .A2(_00008_[2]),
    .ZN(_27192_)
  );
  INV_X1 _35333_ (
    .A(_27192_),
    .ZN(_27193_)
  );
  AND2_X1 _35334_ (
    .A1(_22147_),
    .A2(_27193_),
    .ZN(_27194_)
  );
  AND2_X1 _35335_ (
    .A1(_27191_),
    .A2(_27194_),
    .ZN(_27195_)
  );
  INV_X1 _35336_ (
    .A(_27195_),
    .ZN(_27196_)
  );
  AND2_X1 _35337_ (
    .A1(\cpuregs[3] [24]),
    .A2(_22149_),
    .ZN(_27197_)
  );
  INV_X1 _35338_ (
    .A(_27197_),
    .ZN(_27198_)
  );
  AND2_X1 _35339_ (
    .A1(\cpuregs[7] [24]),
    .A2(_00008_[2]),
    .ZN(_27199_)
  );
  INV_X1 _35340_ (
    .A(_27199_),
    .ZN(_27200_)
  );
  AND2_X1 _35341_ (
    .A1(_00008_[0]),
    .A2(_27200_),
    .ZN(_27201_)
  );
  AND2_X1 _35342_ (
    .A1(_27198_),
    .A2(_27201_),
    .ZN(_27202_)
  );
  INV_X1 _35343_ (
    .A(_27202_),
    .ZN(_27203_)
  );
  AND2_X1 _35344_ (
    .A1(_00008_[3]),
    .A2(_27189_),
    .ZN(_27204_)
  );
  INV_X1 _35345_ (
    .A(_27204_),
    .ZN(_27205_)
  );
  AND2_X1 _35346_ (
    .A1(_22150_),
    .A2(_27203_),
    .ZN(_27206_)
  );
  AND2_X1 _35347_ (
    .A1(_27196_),
    .A2(_27206_),
    .ZN(_27207_)
  );
  INV_X1 _35348_ (
    .A(_27207_),
    .ZN(_27208_)
  );
  AND2_X1 _35349_ (
    .A1(_27205_),
    .A2(_27208_),
    .ZN(_27209_)
  );
  INV_X1 _35350_ (
    .A(_27209_),
    .ZN(_27210_)
  );
  AND2_X1 _35351_ (
    .A1(\cpuregs[8] [24]),
    .A2(_22149_),
    .ZN(_27211_)
  );
  INV_X1 _35352_ (
    .A(_27211_),
    .ZN(_27212_)
  );
  AND2_X1 _35353_ (
    .A1(\cpuregs[12] [24]),
    .A2(_00008_[2]),
    .ZN(_27213_)
  );
  INV_X1 _35354_ (
    .A(_27213_),
    .ZN(_27214_)
  );
  AND2_X1 _35355_ (
    .A1(_22147_),
    .A2(_27214_),
    .ZN(_27215_)
  );
  AND2_X1 _35356_ (
    .A1(_27212_),
    .A2(_27215_),
    .ZN(_27216_)
  );
  INV_X1 _35357_ (
    .A(_27216_),
    .ZN(_27217_)
  );
  AND2_X1 _35358_ (
    .A1(\cpuregs[13] [24]),
    .A2(_00008_[2]),
    .ZN(_27218_)
  );
  INV_X1 _35359_ (
    .A(_27218_),
    .ZN(_27219_)
  );
  AND2_X1 _35360_ (
    .A1(\cpuregs[9] [24]),
    .A2(_22149_),
    .ZN(_27220_)
  );
  INV_X1 _35361_ (
    .A(_27220_),
    .ZN(_27221_)
  );
  AND2_X1 _35362_ (
    .A1(_00008_[0]),
    .A2(_27221_),
    .ZN(_27222_)
  );
  AND2_X1 _35363_ (
    .A1(_27219_),
    .A2(_27222_),
    .ZN(_27223_)
  );
  INV_X1 _35364_ (
    .A(_27223_),
    .ZN(_27224_)
  );
  AND2_X1 _35365_ (
    .A1(_27217_),
    .A2(_27224_),
    .ZN(_27225_)
  );
  AND2_X1 _35366_ (
    .A1(\cpuregs[0] [24]),
    .A2(_22149_),
    .ZN(_27226_)
  );
  INV_X1 _35367_ (
    .A(_27226_),
    .ZN(_27227_)
  );
  AND2_X1 _35368_ (
    .A1(\cpuregs[4] [24]),
    .A2(_00008_[2]),
    .ZN(_27228_)
  );
  INV_X1 _35369_ (
    .A(_27228_),
    .ZN(_27229_)
  );
  AND2_X1 _35370_ (
    .A1(_22147_),
    .A2(_27229_),
    .ZN(_27230_)
  );
  AND2_X1 _35371_ (
    .A1(_27227_),
    .A2(_27230_),
    .ZN(_27231_)
  );
  INV_X1 _35372_ (
    .A(_27231_),
    .ZN(_27232_)
  );
  AND2_X1 _35373_ (
    .A1(\cpuregs[1] [24]),
    .A2(_22149_),
    .ZN(_27233_)
  );
  INV_X1 _35374_ (
    .A(_27233_),
    .ZN(_27234_)
  );
  AND2_X1 _35375_ (
    .A1(\cpuregs[5] [24]),
    .A2(_00008_[2]),
    .ZN(_27235_)
  );
  INV_X1 _35376_ (
    .A(_27235_),
    .ZN(_27236_)
  );
  AND2_X1 _35377_ (
    .A1(_00008_[0]),
    .A2(_27236_),
    .ZN(_27237_)
  );
  AND2_X1 _35378_ (
    .A1(_27234_),
    .A2(_27237_),
    .ZN(_27238_)
  );
  INV_X1 _35379_ (
    .A(_27238_),
    .ZN(_27239_)
  );
  AND2_X1 _35380_ (
    .A1(_00008_[3]),
    .A2(_27225_),
    .ZN(_27240_)
  );
  INV_X1 _35381_ (
    .A(_27240_),
    .ZN(_27241_)
  );
  AND2_X1 _35382_ (
    .A1(_22150_),
    .A2(_27239_),
    .ZN(_27242_)
  );
  AND2_X1 _35383_ (
    .A1(_27232_),
    .A2(_27242_),
    .ZN(_27243_)
  );
  INV_X1 _35384_ (
    .A(_27243_),
    .ZN(_27244_)
  );
  AND2_X1 _35385_ (
    .A1(_27241_),
    .A2(_27244_),
    .ZN(_27245_)
  );
  INV_X1 _35386_ (
    .A(_27245_),
    .ZN(_27246_)
  );
  AND2_X1 _35387_ (
    .A1(_22148_),
    .A2(_27246_),
    .ZN(_27247_)
  );
  INV_X1 _35388_ (
    .A(_27247_),
    .ZN(_27248_)
  );
  AND2_X1 _35389_ (
    .A1(_00008_[1]),
    .A2(_27210_),
    .ZN(_27249_)
  );
  INV_X1 _35390_ (
    .A(_27249_),
    .ZN(_27250_)
  );
  AND2_X1 _35391_ (
    .A1(_27248_),
    .A2(_27250_),
    .ZN(_27251_)
  );
  AND2_X1 _35392_ (
    .A1(_22151_),
    .A2(_27251_),
    .ZN(_27252_)
  );
  INV_X1 _35393_ (
    .A(_27252_),
    .ZN(_27253_)
  );
  AND2_X1 _35394_ (
    .A1(_22546_),
    .A2(_27174_),
    .ZN(_27254_)
  );
  AND2_X1 _35395_ (
    .A1(_27253_),
    .A2(_27254_),
    .ZN(_27255_)
  );
  INV_X1 _35396_ (
    .A(_27255_),
    .ZN(_27256_)
  );
  AND2_X1 _35397_ (
    .A1(_27095_),
    .A2(_27256_),
    .ZN(_27257_)
  );
  INV_X1 _35398_ (
    .A(_27257_),
    .ZN(_27258_)
  );
  AND2_X1 _35399_ (
    .A1(_22271_),
    .A2(_27258_),
    .ZN(_27259_)
  );
  INV_X1 _35400_ (
    .A(_27259_),
    .ZN(_27260_)
  );
  AND2_X1 _35401_ (
    .A1(reg_op1[23]),
    .A2(_22285_),
    .ZN(_27261_)
  );
  INV_X1 _35402_ (
    .A(_27261_),
    .ZN(_27262_)
  );
  AND2_X1 _35403_ (
    .A1(_26661_),
    .A2(_27262_),
    .ZN(_27263_)
  );
  AND2_X1 _35404_ (
    .A1(reg_op1[28]),
    .A2(_22290_),
    .ZN(_27264_)
  );
  INV_X1 _35405_ (
    .A(_27264_),
    .ZN(_27265_)
  );
  AND2_X1 _35406_ (
    .A1(_26658_),
    .A2(_27265_),
    .ZN(_27266_)
  );
  AND2_X1 _35407_ (
    .A1(_22572_),
    .A2(_27263_),
    .ZN(_27267_)
  );
  INV_X1 _35408_ (
    .A(_27267_),
    .ZN(_27268_)
  );
  AND2_X1 _35409_ (
    .A1(_22573_),
    .A2(_27266_),
    .ZN(_27269_)
  );
  INV_X1 _35410_ (
    .A(_27269_),
    .ZN(_27270_)
  );
  AND2_X1 _35411_ (
    .A1(_22295_),
    .A2(_27270_),
    .ZN(_27271_)
  );
  AND2_X1 _35412_ (
    .A1(_27268_),
    .A2(_27271_),
    .ZN(_27272_)
  );
  INV_X1 _35413_ (
    .A(_27272_),
    .ZN(_27273_)
  );
  AND2_X1 _35414_ (
    .A1(_22333_),
    .A2(_27273_),
    .ZN(_27274_)
  );
  AND2_X1 _35415_ (
    .A1(_27260_),
    .A2(_27274_),
    .ZN(_27275_)
  );
  AND2_X1 _35416_ (
    .A1(reg_op1[24]),
    .A2(decoded_imm[24]),
    .ZN(_27276_)
  );
  INV_X1 _35417_ (
    .A(_27276_),
    .ZN(_27277_)
  );
  AND2_X1 _35418_ (
    .A1(_21191_),
    .A2(_21985_),
    .ZN(_27278_)
  );
  INV_X1 _35419_ (
    .A(_27278_),
    .ZN(_27279_)
  );
  AND2_X1 _35420_ (
    .A1(_27277_),
    .A2(_27279_),
    .ZN(_27280_)
  );
  INV_X1 _35421_ (
    .A(_27280_),
    .ZN(_27281_)
  );
  AND2_X1 _35422_ (
    .A1(_26893_),
    .A2(_26898_),
    .ZN(_27282_)
  );
  INV_X1 _35423_ (
    .A(_27282_),
    .ZN(_27283_)
  );
  AND2_X1 _35424_ (
    .A1(_26895_),
    .A2(_26899_),
    .ZN(_27284_)
  );
  INV_X1 _35425_ (
    .A(_27284_),
    .ZN(_27285_)
  );
  AND2_X1 _35426_ (
    .A1(_26895_),
    .A2(_27283_),
    .ZN(_27286_)
  );
  AND2_X1 _35427_ (
    .A1(_26893_),
    .A2(_27285_),
    .ZN(_27287_)
  );
  AND2_X1 _35428_ (
    .A1(_27280_),
    .A2(_27286_),
    .ZN(_27288_)
  );
  INV_X1 _35429_ (
    .A(_27288_),
    .ZN(_27289_)
  );
  AND2_X1 _35430_ (
    .A1(_27281_),
    .A2(_27287_),
    .ZN(_27290_)
  );
  INV_X1 _35431_ (
    .A(_27290_),
    .ZN(_27291_)
  );
  AND2_X1 _35432_ (
    .A1(_27289_),
    .A2(_27291_),
    .ZN(_27292_)
  );
  AND2_X1 _35433_ (
    .A1(_22559_),
    .A2(_27292_),
    .ZN(_27293_)
  );
  INV_X1 _35434_ (
    .A(_27293_),
    .ZN(_27294_)
  );
  AND2_X1 _35435_ (
    .A1(_27275_),
    .A2(_27294_),
    .ZN(_27295_)
  );
  INV_X1 _35436_ (
    .A(_27295_),
    .ZN(_27296_)
  );
  AND2_X1 _35437_ (
    .A1(_27093_),
    .A2(_27296_),
    .ZN(_00081_)
  );
  AND2_X1 _35438_ (
    .A1(_21192_),
    .A2(_22334_),
    .ZN(_27297_)
  );
  INV_X1 _35439_ (
    .A(_27297_),
    .ZN(_27298_)
  );
  AND2_X1 _35440_ (
    .A1(reg_pc[25]),
    .A2(_22335_),
    .ZN(_27299_)
  );
  INV_X1 _35441_ (
    .A(_27299_),
    .ZN(_27300_)
  );
  AND2_X1 _35442_ (
    .A1(\cpuregs[13] [25]),
    .A2(_00008_[2]),
    .ZN(_27301_)
  );
  INV_X1 _35443_ (
    .A(_27301_),
    .ZN(_27302_)
  );
  AND2_X1 _35444_ (
    .A1(\cpuregs[9] [25]),
    .A2(_22149_),
    .ZN(_27303_)
  );
  INV_X1 _35445_ (
    .A(_27303_),
    .ZN(_27304_)
  );
  AND2_X1 _35446_ (
    .A1(_27302_),
    .A2(_27304_),
    .ZN(_27305_)
  );
  INV_X1 _35447_ (
    .A(_27305_),
    .ZN(_27306_)
  );
  AND2_X1 _35448_ (
    .A1(_00008_[0]),
    .A2(_27306_),
    .ZN(_27307_)
  );
  INV_X1 _35449_ (
    .A(_27307_),
    .ZN(_27308_)
  );
  AND2_X1 _35450_ (
    .A1(\cpuregs[12] [25]),
    .A2(_00008_[2]),
    .ZN(_27309_)
  );
  INV_X1 _35451_ (
    .A(_27309_),
    .ZN(_27310_)
  );
  AND2_X1 _35452_ (
    .A1(\cpuregs[8] [25]),
    .A2(_22149_),
    .ZN(_27311_)
  );
  INV_X1 _35453_ (
    .A(_27311_),
    .ZN(_27312_)
  );
  AND2_X1 _35454_ (
    .A1(_27310_),
    .A2(_27312_),
    .ZN(_27313_)
  );
  INV_X1 _35455_ (
    .A(_27313_),
    .ZN(_27314_)
  );
  AND2_X1 _35456_ (
    .A1(_22147_),
    .A2(_27314_),
    .ZN(_27315_)
  );
  INV_X1 _35457_ (
    .A(_27315_),
    .ZN(_27316_)
  );
  AND2_X1 _35458_ (
    .A1(_27308_),
    .A2(_27316_),
    .ZN(_27317_)
  );
  AND2_X1 _35459_ (
    .A1(\cpuregs[5] [25]),
    .A2(_00008_[2]),
    .ZN(_27318_)
  );
  INV_X1 _35460_ (
    .A(_27318_),
    .ZN(_27319_)
  );
  AND2_X1 _35461_ (
    .A1(\cpuregs[1] [25]),
    .A2(_22149_),
    .ZN(_27320_)
  );
  INV_X1 _35462_ (
    .A(_27320_),
    .ZN(_27321_)
  );
  AND2_X1 _35463_ (
    .A1(\cpuregs[4] [25]),
    .A2(_00008_[2]),
    .ZN(_27322_)
  );
  INV_X1 _35464_ (
    .A(_27322_),
    .ZN(_27323_)
  );
  AND2_X1 _35465_ (
    .A1(\cpuregs[0] [25]),
    .A2(_22149_),
    .ZN(_27324_)
  );
  INV_X1 _35466_ (
    .A(_27324_),
    .ZN(_27325_)
  );
  AND2_X1 _35467_ (
    .A1(_27323_),
    .A2(_27325_),
    .ZN(_27326_)
  );
  AND2_X1 _35468_ (
    .A1(_22147_),
    .A2(_27326_),
    .ZN(_27327_)
  );
  INV_X1 _35469_ (
    .A(_27327_),
    .ZN(_27328_)
  );
  AND2_X1 _35470_ (
    .A1(_00008_[0]),
    .A2(_27319_),
    .ZN(_27329_)
  );
  AND2_X1 _35471_ (
    .A1(_27321_),
    .A2(_27329_),
    .ZN(_27330_)
  );
  INV_X1 _35472_ (
    .A(_27330_),
    .ZN(_27331_)
  );
  AND2_X1 _35473_ (
    .A1(_27328_),
    .A2(_27331_),
    .ZN(_27332_)
  );
  INV_X1 _35474_ (
    .A(_27332_),
    .ZN(_27333_)
  );
  AND2_X1 _35475_ (
    .A1(_22150_),
    .A2(_27333_),
    .ZN(_27334_)
  );
  INV_X1 _35476_ (
    .A(_27334_),
    .ZN(_27335_)
  );
  AND2_X1 _35477_ (
    .A1(_00008_[3]),
    .A2(_27317_),
    .ZN(_27336_)
  );
  INV_X1 _35478_ (
    .A(_27336_),
    .ZN(_27337_)
  );
  AND2_X1 _35479_ (
    .A1(_22148_),
    .A2(_27337_),
    .ZN(_27338_)
  );
  AND2_X1 _35480_ (
    .A1(_27335_),
    .A2(_27338_),
    .ZN(_27339_)
  );
  INV_X1 _35481_ (
    .A(_27339_),
    .ZN(_27340_)
  );
  AND2_X1 _35482_ (
    .A1(\cpuregs[7] [25]),
    .A2(_00008_[0]),
    .ZN(_27341_)
  );
  INV_X1 _35483_ (
    .A(_27341_),
    .ZN(_27342_)
  );
  AND2_X1 _35484_ (
    .A1(\cpuregs[6] [25]),
    .A2(_22147_),
    .ZN(_27343_)
  );
  INV_X1 _35485_ (
    .A(_27343_),
    .ZN(_27344_)
  );
  AND2_X1 _35486_ (
    .A1(_00008_[2]),
    .A2(_27344_),
    .ZN(_27345_)
  );
  AND2_X1 _35487_ (
    .A1(_27342_),
    .A2(_27345_),
    .ZN(_27346_)
  );
  INV_X1 _35488_ (
    .A(_27346_),
    .ZN(_27347_)
  );
  AND2_X1 _35489_ (
    .A1(\cpuregs[3] [25]),
    .A2(_00008_[0]),
    .ZN(_27348_)
  );
  INV_X1 _35490_ (
    .A(_27348_),
    .ZN(_27349_)
  );
  AND2_X1 _35491_ (
    .A1(\cpuregs[2] [25]),
    .A2(_22147_),
    .ZN(_27350_)
  );
  INV_X1 _35492_ (
    .A(_27350_),
    .ZN(_27351_)
  );
  AND2_X1 _35493_ (
    .A1(_22149_),
    .A2(_27351_),
    .ZN(_27352_)
  );
  AND2_X1 _35494_ (
    .A1(_27349_),
    .A2(_27352_),
    .ZN(_27353_)
  );
  INV_X1 _35495_ (
    .A(_27353_),
    .ZN(_27354_)
  );
  AND2_X1 _35496_ (
    .A1(_22150_),
    .A2(_27354_),
    .ZN(_27355_)
  );
  AND2_X1 _35497_ (
    .A1(_27347_),
    .A2(_27355_),
    .ZN(_27356_)
  );
  INV_X1 _35498_ (
    .A(_27356_),
    .ZN(_27357_)
  );
  AND2_X1 _35499_ (
    .A1(\cpuregs[15] [25]),
    .A2(_00008_[0]),
    .ZN(_27358_)
  );
  INV_X1 _35500_ (
    .A(_27358_),
    .ZN(_27359_)
  );
  AND2_X1 _35501_ (
    .A1(\cpuregs[14] [25]),
    .A2(_22147_),
    .ZN(_27360_)
  );
  INV_X1 _35502_ (
    .A(_27360_),
    .ZN(_27361_)
  );
  AND2_X1 _35503_ (
    .A1(_00008_[2]),
    .A2(_27361_),
    .ZN(_27362_)
  );
  AND2_X1 _35504_ (
    .A1(_27359_),
    .A2(_27362_),
    .ZN(_27363_)
  );
  INV_X1 _35505_ (
    .A(_27363_),
    .ZN(_27364_)
  );
  AND2_X1 _35506_ (
    .A1(\cpuregs[11] [25]),
    .A2(_00008_[0]),
    .ZN(_27365_)
  );
  INV_X1 _35507_ (
    .A(_27365_),
    .ZN(_27366_)
  );
  AND2_X1 _35508_ (
    .A1(\cpuregs[10] [25]),
    .A2(_22147_),
    .ZN(_27367_)
  );
  INV_X1 _35509_ (
    .A(_27367_),
    .ZN(_27368_)
  );
  AND2_X1 _35510_ (
    .A1(_22149_),
    .A2(_27368_),
    .ZN(_27369_)
  );
  AND2_X1 _35511_ (
    .A1(_27366_),
    .A2(_27369_),
    .ZN(_27370_)
  );
  INV_X1 _35512_ (
    .A(_27370_),
    .ZN(_27371_)
  );
  AND2_X1 _35513_ (
    .A1(_00008_[3]),
    .A2(_27371_),
    .ZN(_27372_)
  );
  AND2_X1 _35514_ (
    .A1(_27364_),
    .A2(_27372_),
    .ZN(_27373_)
  );
  INV_X1 _35515_ (
    .A(_27373_),
    .ZN(_27374_)
  );
  AND2_X1 _35516_ (
    .A1(_27357_),
    .A2(_27374_),
    .ZN(_27375_)
  );
  INV_X1 _35517_ (
    .A(_27375_),
    .ZN(_27376_)
  );
  AND2_X1 _35518_ (
    .A1(_00008_[1]),
    .A2(_27376_),
    .ZN(_27377_)
  );
  INV_X1 _35519_ (
    .A(_27377_),
    .ZN(_27378_)
  );
  AND2_X1 _35520_ (
    .A1(_27340_),
    .A2(_27378_),
    .ZN(_27379_)
  );
  AND2_X1 _35521_ (
    .A1(_22151_),
    .A2(_27379_),
    .ZN(_27380_)
  );
  INV_X1 _35522_ (
    .A(_27380_),
    .ZN(_27381_)
  );
  AND2_X1 _35523_ (
    .A1(\cpuregs[26] [25]),
    .A2(_22149_),
    .ZN(_27382_)
  );
  INV_X1 _35524_ (
    .A(_27382_),
    .ZN(_27383_)
  );
  AND2_X1 _35525_ (
    .A1(\cpuregs[30] [25]),
    .A2(_00008_[2]),
    .ZN(_27384_)
  );
  INV_X1 _35526_ (
    .A(_27384_),
    .ZN(_27385_)
  );
  AND2_X1 _35527_ (
    .A1(_22147_),
    .A2(_27385_),
    .ZN(_27386_)
  );
  AND2_X1 _35528_ (
    .A1(_27383_),
    .A2(_27386_),
    .ZN(_27387_)
  );
  INV_X1 _35529_ (
    .A(_27387_),
    .ZN(_27388_)
  );
  AND2_X1 _35530_ (
    .A1(\cpuregs[31] [25]),
    .A2(_00008_[2]),
    .ZN(_27389_)
  );
  INV_X1 _35531_ (
    .A(_27389_),
    .ZN(_27390_)
  );
  AND2_X1 _35532_ (
    .A1(\cpuregs[27] [25]),
    .A2(_22149_),
    .ZN(_27391_)
  );
  INV_X1 _35533_ (
    .A(_27391_),
    .ZN(_27392_)
  );
  AND2_X1 _35534_ (
    .A1(_00008_[0]),
    .A2(_27392_),
    .ZN(_27393_)
  );
  AND2_X1 _35535_ (
    .A1(_27390_),
    .A2(_27393_),
    .ZN(_27394_)
  );
  INV_X1 _35536_ (
    .A(_27394_),
    .ZN(_27395_)
  );
  AND2_X1 _35537_ (
    .A1(_27388_),
    .A2(_27395_),
    .ZN(_27396_)
  );
  AND2_X1 _35538_ (
    .A1(\cpuregs[18] [25]),
    .A2(_22149_),
    .ZN(_27397_)
  );
  INV_X1 _35539_ (
    .A(_27397_),
    .ZN(_27398_)
  );
  AND2_X1 _35540_ (
    .A1(\cpuregs[22] [25]),
    .A2(_00008_[2]),
    .ZN(_27399_)
  );
  INV_X1 _35541_ (
    .A(_27399_),
    .ZN(_27400_)
  );
  AND2_X1 _35542_ (
    .A1(_22147_),
    .A2(_27400_),
    .ZN(_27401_)
  );
  AND2_X1 _35543_ (
    .A1(_27398_),
    .A2(_27401_),
    .ZN(_27402_)
  );
  INV_X1 _35544_ (
    .A(_27402_),
    .ZN(_27403_)
  );
  AND2_X1 _35545_ (
    .A1(\cpuregs[19] [25]),
    .A2(_22149_),
    .ZN(_27404_)
  );
  INV_X1 _35546_ (
    .A(_27404_),
    .ZN(_27405_)
  );
  AND2_X1 _35547_ (
    .A1(\cpuregs[23] [25]),
    .A2(_00008_[2]),
    .ZN(_27406_)
  );
  INV_X1 _35548_ (
    .A(_27406_),
    .ZN(_27407_)
  );
  AND2_X1 _35549_ (
    .A1(_00008_[0]),
    .A2(_27407_),
    .ZN(_27408_)
  );
  AND2_X1 _35550_ (
    .A1(_27405_),
    .A2(_27408_),
    .ZN(_27409_)
  );
  INV_X1 _35551_ (
    .A(_27409_),
    .ZN(_27410_)
  );
  AND2_X1 _35552_ (
    .A1(_00008_[3]),
    .A2(_27396_),
    .ZN(_27411_)
  );
  INV_X1 _35553_ (
    .A(_27411_),
    .ZN(_27412_)
  );
  AND2_X1 _35554_ (
    .A1(_22150_),
    .A2(_27410_),
    .ZN(_27413_)
  );
  AND2_X1 _35555_ (
    .A1(_27403_),
    .A2(_27413_),
    .ZN(_27414_)
  );
  INV_X1 _35556_ (
    .A(_27414_),
    .ZN(_27415_)
  );
  AND2_X1 _35557_ (
    .A1(_27412_),
    .A2(_27415_),
    .ZN(_27416_)
  );
  AND2_X1 _35558_ (
    .A1(_00008_[1]),
    .A2(_27416_),
    .ZN(_27417_)
  );
  INV_X1 _35559_ (
    .A(_27417_),
    .ZN(_27418_)
  );
  AND2_X1 _35560_ (
    .A1(\cpuregs[24] [25]),
    .A2(_22149_),
    .ZN(_27419_)
  );
  INV_X1 _35561_ (
    .A(_27419_),
    .ZN(_27420_)
  );
  AND2_X1 _35562_ (
    .A1(\cpuregs[28] [25]),
    .A2(_00008_[2]),
    .ZN(_27421_)
  );
  INV_X1 _35563_ (
    .A(_27421_),
    .ZN(_27422_)
  );
  AND2_X1 _35564_ (
    .A1(_22147_),
    .A2(_27422_),
    .ZN(_27423_)
  );
  AND2_X1 _35565_ (
    .A1(_27420_),
    .A2(_27423_),
    .ZN(_27424_)
  );
  INV_X1 _35566_ (
    .A(_27424_),
    .ZN(_27425_)
  );
  AND2_X1 _35567_ (
    .A1(\cpuregs[29] [25]),
    .A2(_00008_[2]),
    .ZN(_27426_)
  );
  INV_X1 _35568_ (
    .A(_27426_),
    .ZN(_27427_)
  );
  AND2_X1 _35569_ (
    .A1(\cpuregs[25] [25]),
    .A2(_22149_),
    .ZN(_27428_)
  );
  INV_X1 _35570_ (
    .A(_27428_),
    .ZN(_27429_)
  );
  AND2_X1 _35571_ (
    .A1(_00008_[0]),
    .A2(_27429_),
    .ZN(_27430_)
  );
  AND2_X1 _35572_ (
    .A1(_27427_),
    .A2(_27430_),
    .ZN(_27431_)
  );
  INV_X1 _35573_ (
    .A(_27431_),
    .ZN(_27432_)
  );
  AND2_X1 _35574_ (
    .A1(_27425_),
    .A2(_27432_),
    .ZN(_27433_)
  );
  AND2_X1 _35575_ (
    .A1(\cpuregs[16] [25]),
    .A2(_22149_),
    .ZN(_27434_)
  );
  INV_X1 _35576_ (
    .A(_27434_),
    .ZN(_27435_)
  );
  AND2_X1 _35577_ (
    .A1(\cpuregs[20] [25]),
    .A2(_00008_[2]),
    .ZN(_27436_)
  );
  INV_X1 _35578_ (
    .A(_27436_),
    .ZN(_27437_)
  );
  AND2_X1 _35579_ (
    .A1(_22147_),
    .A2(_27437_),
    .ZN(_27438_)
  );
  AND2_X1 _35580_ (
    .A1(_27435_),
    .A2(_27438_),
    .ZN(_27439_)
  );
  INV_X1 _35581_ (
    .A(_27439_),
    .ZN(_27440_)
  );
  AND2_X1 _35582_ (
    .A1(\cpuregs[17] [25]),
    .A2(_22149_),
    .ZN(_27441_)
  );
  INV_X1 _35583_ (
    .A(_27441_),
    .ZN(_27442_)
  );
  AND2_X1 _35584_ (
    .A1(\cpuregs[21] [25]),
    .A2(_00008_[2]),
    .ZN(_27443_)
  );
  INV_X1 _35585_ (
    .A(_27443_),
    .ZN(_27444_)
  );
  AND2_X1 _35586_ (
    .A1(_00008_[0]),
    .A2(_27444_),
    .ZN(_27445_)
  );
  AND2_X1 _35587_ (
    .A1(_27442_),
    .A2(_27445_),
    .ZN(_27446_)
  );
  INV_X1 _35588_ (
    .A(_27446_),
    .ZN(_27447_)
  );
  AND2_X1 _35589_ (
    .A1(_00008_[3]),
    .A2(_27433_),
    .ZN(_27448_)
  );
  INV_X1 _35590_ (
    .A(_27448_),
    .ZN(_27449_)
  );
  AND2_X1 _35591_ (
    .A1(_22150_),
    .A2(_27447_),
    .ZN(_27450_)
  );
  AND2_X1 _35592_ (
    .A1(_27440_),
    .A2(_27450_),
    .ZN(_27451_)
  );
  INV_X1 _35593_ (
    .A(_27451_),
    .ZN(_27452_)
  );
  AND2_X1 _35594_ (
    .A1(_27449_),
    .A2(_27452_),
    .ZN(_27453_)
  );
  AND2_X1 _35595_ (
    .A1(_22148_),
    .A2(_27453_),
    .ZN(_27454_)
  );
  INV_X1 _35596_ (
    .A(_27454_),
    .ZN(_27455_)
  );
  AND2_X1 _35597_ (
    .A1(_27418_),
    .A2(_27455_),
    .ZN(_27456_)
  );
  INV_X1 _35598_ (
    .A(_27456_),
    .ZN(_27457_)
  );
  AND2_X1 _35599_ (
    .A1(_00008_[4]),
    .A2(_27457_),
    .ZN(_27458_)
  );
  INV_X1 _35600_ (
    .A(_27458_),
    .ZN(_27459_)
  );
  AND2_X1 _35601_ (
    .A1(_22546_),
    .A2(_27459_),
    .ZN(_27460_)
  );
  AND2_X1 _35602_ (
    .A1(_27381_),
    .A2(_27460_),
    .ZN(_27461_)
  );
  INV_X1 _35603_ (
    .A(_27461_),
    .ZN(_27462_)
  );
  AND2_X1 _35604_ (
    .A1(_27300_),
    .A2(_27462_),
    .ZN(_27463_)
  );
  INV_X1 _35605_ (
    .A(_27463_),
    .ZN(_27464_)
  );
  AND2_X1 _35606_ (
    .A1(_22271_),
    .A2(_27464_),
    .ZN(_27465_)
  );
  INV_X1 _35607_ (
    .A(_27465_),
    .ZN(_27466_)
  );
  AND2_X1 _35608_ (
    .A1(reg_op1[24]),
    .A2(_22285_),
    .ZN(_27467_)
  );
  INV_X1 _35609_ (
    .A(_27467_),
    .ZN(_27468_)
  );
  AND2_X1 _35610_ (
    .A1(_26861_),
    .A2(_27468_),
    .ZN(_27469_)
  );
  AND2_X1 _35611_ (
    .A1(reg_op1[29]),
    .A2(_22290_),
    .ZN(_27470_)
  );
  INV_X1 _35612_ (
    .A(_27470_),
    .ZN(_27471_)
  );
  AND2_X1 _35613_ (
    .A1(_26858_),
    .A2(_27471_),
    .ZN(_27472_)
  );
  AND2_X1 _35614_ (
    .A1(_22572_),
    .A2(_27469_),
    .ZN(_27473_)
  );
  INV_X1 _35615_ (
    .A(_27473_),
    .ZN(_27474_)
  );
  AND2_X1 _35616_ (
    .A1(_22573_),
    .A2(_27472_),
    .ZN(_27475_)
  );
  INV_X1 _35617_ (
    .A(_27475_),
    .ZN(_27476_)
  );
  AND2_X1 _35618_ (
    .A1(_22295_),
    .A2(_27476_),
    .ZN(_27477_)
  );
  AND2_X1 _35619_ (
    .A1(_27474_),
    .A2(_27477_),
    .ZN(_27478_)
  );
  INV_X1 _35620_ (
    .A(_27478_),
    .ZN(_27479_)
  );
  AND2_X1 _35621_ (
    .A1(_22333_),
    .A2(_27479_),
    .ZN(_27480_)
  );
  AND2_X1 _35622_ (
    .A1(_27466_),
    .A2(_27480_),
    .ZN(_27481_)
  );
  AND2_X1 _35623_ (
    .A1(_27277_),
    .A2(_27289_),
    .ZN(_27482_)
  );
  INV_X1 _35624_ (
    .A(_27482_),
    .ZN(_27483_)
  );
  AND2_X1 _35625_ (
    .A1(reg_op1[25]),
    .A2(decoded_imm[25]),
    .ZN(_27484_)
  );
  INV_X1 _35626_ (
    .A(_27484_),
    .ZN(_27485_)
  );
  AND2_X1 _35627_ (
    .A1(_21192_),
    .A2(_21984_),
    .ZN(_27486_)
  );
  INV_X1 _35628_ (
    .A(_27486_),
    .ZN(_27487_)
  );
  AND2_X1 _35629_ (
    .A1(_27485_),
    .A2(_27487_),
    .ZN(_27488_)
  );
  INV_X1 _35630_ (
    .A(_27488_),
    .ZN(_27489_)
  );
  AND2_X1 _35631_ (
    .A1(_27483_),
    .A2(_27488_),
    .ZN(_27490_)
  );
  INV_X1 _35632_ (
    .A(_27490_),
    .ZN(_27491_)
  );
  AND2_X1 _35633_ (
    .A1(_27482_),
    .A2(_27489_),
    .ZN(_27492_)
  );
  INV_X1 _35634_ (
    .A(_27492_),
    .ZN(_27493_)
  );
  AND2_X1 _35635_ (
    .A1(_22559_),
    .A2(_27493_),
    .ZN(_27494_)
  );
  AND2_X1 _35636_ (
    .A1(_27491_),
    .A2(_27494_),
    .ZN(_27495_)
  );
  INV_X1 _35637_ (
    .A(_27495_),
    .ZN(_27496_)
  );
  AND2_X1 _35638_ (
    .A1(_27481_),
    .A2(_27496_),
    .ZN(_27497_)
  );
  INV_X1 _35639_ (
    .A(_27497_),
    .ZN(_27498_)
  );
  AND2_X1 _35640_ (
    .A1(_27298_),
    .A2(_27498_),
    .ZN(_00082_)
  );
  AND2_X1 _35641_ (
    .A1(_21193_),
    .A2(_22334_),
    .ZN(_27499_)
  );
  INV_X1 _35642_ (
    .A(_27499_),
    .ZN(_27500_)
  );
  AND2_X1 _35643_ (
    .A1(reg_pc[26]),
    .A2(_22335_),
    .ZN(_27501_)
  );
  INV_X1 _35644_ (
    .A(_27501_),
    .ZN(_27502_)
  );
  AND2_X1 _35645_ (
    .A1(_21799_),
    .A2(_00008_[2]),
    .ZN(_27503_)
  );
  INV_X1 _35646_ (
    .A(_27503_),
    .ZN(_27504_)
  );
  AND2_X1 _35647_ (
    .A1(_21507_),
    .A2(_22149_),
    .ZN(_27505_)
  );
  INV_X1 _35648_ (
    .A(_27505_),
    .ZN(_27506_)
  );
  AND2_X1 _35649_ (
    .A1(_00008_[0]),
    .A2(_27506_),
    .ZN(_27507_)
  );
  AND2_X1 _35650_ (
    .A1(_27504_),
    .A2(_27507_),
    .ZN(_27508_)
  );
  INV_X1 _35651_ (
    .A(_27508_),
    .ZN(_27509_)
  );
  AND2_X1 _35652_ (
    .A1(_21562_),
    .A2(_22149_),
    .ZN(_27510_)
  );
  INV_X1 _35653_ (
    .A(_27510_),
    .ZN(_27511_)
  );
  AND2_X1 _35654_ (
    .A1(_21828_),
    .A2(_00008_[2]),
    .ZN(_27512_)
  );
  INV_X1 _35655_ (
    .A(_27512_),
    .ZN(_27513_)
  );
  AND2_X1 _35656_ (
    .A1(_27511_),
    .A2(_27513_),
    .ZN(_27514_)
  );
  AND2_X1 _35657_ (
    .A1(_22147_),
    .A2(_27514_),
    .ZN(_27515_)
  );
  INV_X1 _35658_ (
    .A(_27515_),
    .ZN(_27516_)
  );
  AND2_X1 _35659_ (
    .A1(_27509_),
    .A2(_27516_),
    .ZN(_27517_)
  );
  AND2_X1 _35660_ (
    .A1(_21752_),
    .A2(_00008_[2]),
    .ZN(_27518_)
  );
  INV_X1 _35661_ (
    .A(_27518_),
    .ZN(_27519_)
  );
  AND2_X1 _35662_ (
    .A1(_21532_),
    .A2(_22149_),
    .ZN(_27520_)
  );
  INV_X1 _35663_ (
    .A(_27520_),
    .ZN(_27521_)
  );
  AND2_X1 _35664_ (
    .A1(_00008_[0]),
    .A2(_27519_),
    .ZN(_27522_)
  );
  AND2_X1 _35665_ (
    .A1(_27521_),
    .A2(_27522_),
    .ZN(_27523_)
  );
  INV_X1 _35666_ (
    .A(_27523_),
    .ZN(_27524_)
  );
  AND2_X1 _35667_ (
    .A1(_21973_),
    .A2(_22149_),
    .ZN(_27525_)
  );
  INV_X1 _35668_ (
    .A(_27525_),
    .ZN(_27526_)
  );
  AND2_X1 _35669_ (
    .A1(_21689_),
    .A2(_00008_[2]),
    .ZN(_27527_)
  );
  INV_X1 _35670_ (
    .A(_27527_),
    .ZN(_27528_)
  );
  AND2_X1 _35671_ (
    .A1(_27526_),
    .A2(_27528_),
    .ZN(_27529_)
  );
  AND2_X1 _35672_ (
    .A1(_22147_),
    .A2(_27529_),
    .ZN(_27530_)
  );
  INV_X1 _35673_ (
    .A(_27530_),
    .ZN(_27531_)
  );
  AND2_X1 _35674_ (
    .A1(_27524_),
    .A2(_27531_),
    .ZN(_27532_)
  );
  AND2_X1 _35675_ (
    .A1(_00008_[1]),
    .A2(_27517_),
    .ZN(_27533_)
  );
  INV_X1 _35676_ (
    .A(_27533_),
    .ZN(_27534_)
  );
  AND2_X1 _35677_ (
    .A1(_22148_),
    .A2(_27532_),
    .ZN(_27535_)
  );
  INV_X1 _35678_ (
    .A(_27535_),
    .ZN(_27536_)
  );
  AND2_X1 _35679_ (
    .A1(_22150_),
    .A2(_27536_),
    .ZN(_27537_)
  );
  AND2_X1 _35680_ (
    .A1(_27534_),
    .A2(_27537_),
    .ZN(_27538_)
  );
  INV_X1 _35681_ (
    .A(_27538_),
    .ZN(_27539_)
  );
  AND2_X1 _35682_ (
    .A1(\cpuregs[13] [26]),
    .A2(_00008_[0]),
    .ZN(_27540_)
  );
  INV_X1 _35683_ (
    .A(_27540_),
    .ZN(_27541_)
  );
  AND2_X1 _35684_ (
    .A1(\cpuregs[12] [26]),
    .A2(_22147_),
    .ZN(_27542_)
  );
  INV_X1 _35685_ (
    .A(_27542_),
    .ZN(_27543_)
  );
  AND2_X1 _35686_ (
    .A1(_00008_[2]),
    .A2(_27543_),
    .ZN(_27544_)
  );
  AND2_X1 _35687_ (
    .A1(_27541_),
    .A2(_27544_),
    .ZN(_27545_)
  );
  INV_X1 _35688_ (
    .A(_27545_),
    .ZN(_27546_)
  );
  AND2_X1 _35689_ (
    .A1(\cpuregs[9] [26]),
    .A2(_00008_[0]),
    .ZN(_27547_)
  );
  INV_X1 _35690_ (
    .A(_27547_),
    .ZN(_27548_)
  );
  AND2_X1 _35691_ (
    .A1(\cpuregs[8] [26]),
    .A2(_22147_),
    .ZN(_27549_)
  );
  INV_X1 _35692_ (
    .A(_27549_),
    .ZN(_27550_)
  );
  AND2_X1 _35693_ (
    .A1(_22149_),
    .A2(_27550_),
    .ZN(_27551_)
  );
  AND2_X1 _35694_ (
    .A1(_27548_),
    .A2(_27551_),
    .ZN(_27552_)
  );
  INV_X1 _35695_ (
    .A(_27552_),
    .ZN(_27553_)
  );
  AND2_X1 _35696_ (
    .A1(_22148_),
    .A2(_27553_),
    .ZN(_27554_)
  );
  AND2_X1 _35697_ (
    .A1(_27546_),
    .A2(_27554_),
    .ZN(_27555_)
  );
  INV_X1 _35698_ (
    .A(_27555_),
    .ZN(_27556_)
  );
  AND2_X1 _35699_ (
    .A1(\cpuregs[15] [26]),
    .A2(_00008_[0]),
    .ZN(_27557_)
  );
  INV_X1 _35700_ (
    .A(_27557_),
    .ZN(_27558_)
  );
  AND2_X1 _35701_ (
    .A1(\cpuregs[14] [26]),
    .A2(_22147_),
    .ZN(_27559_)
  );
  INV_X1 _35702_ (
    .A(_27559_),
    .ZN(_27560_)
  );
  AND2_X1 _35703_ (
    .A1(_00008_[2]),
    .A2(_27560_),
    .ZN(_27561_)
  );
  AND2_X1 _35704_ (
    .A1(_27558_),
    .A2(_27561_),
    .ZN(_27562_)
  );
  INV_X1 _35705_ (
    .A(_27562_),
    .ZN(_27563_)
  );
  AND2_X1 _35706_ (
    .A1(\cpuregs[11] [26]),
    .A2(_00008_[0]),
    .ZN(_27564_)
  );
  INV_X1 _35707_ (
    .A(_27564_),
    .ZN(_27565_)
  );
  AND2_X1 _35708_ (
    .A1(\cpuregs[10] [26]),
    .A2(_22147_),
    .ZN(_27566_)
  );
  INV_X1 _35709_ (
    .A(_27566_),
    .ZN(_27567_)
  );
  AND2_X1 _35710_ (
    .A1(_22149_),
    .A2(_27567_),
    .ZN(_27568_)
  );
  AND2_X1 _35711_ (
    .A1(_27565_),
    .A2(_27568_),
    .ZN(_27569_)
  );
  INV_X1 _35712_ (
    .A(_27569_),
    .ZN(_27570_)
  );
  AND2_X1 _35713_ (
    .A1(_00008_[1]),
    .A2(_27570_),
    .ZN(_27571_)
  );
  AND2_X1 _35714_ (
    .A1(_27563_),
    .A2(_27571_),
    .ZN(_27572_)
  );
  INV_X1 _35715_ (
    .A(_27572_),
    .ZN(_27573_)
  );
  AND2_X1 _35716_ (
    .A1(_27556_),
    .A2(_27573_),
    .ZN(_27574_)
  );
  INV_X1 _35717_ (
    .A(_27574_),
    .ZN(_27575_)
  );
  AND2_X1 _35718_ (
    .A1(_00008_[3]),
    .A2(_27575_),
    .ZN(_27576_)
  );
  INV_X1 _35719_ (
    .A(_27576_),
    .ZN(_27577_)
  );
  AND2_X1 _35720_ (
    .A1(_22151_),
    .A2(_27539_),
    .ZN(_27578_)
  );
  AND2_X1 _35721_ (
    .A1(_27577_),
    .A2(_27578_),
    .ZN(_27579_)
  );
  INV_X1 _35722_ (
    .A(_27579_),
    .ZN(_27580_)
  );
  AND2_X1 _35723_ (
    .A1(\cpuregs[26] [26]),
    .A2(_22149_),
    .ZN(_27581_)
  );
  INV_X1 _35724_ (
    .A(_27581_),
    .ZN(_27582_)
  );
  AND2_X1 _35725_ (
    .A1(\cpuregs[30] [26]),
    .A2(_00008_[2]),
    .ZN(_27583_)
  );
  INV_X1 _35726_ (
    .A(_27583_),
    .ZN(_27584_)
  );
  AND2_X1 _35727_ (
    .A1(_22147_),
    .A2(_27584_),
    .ZN(_27585_)
  );
  AND2_X1 _35728_ (
    .A1(_27582_),
    .A2(_27585_),
    .ZN(_27586_)
  );
  INV_X1 _35729_ (
    .A(_27586_),
    .ZN(_27587_)
  );
  AND2_X1 _35730_ (
    .A1(\cpuregs[31] [26]),
    .A2(_00008_[2]),
    .ZN(_27588_)
  );
  INV_X1 _35731_ (
    .A(_27588_),
    .ZN(_27589_)
  );
  AND2_X1 _35732_ (
    .A1(\cpuregs[27] [26]),
    .A2(_22149_),
    .ZN(_27590_)
  );
  INV_X1 _35733_ (
    .A(_27590_),
    .ZN(_27591_)
  );
  AND2_X1 _35734_ (
    .A1(_00008_[0]),
    .A2(_27591_),
    .ZN(_27592_)
  );
  AND2_X1 _35735_ (
    .A1(_27589_),
    .A2(_27592_),
    .ZN(_27593_)
  );
  INV_X1 _35736_ (
    .A(_27593_),
    .ZN(_27594_)
  );
  AND2_X1 _35737_ (
    .A1(_27587_),
    .A2(_27594_),
    .ZN(_27595_)
  );
  AND2_X1 _35738_ (
    .A1(\cpuregs[18] [26]),
    .A2(_22149_),
    .ZN(_27596_)
  );
  INV_X1 _35739_ (
    .A(_27596_),
    .ZN(_27597_)
  );
  AND2_X1 _35740_ (
    .A1(\cpuregs[22] [26]),
    .A2(_00008_[2]),
    .ZN(_27598_)
  );
  INV_X1 _35741_ (
    .A(_27598_),
    .ZN(_27599_)
  );
  AND2_X1 _35742_ (
    .A1(_22147_),
    .A2(_27599_),
    .ZN(_27600_)
  );
  AND2_X1 _35743_ (
    .A1(_27597_),
    .A2(_27600_),
    .ZN(_27601_)
  );
  INV_X1 _35744_ (
    .A(_27601_),
    .ZN(_27602_)
  );
  AND2_X1 _35745_ (
    .A1(\cpuregs[19] [26]),
    .A2(_22149_),
    .ZN(_27603_)
  );
  INV_X1 _35746_ (
    .A(_27603_),
    .ZN(_27604_)
  );
  AND2_X1 _35747_ (
    .A1(\cpuregs[23] [26]),
    .A2(_00008_[2]),
    .ZN(_27605_)
  );
  INV_X1 _35748_ (
    .A(_27605_),
    .ZN(_27606_)
  );
  AND2_X1 _35749_ (
    .A1(_00008_[0]),
    .A2(_27606_),
    .ZN(_27607_)
  );
  AND2_X1 _35750_ (
    .A1(_27604_),
    .A2(_27607_),
    .ZN(_27608_)
  );
  INV_X1 _35751_ (
    .A(_27608_),
    .ZN(_27609_)
  );
  AND2_X1 _35752_ (
    .A1(_00008_[3]),
    .A2(_27595_),
    .ZN(_27610_)
  );
  INV_X1 _35753_ (
    .A(_27610_),
    .ZN(_27611_)
  );
  AND2_X1 _35754_ (
    .A1(_22150_),
    .A2(_27609_),
    .ZN(_27612_)
  );
  AND2_X1 _35755_ (
    .A1(_27602_),
    .A2(_27612_),
    .ZN(_27613_)
  );
  INV_X1 _35756_ (
    .A(_27613_),
    .ZN(_27614_)
  );
  AND2_X1 _35757_ (
    .A1(_27611_),
    .A2(_27614_),
    .ZN(_27615_)
  );
  AND2_X1 _35758_ (
    .A1(_00008_[1]),
    .A2(_27615_),
    .ZN(_27616_)
  );
  INV_X1 _35759_ (
    .A(_27616_),
    .ZN(_27617_)
  );
  AND2_X1 _35760_ (
    .A1(\cpuregs[24] [26]),
    .A2(_22149_),
    .ZN(_27618_)
  );
  INV_X1 _35761_ (
    .A(_27618_),
    .ZN(_27619_)
  );
  AND2_X1 _35762_ (
    .A1(\cpuregs[28] [26]),
    .A2(_00008_[2]),
    .ZN(_27620_)
  );
  INV_X1 _35763_ (
    .A(_27620_),
    .ZN(_27621_)
  );
  AND2_X1 _35764_ (
    .A1(_22147_),
    .A2(_27621_),
    .ZN(_27622_)
  );
  AND2_X1 _35765_ (
    .A1(_27619_),
    .A2(_27622_),
    .ZN(_01576_)
  );
  INV_X1 _35766_ (
    .A(_01576_),
    .ZN(_01577_)
  );
  AND2_X1 _35767_ (
    .A1(\cpuregs[29] [26]),
    .A2(_00008_[2]),
    .ZN(_01578_)
  );
  INV_X1 _35768_ (
    .A(_01578_),
    .ZN(_01579_)
  );
  AND2_X1 _35769_ (
    .A1(\cpuregs[25] [26]),
    .A2(_22149_),
    .ZN(_01580_)
  );
  INV_X1 _35770_ (
    .A(_01580_),
    .ZN(_01581_)
  );
  AND2_X1 _35771_ (
    .A1(_00008_[0]),
    .A2(_01581_),
    .ZN(_01582_)
  );
  AND2_X1 _35772_ (
    .A1(_01579_),
    .A2(_01582_),
    .ZN(_01583_)
  );
  INV_X1 _35773_ (
    .A(_01583_),
    .ZN(_01584_)
  );
  AND2_X1 _35774_ (
    .A1(_01577_),
    .A2(_01584_),
    .ZN(_01585_)
  );
  AND2_X1 _35775_ (
    .A1(\cpuregs[16] [26]),
    .A2(_22149_),
    .ZN(_01586_)
  );
  INV_X1 _35776_ (
    .A(_01586_),
    .ZN(_01587_)
  );
  AND2_X1 _35777_ (
    .A1(\cpuregs[20] [26]),
    .A2(_00008_[2]),
    .ZN(_01588_)
  );
  INV_X1 _35778_ (
    .A(_01588_),
    .ZN(_01589_)
  );
  AND2_X1 _35779_ (
    .A1(_22147_),
    .A2(_01589_),
    .ZN(_01590_)
  );
  AND2_X1 _35780_ (
    .A1(_01587_),
    .A2(_01590_),
    .ZN(_01591_)
  );
  INV_X1 _35781_ (
    .A(_01591_),
    .ZN(_01592_)
  );
  AND2_X1 _35782_ (
    .A1(\cpuregs[17] [26]),
    .A2(_22149_),
    .ZN(_01593_)
  );
  INV_X1 _35783_ (
    .A(_01593_),
    .ZN(_01594_)
  );
  AND2_X1 _35784_ (
    .A1(\cpuregs[21] [26]),
    .A2(_00008_[2]),
    .ZN(_01595_)
  );
  INV_X1 _35785_ (
    .A(_01595_),
    .ZN(_01596_)
  );
  AND2_X1 _35786_ (
    .A1(_00008_[0]),
    .A2(_01596_),
    .ZN(_01597_)
  );
  AND2_X1 _35787_ (
    .A1(_01594_),
    .A2(_01597_),
    .ZN(_01598_)
  );
  INV_X1 _35788_ (
    .A(_01598_),
    .ZN(_01599_)
  );
  AND2_X1 _35789_ (
    .A1(_00008_[3]),
    .A2(_01585_),
    .ZN(_01600_)
  );
  INV_X1 _35790_ (
    .A(_01600_),
    .ZN(_01601_)
  );
  AND2_X1 _35791_ (
    .A1(_22150_),
    .A2(_01599_),
    .ZN(_01602_)
  );
  AND2_X1 _35792_ (
    .A1(_01592_),
    .A2(_01602_),
    .ZN(_01603_)
  );
  INV_X1 _35793_ (
    .A(_01603_),
    .ZN(_01604_)
  );
  AND2_X1 _35794_ (
    .A1(_01601_),
    .A2(_01604_),
    .ZN(_01605_)
  );
  AND2_X1 _35795_ (
    .A1(_22148_),
    .A2(_01605_),
    .ZN(_01606_)
  );
  INV_X1 _35796_ (
    .A(_01606_),
    .ZN(_01607_)
  );
  AND2_X1 _35797_ (
    .A1(_27617_),
    .A2(_01607_),
    .ZN(_01608_)
  );
  INV_X1 _35798_ (
    .A(_01608_),
    .ZN(_01609_)
  );
  AND2_X1 _35799_ (
    .A1(_00008_[4]),
    .A2(_01609_),
    .ZN(_01610_)
  );
  INV_X1 _35800_ (
    .A(_01610_),
    .ZN(_01611_)
  );
  AND2_X1 _35801_ (
    .A1(_22546_),
    .A2(_01611_),
    .ZN(_01612_)
  );
  AND2_X1 _35802_ (
    .A1(_27580_),
    .A2(_01612_),
    .ZN(_01613_)
  );
  INV_X1 _35803_ (
    .A(_01613_),
    .ZN(_01614_)
  );
  AND2_X1 _35804_ (
    .A1(_27502_),
    .A2(_01614_),
    .ZN(_01615_)
  );
  INV_X1 _35805_ (
    .A(_01615_),
    .ZN(_01616_)
  );
  AND2_X1 _35806_ (
    .A1(_22271_),
    .A2(_01616_),
    .ZN(_01617_)
  );
  INV_X1 _35807_ (
    .A(_01617_),
    .ZN(_01618_)
  );
  AND2_X1 _35808_ (
    .A1(reg_op1[25]),
    .A2(_22285_),
    .ZN(_01619_)
  );
  INV_X1 _35809_ (
    .A(_01619_),
    .ZN(_01620_)
  );
  AND2_X1 _35810_ (
    .A1(_27079_),
    .A2(_01620_),
    .ZN(_01621_)
  );
  AND2_X1 _35811_ (
    .A1(reg_op1[30]),
    .A2(_22290_),
    .ZN(_01622_)
  );
  INV_X1 _35812_ (
    .A(_01622_),
    .ZN(_01623_)
  );
  AND2_X1 _35813_ (
    .A1(_27073_),
    .A2(_01623_),
    .ZN(_01624_)
  );
  AND2_X1 _35814_ (
    .A1(_22572_),
    .A2(_01621_),
    .ZN(_01625_)
  );
  INV_X1 _35815_ (
    .A(_01625_),
    .ZN(_01626_)
  );
  AND2_X1 _35816_ (
    .A1(_22573_),
    .A2(_01624_),
    .ZN(_01627_)
  );
  INV_X1 _35817_ (
    .A(_01627_),
    .ZN(_01628_)
  );
  AND2_X1 _35818_ (
    .A1(_22295_),
    .A2(_01628_),
    .ZN(_01629_)
  );
  AND2_X1 _35819_ (
    .A1(_01626_),
    .A2(_01629_),
    .ZN(_01630_)
  );
  INV_X1 _35820_ (
    .A(_01630_),
    .ZN(_01631_)
  );
  AND2_X1 _35821_ (
    .A1(_22333_),
    .A2(_01631_),
    .ZN(_01632_)
  );
  AND2_X1 _35822_ (
    .A1(_01618_),
    .A2(_01632_),
    .ZN(_01633_)
  );
  AND2_X1 _35823_ (
    .A1(reg_op1[26]),
    .A2(decoded_imm[26]),
    .ZN(_01634_)
  );
  INV_X1 _35824_ (
    .A(_01634_),
    .ZN(_01635_)
  );
  AND2_X1 _35825_ (
    .A1(_21193_),
    .A2(_21983_),
    .ZN(_01636_)
  );
  INV_X1 _35826_ (
    .A(_01636_),
    .ZN(_01637_)
  );
  AND2_X1 _35827_ (
    .A1(_01635_),
    .A2(_01637_),
    .ZN(_01638_)
  );
  INV_X1 _35828_ (
    .A(_01638_),
    .ZN(_01639_)
  );
  AND2_X1 _35829_ (
    .A1(_27483_),
    .A2(_27487_),
    .ZN(_01640_)
  );
  INV_X1 _35830_ (
    .A(_01640_),
    .ZN(_01641_)
  );
  AND2_X1 _35831_ (
    .A1(_27482_),
    .A2(_27485_),
    .ZN(_01642_)
  );
  INV_X1 _35832_ (
    .A(_01642_),
    .ZN(_01643_)
  );
  AND2_X1 _35833_ (
    .A1(_27485_),
    .A2(_01641_),
    .ZN(_01644_)
  );
  AND2_X1 _35834_ (
    .A1(_27487_),
    .A2(_01643_),
    .ZN(_01645_)
  );
  AND2_X1 _35835_ (
    .A1(_01638_),
    .A2(_01645_),
    .ZN(_01646_)
  );
  INV_X1 _35836_ (
    .A(_01646_),
    .ZN(_01647_)
  );
  AND2_X1 _35837_ (
    .A1(_01639_),
    .A2(_01644_),
    .ZN(_01648_)
  );
  INV_X1 _35838_ (
    .A(_01648_),
    .ZN(_01649_)
  );
  AND2_X1 _35839_ (
    .A1(_22559_),
    .A2(_01649_),
    .ZN(_01650_)
  );
  AND2_X1 _35840_ (
    .A1(_01647_),
    .A2(_01650_),
    .ZN(_01651_)
  );
  INV_X1 _35841_ (
    .A(_01651_),
    .ZN(_01652_)
  );
  AND2_X1 _35842_ (
    .A1(_01633_),
    .A2(_01652_),
    .ZN(_01653_)
  );
  INV_X1 _35843_ (
    .A(_01653_),
    .ZN(_01654_)
  );
  AND2_X1 _35844_ (
    .A1(_27500_),
    .A2(_01654_),
    .ZN(_00083_)
  );
  AND2_X1 _35845_ (
    .A1(_21194_),
    .A2(_22334_),
    .ZN(_01655_)
  );
  INV_X1 _35846_ (
    .A(_01655_),
    .ZN(_01656_)
  );
  AND2_X1 _35847_ (
    .A1(reg_pc[27]),
    .A2(_22335_),
    .ZN(_01657_)
  );
  INV_X1 _35848_ (
    .A(_01657_),
    .ZN(_01658_)
  );
  AND2_X1 _35849_ (
    .A1(\cpuregs[21] [27]),
    .A2(_00008_[2]),
    .ZN(_01659_)
  );
  INV_X1 _35850_ (
    .A(_01659_),
    .ZN(_01660_)
  );
  AND2_X1 _35851_ (
    .A1(\cpuregs[17] [27]),
    .A2(_22149_),
    .ZN(_01661_)
  );
  INV_X1 _35852_ (
    .A(_01661_),
    .ZN(_01662_)
  );
  AND2_X1 _35853_ (
    .A1(_01660_),
    .A2(_01662_),
    .ZN(_01663_)
  );
  INV_X1 _35854_ (
    .A(_01663_),
    .ZN(_01664_)
  );
  AND2_X1 _35855_ (
    .A1(_00008_[0]),
    .A2(_01664_),
    .ZN(_01665_)
  );
  INV_X1 _35856_ (
    .A(_01665_),
    .ZN(_01666_)
  );
  AND2_X1 _35857_ (
    .A1(\cpuregs[20] [27]),
    .A2(_00008_[2]),
    .ZN(_01667_)
  );
  INV_X1 _35858_ (
    .A(_01667_),
    .ZN(_01668_)
  );
  AND2_X1 _35859_ (
    .A1(\cpuregs[16] [27]),
    .A2(_22149_),
    .ZN(_01669_)
  );
  INV_X1 _35860_ (
    .A(_01669_),
    .ZN(_01670_)
  );
  AND2_X1 _35861_ (
    .A1(_01668_),
    .A2(_01670_),
    .ZN(_01671_)
  );
  INV_X1 _35862_ (
    .A(_01671_),
    .ZN(_01672_)
  );
  AND2_X1 _35863_ (
    .A1(_22147_),
    .A2(_01672_),
    .ZN(_01673_)
  );
  INV_X1 _35864_ (
    .A(_01673_),
    .ZN(_01674_)
  );
  AND2_X1 _35865_ (
    .A1(_01666_),
    .A2(_01674_),
    .ZN(_01675_)
  );
  AND2_X1 _35866_ (
    .A1(_21690_),
    .A2(_00008_[2]),
    .ZN(_01676_)
  );
  INV_X1 _35867_ (
    .A(_01676_),
    .ZN(_01677_)
  );
  AND2_X1 _35868_ (
    .A1(_21974_),
    .A2(_22149_),
    .ZN(_01678_)
  );
  INV_X1 _35869_ (
    .A(_01678_),
    .ZN(_01679_)
  );
  AND2_X1 _35870_ (
    .A1(_01677_),
    .A2(_01679_),
    .ZN(_01680_)
  );
  AND2_X1 _35871_ (
    .A1(_22147_),
    .A2(_01680_),
    .ZN(_01681_)
  );
  INV_X1 _35872_ (
    .A(_01681_),
    .ZN(_01682_)
  );
  AND2_X1 _35873_ (
    .A1(_21753_),
    .A2(_00008_[2]),
    .ZN(_01683_)
  );
  INV_X1 _35874_ (
    .A(_01683_),
    .ZN(_01684_)
  );
  AND2_X1 _35875_ (
    .A1(_21533_),
    .A2(_22149_),
    .ZN(_01685_)
  );
  INV_X1 _35876_ (
    .A(_01685_),
    .ZN(_01686_)
  );
  AND2_X1 _35877_ (
    .A1(_00008_[0]),
    .A2(_01686_),
    .ZN(_01687_)
  );
  AND2_X1 _35878_ (
    .A1(_01684_),
    .A2(_01687_),
    .ZN(_01688_)
  );
  INV_X1 _35879_ (
    .A(_01688_),
    .ZN(_01689_)
  );
  AND2_X1 _35880_ (
    .A1(_01682_),
    .A2(_01689_),
    .ZN(_01690_)
  );
  AND2_X1 _35881_ (
    .A1(\cpuregs[23] [27]),
    .A2(_00008_[2]),
    .ZN(_01691_)
  );
  INV_X1 _35882_ (
    .A(_01691_),
    .ZN(_01692_)
  );
  AND2_X1 _35883_ (
    .A1(\cpuregs[19] [27]),
    .A2(_22149_),
    .ZN(_01693_)
  );
  INV_X1 _35884_ (
    .A(_01693_),
    .ZN(_01694_)
  );
  AND2_X1 _35885_ (
    .A1(_01692_),
    .A2(_01694_),
    .ZN(_01695_)
  );
  INV_X1 _35886_ (
    .A(_01695_),
    .ZN(_01696_)
  );
  AND2_X1 _35887_ (
    .A1(_00008_[0]),
    .A2(_01696_),
    .ZN(_01697_)
  );
  INV_X1 _35888_ (
    .A(_01697_),
    .ZN(_01698_)
  );
  AND2_X1 _35889_ (
    .A1(_21612_),
    .A2(_22149_),
    .ZN(_01699_)
  );
  INV_X1 _35890_ (
    .A(_01699_),
    .ZN(_01700_)
  );
  AND2_X1 _35891_ (
    .A1(_21432_),
    .A2(_00008_[2]),
    .ZN(_01701_)
  );
  INV_X1 _35892_ (
    .A(_01701_),
    .ZN(_01702_)
  );
  AND2_X1 _35893_ (
    .A1(_01700_),
    .A2(_01702_),
    .ZN(_01703_)
  );
  AND2_X1 _35894_ (
    .A1(_22147_),
    .A2(_01703_),
    .ZN(_01704_)
  );
  INV_X1 _35895_ (
    .A(_01704_),
    .ZN(_01705_)
  );
  AND2_X1 _35896_ (
    .A1(_21829_),
    .A2(_00008_[2]),
    .ZN(_01706_)
  );
  INV_X1 _35897_ (
    .A(_01706_),
    .ZN(_01707_)
  );
  AND2_X1 _35898_ (
    .A1(_21563_),
    .A2(_22149_),
    .ZN(_01708_)
  );
  INV_X1 _35899_ (
    .A(_01708_),
    .ZN(_01709_)
  );
  AND2_X1 _35900_ (
    .A1(_01707_),
    .A2(_01709_),
    .ZN(_01710_)
  );
  AND2_X1 _35901_ (
    .A1(_22147_),
    .A2(_01710_),
    .ZN(_01711_)
  );
  INV_X1 _35902_ (
    .A(_01711_),
    .ZN(_01712_)
  );
  AND2_X1 _35903_ (
    .A1(_21800_),
    .A2(_00008_[2]),
    .ZN(_01713_)
  );
  INV_X1 _35904_ (
    .A(_01713_),
    .ZN(_01714_)
  );
  AND2_X1 _35905_ (
    .A1(_21508_),
    .A2(_22149_),
    .ZN(_01715_)
  );
  INV_X1 _35906_ (
    .A(_01715_),
    .ZN(_01716_)
  );
  AND2_X1 _35907_ (
    .A1(_00008_[0]),
    .A2(_01716_),
    .ZN(_01717_)
  );
  AND2_X1 _35908_ (
    .A1(_01714_),
    .A2(_01717_),
    .ZN(_01718_)
  );
  INV_X1 _35909_ (
    .A(_01718_),
    .ZN(_01719_)
  );
  AND2_X1 _35910_ (
    .A1(_01712_),
    .A2(_01719_),
    .ZN(_01720_)
  );
  AND2_X1 _35911_ (
    .A1(_00008_[1]),
    .A2(_01720_),
    .ZN(_01721_)
  );
  INV_X1 _35912_ (
    .A(_01721_),
    .ZN(_01722_)
  );
  AND2_X1 _35913_ (
    .A1(_22148_),
    .A2(_01690_),
    .ZN(_01723_)
  );
  INV_X1 _35914_ (
    .A(_01723_),
    .ZN(_01724_)
  );
  AND2_X1 _35915_ (
    .A1(_01722_),
    .A2(_01724_),
    .ZN(_01725_)
  );
  AND2_X1 _35916_ (
    .A1(_22151_),
    .A2(_01725_),
    .ZN(_01726_)
  );
  INV_X1 _35917_ (
    .A(_01726_),
    .ZN(_01727_)
  );
  AND2_X1 _35918_ (
    .A1(_00008_[1]),
    .A2(_01705_),
    .ZN(_01728_)
  );
  AND2_X1 _35919_ (
    .A1(_01698_),
    .A2(_01728_),
    .ZN(_01729_)
  );
  INV_X1 _35920_ (
    .A(_01729_),
    .ZN(_01730_)
  );
  AND2_X1 _35921_ (
    .A1(_22148_),
    .A2(_01675_),
    .ZN(_01731_)
  );
  INV_X1 _35922_ (
    .A(_01731_),
    .ZN(_01732_)
  );
  AND2_X1 _35923_ (
    .A1(_00008_[4]),
    .A2(_01732_),
    .ZN(_01733_)
  );
  AND2_X1 _35924_ (
    .A1(_01730_),
    .A2(_01733_),
    .ZN(_01734_)
  );
  INV_X1 _35925_ (
    .A(_01734_),
    .ZN(_01735_)
  );
  AND2_X1 _35926_ (
    .A1(_01727_),
    .A2(_01735_),
    .ZN(_01736_)
  );
  AND2_X1 _35927_ (
    .A1(_22150_),
    .A2(_01736_),
    .ZN(_01737_)
  );
  INV_X1 _35928_ (
    .A(_01737_),
    .ZN(_01738_)
  );
  AND2_X1 _35929_ (
    .A1(\cpuregs[29] [27]),
    .A2(_00008_[2]),
    .ZN(_01739_)
  );
  INV_X1 _35930_ (
    .A(_01739_),
    .ZN(_01740_)
  );
  AND2_X1 _35931_ (
    .A1(\cpuregs[25] [27]),
    .A2(_22149_),
    .ZN(_01741_)
  );
  INV_X1 _35932_ (
    .A(_01741_),
    .ZN(_01742_)
  );
  AND2_X1 _35933_ (
    .A1(_22148_),
    .A2(_01742_),
    .ZN(_01743_)
  );
  AND2_X1 _35934_ (
    .A1(_01740_),
    .A2(_01743_),
    .ZN(_01744_)
  );
  INV_X1 _35935_ (
    .A(_01744_),
    .ZN(_01745_)
  );
  AND2_X1 _35936_ (
    .A1(\cpuregs[27] [27]),
    .A2(_22149_),
    .ZN(_01746_)
  );
  INV_X1 _35937_ (
    .A(_01746_),
    .ZN(_01747_)
  );
  AND2_X1 _35938_ (
    .A1(\cpuregs[31] [27]),
    .A2(_00008_[2]),
    .ZN(_01748_)
  );
  INV_X1 _35939_ (
    .A(_01748_),
    .ZN(_01749_)
  );
  AND2_X1 _35940_ (
    .A1(_00008_[1]),
    .A2(_01749_),
    .ZN(_01750_)
  );
  AND2_X1 _35941_ (
    .A1(_01747_),
    .A2(_01750_),
    .ZN(_01751_)
  );
  INV_X1 _35942_ (
    .A(_01751_),
    .ZN(_01752_)
  );
  AND2_X1 _35943_ (
    .A1(_01745_),
    .A2(_01752_),
    .ZN(_01753_)
  );
  INV_X1 _35944_ (
    .A(_01753_),
    .ZN(_01754_)
  );
  AND2_X1 _35945_ (
    .A1(_00008_[0]),
    .A2(_01754_),
    .ZN(_01755_)
  );
  INV_X1 _35946_ (
    .A(_01755_),
    .ZN(_01756_)
  );
  AND2_X1 _35947_ (
    .A1(\cpuregs[24] [27]),
    .A2(_22149_),
    .ZN(_01757_)
  );
  INV_X1 _35948_ (
    .A(_01757_),
    .ZN(_01758_)
  );
  AND2_X1 _35949_ (
    .A1(\cpuregs[28] [27]),
    .A2(_00008_[2]),
    .ZN(_01759_)
  );
  INV_X1 _35950_ (
    .A(_01759_),
    .ZN(_01760_)
  );
  AND2_X1 _35951_ (
    .A1(_22148_),
    .A2(_01760_),
    .ZN(_01761_)
  );
  AND2_X1 _35952_ (
    .A1(_01758_),
    .A2(_01761_),
    .ZN(_01762_)
  );
  INV_X1 _35953_ (
    .A(_01762_),
    .ZN(_01763_)
  );
  AND2_X1 _35954_ (
    .A1(\cpuregs[26] [27]),
    .A2(_22149_),
    .ZN(_01764_)
  );
  INV_X1 _35955_ (
    .A(_01764_),
    .ZN(_01765_)
  );
  AND2_X1 _35956_ (
    .A1(\cpuregs[30] [27]),
    .A2(_00008_[2]),
    .ZN(_01766_)
  );
  INV_X1 _35957_ (
    .A(_01766_),
    .ZN(_01767_)
  );
  AND2_X1 _35958_ (
    .A1(_00008_[1]),
    .A2(_01767_),
    .ZN(_01768_)
  );
  AND2_X1 _35959_ (
    .A1(_01765_),
    .A2(_01768_),
    .ZN(_01769_)
  );
  INV_X1 _35960_ (
    .A(_01769_),
    .ZN(_01770_)
  );
  AND2_X1 _35961_ (
    .A1(_01763_),
    .A2(_01770_),
    .ZN(_01771_)
  );
  INV_X1 _35962_ (
    .A(_01771_),
    .ZN(_01772_)
  );
  AND2_X1 _35963_ (
    .A1(_22147_),
    .A2(_01772_),
    .ZN(_01773_)
  );
  INV_X1 _35964_ (
    .A(_01773_),
    .ZN(_01774_)
  );
  AND2_X1 _35965_ (
    .A1(_01756_),
    .A2(_01774_),
    .ZN(_01775_)
  );
  INV_X1 _35966_ (
    .A(_01775_),
    .ZN(_01776_)
  );
  AND2_X1 _35967_ (
    .A1(_00008_[4]),
    .A2(_01776_),
    .ZN(_01777_)
  );
  INV_X1 _35968_ (
    .A(_01777_),
    .ZN(_01778_)
  );
  AND2_X1 _35969_ (
    .A1(\cpuregs[9] [27]),
    .A2(_22148_),
    .ZN(_01779_)
  );
  INV_X1 _35970_ (
    .A(_01779_),
    .ZN(_01780_)
  );
  AND2_X1 _35971_ (
    .A1(\cpuregs[11] [27]),
    .A2(_00008_[1]),
    .ZN(_01781_)
  );
  INV_X1 _35972_ (
    .A(_01781_),
    .ZN(_01782_)
  );
  AND2_X1 _35973_ (
    .A1(_22149_),
    .A2(_01782_),
    .ZN(_01783_)
  );
  AND2_X1 _35974_ (
    .A1(_01780_),
    .A2(_01783_),
    .ZN(_01784_)
  );
  INV_X1 _35975_ (
    .A(_01784_),
    .ZN(_01785_)
  );
  AND2_X1 _35976_ (
    .A1(\cpuregs[13] [27]),
    .A2(_22148_),
    .ZN(_01786_)
  );
  INV_X1 _35977_ (
    .A(_01786_),
    .ZN(_01787_)
  );
  AND2_X1 _35978_ (
    .A1(\cpuregs[15] [27]),
    .A2(_00008_[1]),
    .ZN(_01788_)
  );
  INV_X1 _35979_ (
    .A(_01788_),
    .ZN(_01789_)
  );
  AND2_X1 _35980_ (
    .A1(_00008_[2]),
    .A2(_01789_),
    .ZN(_01790_)
  );
  AND2_X1 _35981_ (
    .A1(_01787_),
    .A2(_01790_),
    .ZN(_01791_)
  );
  INV_X1 _35982_ (
    .A(_01791_),
    .ZN(_01792_)
  );
  AND2_X1 _35983_ (
    .A1(_01785_),
    .A2(_01792_),
    .ZN(_01793_)
  );
  INV_X1 _35984_ (
    .A(_01793_),
    .ZN(_01794_)
  );
  AND2_X1 _35985_ (
    .A1(_00008_[0]),
    .A2(_01794_),
    .ZN(_01795_)
  );
  INV_X1 _35986_ (
    .A(_01795_),
    .ZN(_01796_)
  );
  AND2_X1 _35987_ (
    .A1(\cpuregs[8] [27]),
    .A2(_22148_),
    .ZN(_01797_)
  );
  INV_X1 _35988_ (
    .A(_01797_),
    .ZN(_01798_)
  );
  AND2_X1 _35989_ (
    .A1(\cpuregs[10] [27]),
    .A2(_00008_[1]),
    .ZN(_01799_)
  );
  INV_X1 _35990_ (
    .A(_01799_),
    .ZN(_01800_)
  );
  AND2_X1 _35991_ (
    .A1(_22149_),
    .A2(_01800_),
    .ZN(_01801_)
  );
  AND2_X1 _35992_ (
    .A1(_01798_),
    .A2(_01801_),
    .ZN(_01802_)
  );
  INV_X1 _35993_ (
    .A(_01802_),
    .ZN(_01803_)
  );
  AND2_X1 _35994_ (
    .A1(\cpuregs[12] [27]),
    .A2(_22148_),
    .ZN(_01804_)
  );
  INV_X1 _35995_ (
    .A(_01804_),
    .ZN(_01805_)
  );
  AND2_X1 _35996_ (
    .A1(\cpuregs[14] [27]),
    .A2(_00008_[1]),
    .ZN(_01806_)
  );
  INV_X1 _35997_ (
    .A(_01806_),
    .ZN(_01807_)
  );
  AND2_X1 _35998_ (
    .A1(_00008_[2]),
    .A2(_01807_),
    .ZN(_01808_)
  );
  AND2_X1 _35999_ (
    .A1(_01805_),
    .A2(_01808_),
    .ZN(_01809_)
  );
  INV_X1 _36000_ (
    .A(_01809_),
    .ZN(_01810_)
  );
  AND2_X1 _36001_ (
    .A1(_01803_),
    .A2(_01810_),
    .ZN(_01811_)
  );
  INV_X1 _36002_ (
    .A(_01811_),
    .ZN(_01812_)
  );
  AND2_X1 _36003_ (
    .A1(_22147_),
    .A2(_01812_),
    .ZN(_01813_)
  );
  INV_X1 _36004_ (
    .A(_01813_),
    .ZN(_01814_)
  );
  AND2_X1 _36005_ (
    .A1(_01796_),
    .A2(_01814_),
    .ZN(_01815_)
  );
  INV_X1 _36006_ (
    .A(_01815_),
    .ZN(_01816_)
  );
  AND2_X1 _36007_ (
    .A1(_22151_),
    .A2(_01816_),
    .ZN(_01817_)
  );
  INV_X1 _36008_ (
    .A(_01817_),
    .ZN(_01818_)
  );
  AND2_X1 _36009_ (
    .A1(_01778_),
    .A2(_01818_),
    .ZN(_01819_)
  );
  INV_X1 _36010_ (
    .A(_01819_),
    .ZN(_01820_)
  );
  AND2_X1 _36011_ (
    .A1(_00008_[3]),
    .A2(_01820_),
    .ZN(_01821_)
  );
  INV_X1 _36012_ (
    .A(_01821_),
    .ZN(_01822_)
  );
  AND2_X1 _36013_ (
    .A1(_22546_),
    .A2(_01738_),
    .ZN(_01823_)
  );
  AND2_X1 _36014_ (
    .A1(_01822_),
    .A2(_01823_),
    .ZN(_01824_)
  );
  INV_X1 _36015_ (
    .A(_01824_),
    .ZN(_01825_)
  );
  AND2_X1 _36016_ (
    .A1(_01658_),
    .A2(_01825_),
    .ZN(_01826_)
  );
  INV_X1 _36017_ (
    .A(_01826_),
    .ZN(_01827_)
  );
  AND2_X1 _36018_ (
    .A1(_22271_),
    .A2(_01827_),
    .ZN(_01828_)
  );
  INV_X1 _36019_ (
    .A(_01828_),
    .ZN(_01829_)
  );
  AND2_X1 _36020_ (
    .A1(reg_op1[26]),
    .A2(_22285_),
    .ZN(_01830_)
  );
  INV_X1 _36021_ (
    .A(_01830_),
    .ZN(_01831_)
  );
  AND2_X1 _36022_ (
    .A1(_27265_),
    .A2(_01831_),
    .ZN(_01832_)
  );
  AND2_X1 _36023_ (
    .A1(reg_op1[31]),
    .A2(_22290_),
    .ZN(_01833_)
  );
  INV_X1 _36024_ (
    .A(_01833_),
    .ZN(_01834_)
  );
  AND2_X1 _36025_ (
    .A1(_27262_),
    .A2(_01834_),
    .ZN(_01835_)
  );
  AND2_X1 _36026_ (
    .A1(_22573_),
    .A2(_01835_),
    .ZN(_01836_)
  );
  INV_X1 _36027_ (
    .A(_01836_),
    .ZN(_01837_)
  );
  AND2_X1 _36028_ (
    .A1(_22572_),
    .A2(_01832_),
    .ZN(_01838_)
  );
  INV_X1 _36029_ (
    .A(_01838_),
    .ZN(_01839_)
  );
  AND2_X1 _36030_ (
    .A1(_22295_),
    .A2(_01839_),
    .ZN(_01840_)
  );
  AND2_X1 _36031_ (
    .A1(_01837_),
    .A2(_01840_),
    .ZN(_01841_)
  );
  INV_X1 _36032_ (
    .A(_01841_),
    .ZN(_01842_)
  );
  AND2_X1 _36033_ (
    .A1(_22333_),
    .A2(_01842_),
    .ZN(_01843_)
  );
  AND2_X1 _36034_ (
    .A1(_01829_),
    .A2(_01843_),
    .ZN(_01844_)
  );
  AND2_X1 _36035_ (
    .A1(_01635_),
    .A2(_01647_),
    .ZN(_01845_)
  );
  INV_X1 _36036_ (
    .A(_01845_),
    .ZN(_01846_)
  );
  AND2_X1 _36037_ (
    .A1(reg_op1[27]),
    .A2(decoded_imm[27]),
    .ZN(_01847_)
  );
  INV_X1 _36038_ (
    .A(_01847_),
    .ZN(_01848_)
  );
  AND2_X1 _36039_ (
    .A1(_21194_),
    .A2(_21982_),
    .ZN(_01849_)
  );
  INV_X1 _36040_ (
    .A(_01849_),
    .ZN(_01850_)
  );
  AND2_X1 _36041_ (
    .A1(_01848_),
    .A2(_01850_),
    .ZN(_01851_)
  );
  INV_X1 _36042_ (
    .A(_01851_),
    .ZN(_01852_)
  );
  AND2_X1 _36043_ (
    .A1(_01846_),
    .A2(_01851_),
    .ZN(_01853_)
  );
  INV_X1 _36044_ (
    .A(_01853_),
    .ZN(_01854_)
  );
  AND2_X1 _36045_ (
    .A1(_01845_),
    .A2(_01852_),
    .ZN(_01855_)
  );
  INV_X1 _36046_ (
    .A(_01855_),
    .ZN(_01856_)
  );
  AND2_X1 _36047_ (
    .A1(_22559_),
    .A2(_01856_),
    .ZN(_01857_)
  );
  AND2_X1 _36048_ (
    .A1(_01854_),
    .A2(_01857_),
    .ZN(_01858_)
  );
  INV_X1 _36049_ (
    .A(_01858_),
    .ZN(_01859_)
  );
  AND2_X1 _36050_ (
    .A1(_01844_),
    .A2(_01859_),
    .ZN(_01860_)
  );
  INV_X1 _36051_ (
    .A(_01860_),
    .ZN(_01861_)
  );
  AND2_X1 _36052_ (
    .A1(_01656_),
    .A2(_01861_),
    .ZN(_00084_)
  );
  AND2_X1 _36053_ (
    .A1(_21195_),
    .A2(_22334_),
    .ZN(_01862_)
  );
  INV_X1 _36054_ (
    .A(_01862_),
    .ZN(_01863_)
  );
  AND2_X1 _36055_ (
    .A1(reg_pc[28]),
    .A2(_22335_),
    .ZN(_01864_)
  );
  INV_X1 _36056_ (
    .A(_01864_),
    .ZN(_01865_)
  );
  AND2_X1 _36057_ (
    .A1(_21801_),
    .A2(_00008_[2]),
    .ZN(_01866_)
  );
  INV_X1 _36058_ (
    .A(_01866_),
    .ZN(_01867_)
  );
  AND2_X1 _36059_ (
    .A1(_21509_),
    .A2(_22149_),
    .ZN(_01868_)
  );
  INV_X1 _36060_ (
    .A(_01868_),
    .ZN(_01869_)
  );
  AND2_X1 _36061_ (
    .A1(_00008_[0]),
    .A2(_01869_),
    .ZN(_01870_)
  );
  AND2_X1 _36062_ (
    .A1(_01867_),
    .A2(_01870_),
    .ZN(_01871_)
  );
  INV_X1 _36063_ (
    .A(_01871_),
    .ZN(_01872_)
  );
  AND2_X1 _36064_ (
    .A1(_21564_),
    .A2(_22149_),
    .ZN(_01873_)
  );
  INV_X1 _36065_ (
    .A(_01873_),
    .ZN(_01874_)
  );
  AND2_X1 _36066_ (
    .A1(_21830_),
    .A2(_00008_[2]),
    .ZN(_01875_)
  );
  INV_X1 _36067_ (
    .A(_01875_),
    .ZN(_01876_)
  );
  AND2_X1 _36068_ (
    .A1(_01874_),
    .A2(_01876_),
    .ZN(_01877_)
  );
  AND2_X1 _36069_ (
    .A1(_22147_),
    .A2(_01877_),
    .ZN(_01878_)
  );
  INV_X1 _36070_ (
    .A(_01878_),
    .ZN(_01879_)
  );
  AND2_X1 _36071_ (
    .A1(_01872_),
    .A2(_01879_),
    .ZN(_01880_)
  );
  AND2_X1 _36072_ (
    .A1(_21754_),
    .A2(_00008_[2]),
    .ZN(_01881_)
  );
  INV_X1 _36073_ (
    .A(_01881_),
    .ZN(_01882_)
  );
  AND2_X1 _36074_ (
    .A1(_21534_),
    .A2(_22149_),
    .ZN(_01883_)
  );
  INV_X1 _36075_ (
    .A(_01883_),
    .ZN(_01884_)
  );
  AND2_X1 _36076_ (
    .A1(_00008_[0]),
    .A2(_01882_),
    .ZN(_01885_)
  );
  AND2_X1 _36077_ (
    .A1(_01884_),
    .A2(_01885_),
    .ZN(_01886_)
  );
  INV_X1 _36078_ (
    .A(_01886_),
    .ZN(_01887_)
  );
  AND2_X1 _36079_ (
    .A1(_21975_),
    .A2(_22149_),
    .ZN(_01888_)
  );
  INV_X1 _36080_ (
    .A(_01888_),
    .ZN(_01889_)
  );
  AND2_X1 _36081_ (
    .A1(_21691_),
    .A2(_00008_[2]),
    .ZN(_01890_)
  );
  INV_X1 _36082_ (
    .A(_01890_),
    .ZN(_01891_)
  );
  AND2_X1 _36083_ (
    .A1(_01889_),
    .A2(_01891_),
    .ZN(_01892_)
  );
  AND2_X1 _36084_ (
    .A1(_22147_),
    .A2(_01892_),
    .ZN(_01893_)
  );
  INV_X1 _36085_ (
    .A(_01893_),
    .ZN(_01894_)
  );
  AND2_X1 _36086_ (
    .A1(_01887_),
    .A2(_01894_),
    .ZN(_01895_)
  );
  AND2_X1 _36087_ (
    .A1(_00008_[1]),
    .A2(_01880_),
    .ZN(_01896_)
  );
  INV_X1 _36088_ (
    .A(_01896_),
    .ZN(_01897_)
  );
  AND2_X1 _36089_ (
    .A1(_22148_),
    .A2(_01895_),
    .ZN(_01898_)
  );
  INV_X1 _36090_ (
    .A(_01898_),
    .ZN(_01899_)
  );
  AND2_X1 _36091_ (
    .A1(_01897_),
    .A2(_01899_),
    .ZN(_01900_)
  );
  AND2_X1 _36092_ (
    .A1(_22150_),
    .A2(_01900_),
    .ZN(_01901_)
  );
  INV_X1 _36093_ (
    .A(_01901_),
    .ZN(_01902_)
  );
  AND2_X1 _36094_ (
    .A1(\cpuregs[13] [28]),
    .A2(_00008_[0]),
    .ZN(_01903_)
  );
  INV_X1 _36095_ (
    .A(_01903_),
    .ZN(_01904_)
  );
  AND2_X1 _36096_ (
    .A1(\cpuregs[12] [28]),
    .A2(_22147_),
    .ZN(_01905_)
  );
  INV_X1 _36097_ (
    .A(_01905_),
    .ZN(_01906_)
  );
  AND2_X1 _36098_ (
    .A1(_00008_[2]),
    .A2(_01906_),
    .ZN(_01907_)
  );
  AND2_X1 _36099_ (
    .A1(_01904_),
    .A2(_01907_),
    .ZN(_01908_)
  );
  INV_X1 _36100_ (
    .A(_01908_),
    .ZN(_01909_)
  );
  AND2_X1 _36101_ (
    .A1(\cpuregs[9] [28]),
    .A2(_00008_[0]),
    .ZN(_01910_)
  );
  INV_X1 _36102_ (
    .A(_01910_),
    .ZN(_01911_)
  );
  AND2_X1 _36103_ (
    .A1(\cpuregs[8] [28]),
    .A2(_22147_),
    .ZN(_01912_)
  );
  INV_X1 _36104_ (
    .A(_01912_),
    .ZN(_01913_)
  );
  AND2_X1 _36105_ (
    .A1(_22149_),
    .A2(_01913_),
    .ZN(_01914_)
  );
  AND2_X1 _36106_ (
    .A1(_01911_),
    .A2(_01914_),
    .ZN(_01915_)
  );
  INV_X1 _36107_ (
    .A(_01915_),
    .ZN(_01916_)
  );
  AND2_X1 _36108_ (
    .A1(_22148_),
    .A2(_01916_),
    .ZN(_01917_)
  );
  AND2_X1 _36109_ (
    .A1(_01909_),
    .A2(_01917_),
    .ZN(_01918_)
  );
  INV_X1 _36110_ (
    .A(_01918_),
    .ZN(_01919_)
  );
  AND2_X1 _36111_ (
    .A1(\cpuregs[15] [28]),
    .A2(_00008_[0]),
    .ZN(_01920_)
  );
  INV_X1 _36112_ (
    .A(_01920_),
    .ZN(_01921_)
  );
  AND2_X1 _36113_ (
    .A1(\cpuregs[14] [28]),
    .A2(_22147_),
    .ZN(_01922_)
  );
  INV_X1 _36114_ (
    .A(_01922_),
    .ZN(_01923_)
  );
  AND2_X1 _36115_ (
    .A1(_00008_[2]),
    .A2(_01923_),
    .ZN(_01924_)
  );
  AND2_X1 _36116_ (
    .A1(_01921_),
    .A2(_01924_),
    .ZN(_01925_)
  );
  INV_X1 _36117_ (
    .A(_01925_),
    .ZN(_01926_)
  );
  AND2_X1 _36118_ (
    .A1(\cpuregs[11] [28]),
    .A2(_00008_[0]),
    .ZN(_01927_)
  );
  INV_X1 _36119_ (
    .A(_01927_),
    .ZN(_01928_)
  );
  AND2_X1 _36120_ (
    .A1(\cpuregs[10] [28]),
    .A2(_22147_),
    .ZN(_01929_)
  );
  INV_X1 _36121_ (
    .A(_01929_),
    .ZN(_01930_)
  );
  AND2_X1 _36122_ (
    .A1(_22149_),
    .A2(_01930_),
    .ZN(_01931_)
  );
  AND2_X1 _36123_ (
    .A1(_01928_),
    .A2(_01931_),
    .ZN(_01932_)
  );
  INV_X1 _36124_ (
    .A(_01932_),
    .ZN(_01933_)
  );
  AND2_X1 _36125_ (
    .A1(_00008_[1]),
    .A2(_01933_),
    .ZN(_01934_)
  );
  AND2_X1 _36126_ (
    .A1(_01926_),
    .A2(_01934_),
    .ZN(_01935_)
  );
  INV_X1 _36127_ (
    .A(_01935_),
    .ZN(_01936_)
  );
  AND2_X1 _36128_ (
    .A1(_01919_),
    .A2(_01936_),
    .ZN(_01937_)
  );
  INV_X1 _36129_ (
    .A(_01937_),
    .ZN(_01938_)
  );
  AND2_X1 _36130_ (
    .A1(_00008_[3]),
    .A2(_01938_),
    .ZN(_01939_)
  );
  INV_X1 _36131_ (
    .A(_01939_),
    .ZN(_01940_)
  );
  AND2_X1 _36132_ (
    .A1(_22151_),
    .A2(_01902_),
    .ZN(_01941_)
  );
  AND2_X1 _36133_ (
    .A1(_01940_),
    .A2(_01941_),
    .ZN(_01942_)
  );
  INV_X1 _36134_ (
    .A(_01942_),
    .ZN(_01943_)
  );
  AND2_X1 _36135_ (
    .A1(_21391_),
    .A2(_00008_[2]),
    .ZN(_01944_)
  );
  INV_X1 _36136_ (
    .A(_01944_),
    .ZN(_01945_)
  );
  AND2_X1 _36137_ (
    .A1(_21637_),
    .A2(_22149_),
    .ZN(_01946_)
  );
  INV_X1 _36138_ (
    .A(_01946_),
    .ZN(_01947_)
  );
  AND2_X1 _36139_ (
    .A1(_00008_[0]),
    .A2(_01947_),
    .ZN(_01948_)
  );
  AND2_X1 _36140_ (
    .A1(_01945_),
    .A2(_01948_),
    .ZN(_01949_)
  );
  INV_X1 _36141_ (
    .A(_01949_),
    .ZN(_01950_)
  );
  AND2_X1 _36142_ (
    .A1(_21613_),
    .A2(_22149_),
    .ZN(_01951_)
  );
  INV_X1 _36143_ (
    .A(_01951_),
    .ZN(_01952_)
  );
  AND2_X1 _36144_ (
    .A1(_21433_),
    .A2(_00008_[2]),
    .ZN(_01953_)
  );
  INV_X1 _36145_ (
    .A(_01953_),
    .ZN(_01954_)
  );
  AND2_X1 _36146_ (
    .A1(_01952_),
    .A2(_01954_),
    .ZN(_01955_)
  );
  AND2_X1 _36147_ (
    .A1(_22147_),
    .A2(_01955_),
    .ZN(_01956_)
  );
  INV_X1 _36148_ (
    .A(_01956_),
    .ZN(_01957_)
  );
  AND2_X1 _36149_ (
    .A1(_01950_),
    .A2(_01957_),
    .ZN(_01958_)
  );
  AND2_X1 _36150_ (
    .A1(_00008_[1]),
    .A2(_01958_),
    .ZN(_01959_)
  );
  INV_X1 _36151_ (
    .A(_01959_),
    .ZN(_01960_)
  );
  AND2_X1 _36152_ (
    .A1(_21777_),
    .A2(_00008_[2]),
    .ZN(_01961_)
  );
  INV_X1 _36153_ (
    .A(_01961_),
    .ZN(_01962_)
  );
  AND2_X1 _36154_ (
    .A1(_21478_),
    .A2(_22149_),
    .ZN(_01963_)
  );
  INV_X1 _36155_ (
    .A(_01963_),
    .ZN(_01964_)
  );
  AND2_X1 _36156_ (
    .A1(_00008_[0]),
    .A2(_01964_),
    .ZN(_01965_)
  );
  AND2_X1 _36157_ (
    .A1(_01962_),
    .A2(_01965_),
    .ZN(_01966_)
  );
  INV_X1 _36158_ (
    .A(_01966_),
    .ZN(_01967_)
  );
  AND2_X1 _36159_ (
    .A1(_21456_),
    .A2(_22149_),
    .ZN(_01968_)
  );
  INV_X1 _36160_ (
    .A(_01968_),
    .ZN(_01969_)
  );
  AND2_X1 _36161_ (
    .A1(_21667_),
    .A2(_00008_[2]),
    .ZN(_01970_)
  );
  INV_X1 _36162_ (
    .A(_01970_),
    .ZN(_01971_)
  );
  AND2_X1 _36163_ (
    .A1(_01969_),
    .A2(_01971_),
    .ZN(_01972_)
  );
  AND2_X1 _36164_ (
    .A1(_22147_),
    .A2(_01972_),
    .ZN(_01973_)
  );
  INV_X1 _36165_ (
    .A(_01973_),
    .ZN(_01974_)
  );
  AND2_X1 _36166_ (
    .A1(_01967_),
    .A2(_01974_),
    .ZN(_01975_)
  );
  AND2_X1 _36167_ (
    .A1(_22148_),
    .A2(_01975_),
    .ZN(_01976_)
  );
  INV_X1 _36168_ (
    .A(_01976_),
    .ZN(_01977_)
  );
  AND2_X1 _36169_ (
    .A1(_01960_),
    .A2(_01977_),
    .ZN(_01978_)
  );
  AND2_X1 _36170_ (
    .A1(_21886_),
    .A2(_22149_),
    .ZN(_01979_)
  );
  INV_X1 _36171_ (
    .A(_01979_),
    .ZN(_01980_)
  );
  AND2_X1 _36172_ (
    .A1(_21863_),
    .A2(_00008_[2]),
    .ZN(_01981_)
  );
  INV_X1 _36173_ (
    .A(_01981_),
    .ZN(_01982_)
  );
  AND2_X1 _36174_ (
    .A1(_01980_),
    .A2(_01982_),
    .ZN(_01983_)
  );
  AND2_X1 _36175_ (
    .A1(_22147_),
    .A2(_01983_),
    .ZN(_01984_)
  );
  INV_X1 _36176_ (
    .A(_01984_),
    .ZN(_01985_)
  );
  AND2_X1 _36177_ (
    .A1(_21951_),
    .A2(_00008_[2]),
    .ZN(_01986_)
  );
  INV_X1 _36178_ (
    .A(_01986_),
    .ZN(_01987_)
  );
  AND2_X1 _36179_ (
    .A1(_21935_),
    .A2(_22149_),
    .ZN(_01988_)
  );
  INV_X1 _36180_ (
    .A(_01988_),
    .ZN(_01989_)
  );
  AND2_X1 _36181_ (
    .A1(_00008_[0]),
    .A2(_01989_),
    .ZN(_01990_)
  );
  AND2_X1 _36182_ (
    .A1(_01987_),
    .A2(_01990_),
    .ZN(_01991_)
  );
  INV_X1 _36183_ (
    .A(_01991_),
    .ZN(_01992_)
  );
  AND2_X1 _36184_ (
    .A1(_01985_),
    .A2(_01992_),
    .ZN(_01993_)
  );
  AND2_X1 _36185_ (
    .A1(_00008_[1]),
    .A2(_01993_),
    .ZN(_01994_)
  );
  INV_X1 _36186_ (
    .A(_01994_),
    .ZN(_01995_)
  );
  AND2_X1 _36187_ (
    .A1(_21903_),
    .A2(_00008_[2]),
    .ZN(_01996_)
  );
  INV_X1 _36188_ (
    .A(_01996_),
    .ZN(_01997_)
  );
  AND2_X1 _36189_ (
    .A1(_21847_),
    .A2(_22149_),
    .ZN(_01998_)
  );
  INV_X1 _36190_ (
    .A(_01998_),
    .ZN(_01999_)
  );
  AND2_X1 _36191_ (
    .A1(_00008_[0]),
    .A2(_01999_),
    .ZN(_02000_)
  );
  AND2_X1 _36192_ (
    .A1(_01997_),
    .A2(_02000_),
    .ZN(_02001_)
  );
  INV_X1 _36193_ (
    .A(_02001_),
    .ZN(_02002_)
  );
  AND2_X1 _36194_ (
    .A1(_21581_),
    .A2(_22149_),
    .ZN(_02003_)
  );
  INV_X1 _36195_ (
    .A(_02003_),
    .ZN(_02004_)
  );
  AND2_X1 _36196_ (
    .A1(_21919_),
    .A2(_00008_[2]),
    .ZN(_02005_)
  );
  INV_X1 _36197_ (
    .A(_02005_),
    .ZN(_02006_)
  );
  AND2_X1 _36198_ (
    .A1(_02004_),
    .A2(_02006_),
    .ZN(_02007_)
  );
  AND2_X1 _36199_ (
    .A1(_22147_),
    .A2(_02007_),
    .ZN(_02008_)
  );
  INV_X1 _36200_ (
    .A(_02008_),
    .ZN(_02009_)
  );
  AND2_X1 _36201_ (
    .A1(_02002_),
    .A2(_02009_),
    .ZN(_02010_)
  );
  AND2_X1 _36202_ (
    .A1(_22148_),
    .A2(_02010_),
    .ZN(_02011_)
  );
  INV_X1 _36203_ (
    .A(_02011_),
    .ZN(_02012_)
  );
  AND2_X1 _36204_ (
    .A1(_00008_[3]),
    .A2(_02012_),
    .ZN(_02013_)
  );
  AND2_X1 _36205_ (
    .A1(_01995_),
    .A2(_02013_),
    .ZN(_02014_)
  );
  INV_X1 _36206_ (
    .A(_02014_),
    .ZN(_02015_)
  );
  AND2_X1 _36207_ (
    .A1(_22150_),
    .A2(_01978_),
    .ZN(_02016_)
  );
  INV_X1 _36208_ (
    .A(_02016_),
    .ZN(_02017_)
  );
  AND2_X1 _36209_ (
    .A1(_00008_[4]),
    .A2(_02015_),
    .ZN(_02018_)
  );
  AND2_X1 _36210_ (
    .A1(_02017_),
    .A2(_02018_),
    .ZN(_02019_)
  );
  INV_X1 _36211_ (
    .A(_02019_),
    .ZN(_02020_)
  );
  AND2_X1 _36212_ (
    .A1(_22546_),
    .A2(_02020_),
    .ZN(_02021_)
  );
  AND2_X1 _36213_ (
    .A1(_01943_),
    .A2(_02021_),
    .ZN(_02022_)
  );
  INV_X1 _36214_ (
    .A(_02022_),
    .ZN(_02023_)
  );
  AND2_X1 _36215_ (
    .A1(_01865_),
    .A2(_02023_),
    .ZN(_02024_)
  );
  INV_X1 _36216_ (
    .A(_02024_),
    .ZN(_02025_)
  );
  AND2_X1 _36217_ (
    .A1(_22271_),
    .A2(_02025_),
    .ZN(_02026_)
  );
  INV_X1 _36218_ (
    .A(_02026_),
    .ZN(_02027_)
  );
  AND2_X1 _36219_ (
    .A1(reg_op1[27]),
    .A2(_22285_),
    .ZN(_02028_)
  );
  INV_X1 _36220_ (
    .A(_02028_),
    .ZN(_02029_)
  );
  AND2_X1 _36221_ (
    .A1(_27471_),
    .A2(_02029_),
    .ZN(_02030_)
  );
  AND2_X1 _36222_ (
    .A1(reg_op1[31]),
    .A2(_22288_),
    .ZN(_02031_)
  );
  INV_X1 _36223_ (
    .A(_02031_),
    .ZN(_02032_)
  );
  AND2_X1 _36224_ (
    .A1(_27468_),
    .A2(_02032_),
    .ZN(_02033_)
  );
  AND2_X1 _36225_ (
    .A1(_22572_),
    .A2(_02030_),
    .ZN(_02034_)
  );
  INV_X1 _36226_ (
    .A(_02034_),
    .ZN(_02035_)
  );
  AND2_X1 _36227_ (
    .A1(_22573_),
    .A2(_02033_),
    .ZN(_02036_)
  );
  INV_X1 _36228_ (
    .A(_02036_),
    .ZN(_02037_)
  );
  AND2_X1 _36229_ (
    .A1(_22295_),
    .A2(_02037_),
    .ZN(_02038_)
  );
  AND2_X1 _36230_ (
    .A1(_02035_),
    .A2(_02038_),
    .ZN(_02039_)
  );
  INV_X1 _36231_ (
    .A(_02039_),
    .ZN(_02040_)
  );
  AND2_X1 _36232_ (
    .A1(_22333_),
    .A2(_02040_),
    .ZN(_02041_)
  );
  AND2_X1 _36233_ (
    .A1(_02027_),
    .A2(_02041_),
    .ZN(_02042_)
  );
  AND2_X1 _36234_ (
    .A1(reg_op1[28]),
    .A2(decoded_imm[28]),
    .ZN(_02043_)
  );
  INV_X1 _36235_ (
    .A(_02043_),
    .ZN(_02044_)
  );
  AND2_X1 _36236_ (
    .A1(_21195_),
    .A2(_21981_),
    .ZN(_02045_)
  );
  INV_X1 _36237_ (
    .A(_02045_),
    .ZN(_02046_)
  );
  AND2_X1 _36238_ (
    .A1(_02044_),
    .A2(_02046_),
    .ZN(_02047_)
  );
  INV_X1 _36239_ (
    .A(_02047_),
    .ZN(_02048_)
  );
  AND2_X1 _36240_ (
    .A1(_01846_),
    .A2(_01850_),
    .ZN(_02049_)
  );
  INV_X1 _36241_ (
    .A(_02049_),
    .ZN(_02050_)
  );
  AND2_X1 _36242_ (
    .A1(_01845_),
    .A2(_01848_),
    .ZN(_02051_)
  );
  INV_X1 _36243_ (
    .A(_02051_),
    .ZN(_02052_)
  );
  AND2_X1 _36244_ (
    .A1(_01848_),
    .A2(_02050_),
    .ZN(_02053_)
  );
  AND2_X1 _36245_ (
    .A1(_01850_),
    .A2(_02052_),
    .ZN(_02054_)
  );
  AND2_X1 _36246_ (
    .A1(_02047_),
    .A2(_02054_),
    .ZN(_02055_)
  );
  INV_X1 _36247_ (
    .A(_02055_),
    .ZN(_02056_)
  );
  AND2_X1 _36248_ (
    .A1(_02048_),
    .A2(_02053_),
    .ZN(_02057_)
  );
  INV_X1 _36249_ (
    .A(_02057_),
    .ZN(_02058_)
  );
  AND2_X1 _36250_ (
    .A1(_22559_),
    .A2(_02058_),
    .ZN(_02059_)
  );
  AND2_X1 _36251_ (
    .A1(_02056_),
    .A2(_02059_),
    .ZN(_02060_)
  );
  INV_X1 _36252_ (
    .A(_02060_),
    .ZN(_02061_)
  );
  AND2_X1 _36253_ (
    .A1(_02042_),
    .A2(_02061_),
    .ZN(_02062_)
  );
  INV_X1 _36254_ (
    .A(_02062_),
    .ZN(_02063_)
  );
  AND2_X1 _36255_ (
    .A1(_01863_),
    .A2(_02063_),
    .ZN(_00085_)
  );
  AND2_X1 _36256_ (
    .A1(_21196_),
    .A2(_22334_),
    .ZN(_02064_)
  );
  INV_X1 _36257_ (
    .A(_02064_),
    .ZN(_02065_)
  );
  AND2_X1 _36258_ (
    .A1(reg_pc[29]),
    .A2(_22335_),
    .ZN(_02066_)
  );
  INV_X1 _36259_ (
    .A(_02066_),
    .ZN(_02067_)
  );
  AND2_X1 _36260_ (
    .A1(_21565_),
    .A2(_22149_),
    .ZN(_02068_)
  );
  INV_X1 _36261_ (
    .A(_02068_),
    .ZN(_02069_)
  );
  AND2_X1 _36262_ (
    .A1(_21831_),
    .A2(_00008_[2]),
    .ZN(_02070_)
  );
  INV_X1 _36263_ (
    .A(_02070_),
    .ZN(_02071_)
  );
  AND2_X1 _36264_ (
    .A1(_02069_),
    .A2(_02071_),
    .ZN(_02072_)
  );
  AND2_X1 _36265_ (
    .A1(_22147_),
    .A2(_02072_),
    .ZN(_02073_)
  );
  INV_X1 _36266_ (
    .A(_02073_),
    .ZN(_02074_)
  );
  AND2_X1 _36267_ (
    .A1(_21802_),
    .A2(_00008_[2]),
    .ZN(_02075_)
  );
  INV_X1 _36268_ (
    .A(_02075_),
    .ZN(_02076_)
  );
  AND2_X1 _36269_ (
    .A1(_21510_),
    .A2(_22149_),
    .ZN(_02077_)
  );
  INV_X1 _36270_ (
    .A(_02077_),
    .ZN(_02078_)
  );
  AND2_X1 _36271_ (
    .A1(_00008_[0]),
    .A2(_02078_),
    .ZN(_02079_)
  );
  AND2_X1 _36272_ (
    .A1(_02076_),
    .A2(_02079_),
    .ZN(_02080_)
  );
  INV_X1 _36273_ (
    .A(_02080_),
    .ZN(_02081_)
  );
  AND2_X1 _36274_ (
    .A1(_02074_),
    .A2(_02081_),
    .ZN(_02082_)
  );
  AND2_X1 _36275_ (
    .A1(_21755_),
    .A2(_00008_[2]),
    .ZN(_02083_)
  );
  INV_X1 _36276_ (
    .A(_02083_),
    .ZN(_02084_)
  );
  AND2_X1 _36277_ (
    .A1(_21535_),
    .A2(_22149_),
    .ZN(_02085_)
  );
  INV_X1 _36278_ (
    .A(_02085_),
    .ZN(_02086_)
  );
  AND2_X1 _36279_ (
    .A1(_00008_[0]),
    .A2(_02084_),
    .ZN(_02087_)
  );
  AND2_X1 _36280_ (
    .A1(_02086_),
    .A2(_02087_),
    .ZN(_02088_)
  );
  INV_X1 _36281_ (
    .A(_02088_),
    .ZN(_02089_)
  );
  AND2_X1 _36282_ (
    .A1(_21976_),
    .A2(_22149_),
    .ZN(_02090_)
  );
  INV_X1 _36283_ (
    .A(_02090_),
    .ZN(_02091_)
  );
  AND2_X1 _36284_ (
    .A1(_21692_),
    .A2(_00008_[2]),
    .ZN(_02092_)
  );
  INV_X1 _36285_ (
    .A(_02092_),
    .ZN(_02093_)
  );
  AND2_X1 _36286_ (
    .A1(_02091_),
    .A2(_02093_),
    .ZN(_02094_)
  );
  AND2_X1 _36287_ (
    .A1(_22147_),
    .A2(_02094_),
    .ZN(_02095_)
  );
  INV_X1 _36288_ (
    .A(_02095_),
    .ZN(_02096_)
  );
  AND2_X1 _36289_ (
    .A1(_02089_),
    .A2(_02096_),
    .ZN(_02097_)
  );
  AND2_X1 _36290_ (
    .A1(_00008_[1]),
    .A2(_02082_),
    .ZN(_02098_)
  );
  INV_X1 _36291_ (
    .A(_02098_),
    .ZN(_02099_)
  );
  AND2_X1 _36292_ (
    .A1(_22148_),
    .A2(_02097_),
    .ZN(_02100_)
  );
  INV_X1 _36293_ (
    .A(_02100_),
    .ZN(_02101_)
  );
  AND2_X1 _36294_ (
    .A1(_02099_),
    .A2(_02101_),
    .ZN(_02102_)
  );
  AND2_X1 _36295_ (
    .A1(_22151_),
    .A2(_02102_),
    .ZN(_02103_)
  );
  INV_X1 _36296_ (
    .A(_02103_),
    .ZN(_02104_)
  );
  AND2_X1 _36297_ (
    .A1(_21392_),
    .A2(_00008_[2]),
    .ZN(_02105_)
  );
  INV_X1 _36298_ (
    .A(_02105_),
    .ZN(_02106_)
  );
  AND2_X1 _36299_ (
    .A1(_21638_),
    .A2(_22149_),
    .ZN(_02107_)
  );
  INV_X1 _36300_ (
    .A(_02107_),
    .ZN(_02108_)
  );
  AND2_X1 _36301_ (
    .A1(_00008_[0]),
    .A2(_02108_),
    .ZN(_02109_)
  );
  AND2_X1 _36302_ (
    .A1(_02106_),
    .A2(_02109_),
    .ZN(_02110_)
  );
  INV_X1 _36303_ (
    .A(_02110_),
    .ZN(_02111_)
  );
  AND2_X1 _36304_ (
    .A1(_21614_),
    .A2(_22149_),
    .ZN(_02112_)
  );
  INV_X1 _36305_ (
    .A(_02112_),
    .ZN(_02113_)
  );
  AND2_X1 _36306_ (
    .A1(_21434_),
    .A2(_00008_[2]),
    .ZN(_02114_)
  );
  INV_X1 _36307_ (
    .A(_02114_),
    .ZN(_02115_)
  );
  AND2_X1 _36308_ (
    .A1(_02113_),
    .A2(_02115_),
    .ZN(_02116_)
  );
  AND2_X1 _36309_ (
    .A1(_22147_),
    .A2(_02116_),
    .ZN(_02117_)
  );
  INV_X1 _36310_ (
    .A(_02117_),
    .ZN(_02118_)
  );
  AND2_X1 _36311_ (
    .A1(_02111_),
    .A2(_02118_),
    .ZN(_02119_)
  );
  AND2_X1 _36312_ (
    .A1(_21778_),
    .A2(_00008_[2]),
    .ZN(_02120_)
  );
  INV_X1 _36313_ (
    .A(_02120_),
    .ZN(_02121_)
  );
  AND2_X1 _36314_ (
    .A1(_21479_),
    .A2(_22149_),
    .ZN(_02122_)
  );
  INV_X1 _36315_ (
    .A(_02122_),
    .ZN(_02123_)
  );
  AND2_X1 _36316_ (
    .A1(_00008_[0]),
    .A2(_02121_),
    .ZN(_02124_)
  );
  AND2_X1 _36317_ (
    .A1(_02123_),
    .A2(_02124_),
    .ZN(_02125_)
  );
  INV_X1 _36318_ (
    .A(_02125_),
    .ZN(_02126_)
  );
  AND2_X1 _36319_ (
    .A1(_21457_),
    .A2(_22149_),
    .ZN(_02127_)
  );
  INV_X1 _36320_ (
    .A(_02127_),
    .ZN(_02128_)
  );
  AND2_X1 _36321_ (
    .A1(_21668_),
    .A2(_00008_[2]),
    .ZN(_02129_)
  );
  INV_X1 _36322_ (
    .A(_02129_),
    .ZN(_02130_)
  );
  AND2_X1 _36323_ (
    .A1(_02128_),
    .A2(_02130_),
    .ZN(_02131_)
  );
  AND2_X1 _36324_ (
    .A1(_22147_),
    .A2(_02131_),
    .ZN(_02132_)
  );
  INV_X1 _36325_ (
    .A(_02132_),
    .ZN(_02133_)
  );
  AND2_X1 _36326_ (
    .A1(_02126_),
    .A2(_02133_),
    .ZN(_02134_)
  );
  AND2_X1 _36327_ (
    .A1(_22148_),
    .A2(_02134_),
    .ZN(_02135_)
  );
  INV_X1 _36328_ (
    .A(_02135_),
    .ZN(_02136_)
  );
  AND2_X1 _36329_ (
    .A1(_00008_[1]),
    .A2(_02119_),
    .ZN(_02137_)
  );
  INV_X1 _36330_ (
    .A(_02137_),
    .ZN(_02138_)
  );
  AND2_X1 _36331_ (
    .A1(_00008_[4]),
    .A2(_02136_),
    .ZN(_02139_)
  );
  AND2_X1 _36332_ (
    .A1(_02138_),
    .A2(_02139_),
    .ZN(_02140_)
  );
  INV_X1 _36333_ (
    .A(_02140_),
    .ZN(_02141_)
  );
  AND2_X1 _36334_ (
    .A1(_02104_),
    .A2(_02141_),
    .ZN(_02142_)
  );
  AND2_X1 _36335_ (
    .A1(_22150_),
    .A2(_02142_),
    .ZN(_02143_)
  );
  INV_X1 _36336_ (
    .A(_02143_),
    .ZN(_02144_)
  );
  AND2_X1 _36337_ (
    .A1(_21588_),
    .A2(_22149_),
    .ZN(_02145_)
  );
  INV_X1 _36338_ (
    .A(_02145_),
    .ZN(_02146_)
  );
  AND2_X1 _36339_ (
    .A1(_21406_),
    .A2(_00008_[2]),
    .ZN(_02147_)
  );
  INV_X1 _36340_ (
    .A(_02147_),
    .ZN(_02148_)
  );
  AND2_X1 _36341_ (
    .A1(_21715_),
    .A2(_22149_),
    .ZN(_02149_)
  );
  INV_X1 _36342_ (
    .A(_02149_),
    .ZN(_02150_)
  );
  AND2_X1 _36343_ (
    .A1(_21399_),
    .A2(_00008_[2]),
    .ZN(_02151_)
  );
  INV_X1 _36344_ (
    .A(_02151_),
    .ZN(_02152_)
  );
  AND2_X1 _36345_ (
    .A1(_02150_),
    .A2(_02152_),
    .ZN(_02153_)
  );
  AND2_X1 _36346_ (
    .A1(_22147_),
    .A2(_02153_),
    .ZN(_02154_)
  );
  INV_X1 _36347_ (
    .A(_02154_),
    .ZN(_02155_)
  );
  AND2_X1 _36348_ (
    .A1(_00008_[0]),
    .A2(_02146_),
    .ZN(_02156_)
  );
  AND2_X1 _36349_ (
    .A1(_02148_),
    .A2(_02156_),
    .ZN(_02157_)
  );
  INV_X1 _36350_ (
    .A(_02157_),
    .ZN(_02158_)
  );
  AND2_X1 _36351_ (
    .A1(_02155_),
    .A2(_02158_),
    .ZN(_02159_)
  );
  AND2_X1 _36352_ (
    .A1(_00008_[1]),
    .A2(_02159_),
    .ZN(_02160_)
  );
  INV_X1 _36353_ (
    .A(_02160_),
    .ZN(_02161_)
  );
  AND2_X1 _36354_ (
    .A1(_21723_),
    .A2(_22149_),
    .ZN(_02162_)
  );
  INV_X1 _36355_ (
    .A(_02162_),
    .ZN(_02163_)
  );
  AND2_X1 _36356_ (
    .A1(_21645_),
    .A2(_00008_[2]),
    .ZN(_02164_)
  );
  INV_X1 _36357_ (
    .A(_02164_),
    .ZN(_02165_)
  );
  AND2_X1 _36358_ (
    .A1(_21730_),
    .A2(_22149_),
    .ZN(_02166_)
  );
  INV_X1 _36359_ (
    .A(_02166_),
    .ZN(_02167_)
  );
  AND2_X1 _36360_ (
    .A1(_21485_),
    .A2(_00008_[2]),
    .ZN(_02168_)
  );
  INV_X1 _36361_ (
    .A(_02168_),
    .ZN(_02169_)
  );
  AND2_X1 _36362_ (
    .A1(_02167_),
    .A2(_02169_),
    .ZN(_02170_)
  );
  AND2_X1 _36363_ (
    .A1(_00008_[0]),
    .A2(_02163_),
    .ZN(_02171_)
  );
  AND2_X1 _36364_ (
    .A1(_02165_),
    .A2(_02171_),
    .ZN(_02172_)
  );
  INV_X1 _36365_ (
    .A(_02172_),
    .ZN(_02173_)
  );
  AND2_X1 _36366_ (
    .A1(_22147_),
    .A2(_02170_),
    .ZN(_02174_)
  );
  INV_X1 _36367_ (
    .A(_02174_),
    .ZN(_02175_)
  );
  AND2_X1 _36368_ (
    .A1(_02173_),
    .A2(_02175_),
    .ZN(_02176_)
  );
  AND2_X1 _36369_ (
    .A1(_22148_),
    .A2(_02176_),
    .ZN(_02177_)
  );
  INV_X1 _36370_ (
    .A(_02177_),
    .ZN(_02178_)
  );
  AND2_X1 _36371_ (
    .A1(_22151_),
    .A2(_02178_),
    .ZN(_02179_)
  );
  AND2_X1 _36372_ (
    .A1(_02161_),
    .A2(_02179_),
    .ZN(_02180_)
  );
  INV_X1 _36373_ (
    .A(_02180_),
    .ZN(_02181_)
  );
  AND2_X1 _36374_ (
    .A1(_21904_),
    .A2(_00008_[2]),
    .ZN(_02182_)
  );
  INV_X1 _36375_ (
    .A(_02182_),
    .ZN(_02183_)
  );
  AND2_X1 _36376_ (
    .A1(_21848_),
    .A2(_22149_),
    .ZN(_02184_)
  );
  INV_X1 _36377_ (
    .A(_02184_),
    .ZN(_02185_)
  );
  AND2_X1 _36378_ (
    .A1(_00008_[0]),
    .A2(_02185_),
    .ZN(_02186_)
  );
  AND2_X1 _36379_ (
    .A1(_02183_),
    .A2(_02186_),
    .ZN(_02187_)
  );
  INV_X1 _36380_ (
    .A(_02187_),
    .ZN(_02188_)
  );
  AND2_X1 _36381_ (
    .A1(_21582_),
    .A2(_22149_),
    .ZN(_02189_)
  );
  INV_X1 _36382_ (
    .A(_02189_),
    .ZN(_02190_)
  );
  AND2_X1 _36383_ (
    .A1(_21920_),
    .A2(_00008_[2]),
    .ZN(_02191_)
  );
  INV_X1 _36384_ (
    .A(_02191_),
    .ZN(_02192_)
  );
  AND2_X1 _36385_ (
    .A1(_02190_),
    .A2(_02192_),
    .ZN(_02193_)
  );
  AND2_X1 _36386_ (
    .A1(_22147_),
    .A2(_02193_),
    .ZN(_02194_)
  );
  INV_X1 _36387_ (
    .A(_02194_),
    .ZN(_02195_)
  );
  AND2_X1 _36388_ (
    .A1(_02188_),
    .A2(_02195_),
    .ZN(_02196_)
  );
  AND2_X1 _36389_ (
    .A1(_22148_),
    .A2(_02196_),
    .ZN(_02197_)
  );
  INV_X1 _36390_ (
    .A(_02197_),
    .ZN(_02198_)
  );
  AND2_X1 _36391_ (
    .A1(_21887_),
    .A2(_22149_),
    .ZN(_02199_)
  );
  INV_X1 _36392_ (
    .A(_02199_),
    .ZN(_02200_)
  );
  AND2_X1 _36393_ (
    .A1(_21864_),
    .A2(_00008_[2]),
    .ZN(_02201_)
  );
  INV_X1 _36394_ (
    .A(_02201_),
    .ZN(_02202_)
  );
  AND2_X1 _36395_ (
    .A1(_02200_),
    .A2(_02202_),
    .ZN(_02203_)
  );
  AND2_X1 _36396_ (
    .A1(_22147_),
    .A2(_02203_),
    .ZN(_02204_)
  );
  INV_X1 _36397_ (
    .A(_02204_),
    .ZN(_02205_)
  );
  AND2_X1 _36398_ (
    .A1(_21952_),
    .A2(_00008_[2]),
    .ZN(_02206_)
  );
  INV_X1 _36399_ (
    .A(_02206_),
    .ZN(_02207_)
  );
  AND2_X1 _36400_ (
    .A1(_21936_),
    .A2(_22149_),
    .ZN(_02208_)
  );
  INV_X1 _36401_ (
    .A(_02208_),
    .ZN(_02209_)
  );
  AND2_X1 _36402_ (
    .A1(_00008_[0]),
    .A2(_02209_),
    .ZN(_02210_)
  );
  AND2_X1 _36403_ (
    .A1(_02207_),
    .A2(_02210_),
    .ZN(_02211_)
  );
  INV_X1 _36404_ (
    .A(_02211_),
    .ZN(_02212_)
  );
  AND2_X1 _36405_ (
    .A1(_02205_),
    .A2(_02212_),
    .ZN(_02213_)
  );
  AND2_X1 _36406_ (
    .A1(_00008_[1]),
    .A2(_02213_),
    .ZN(_02214_)
  );
  INV_X1 _36407_ (
    .A(_02214_),
    .ZN(_02215_)
  );
  AND2_X1 _36408_ (
    .A1(_00008_[4]),
    .A2(_02215_),
    .ZN(_02216_)
  );
  AND2_X1 _36409_ (
    .A1(_02198_),
    .A2(_02216_),
    .ZN(_02217_)
  );
  INV_X1 _36410_ (
    .A(_02217_),
    .ZN(_02218_)
  );
  AND2_X1 _36411_ (
    .A1(_02181_),
    .A2(_02218_),
    .ZN(_02219_)
  );
  AND2_X1 _36412_ (
    .A1(_00008_[3]),
    .A2(_02219_),
    .ZN(_02220_)
  );
  INV_X1 _36413_ (
    .A(_02220_),
    .ZN(_02221_)
  );
  AND2_X1 _36414_ (
    .A1(_22546_),
    .A2(_02221_),
    .ZN(_02222_)
  );
  AND2_X1 _36415_ (
    .A1(_02144_),
    .A2(_02222_),
    .ZN(_02223_)
  );
  INV_X1 _36416_ (
    .A(_02223_),
    .ZN(_02224_)
  );
  AND2_X1 _36417_ (
    .A1(_02067_),
    .A2(_02224_),
    .ZN(_02225_)
  );
  INV_X1 _36418_ (
    .A(_02225_),
    .ZN(_02226_)
  );
  AND2_X1 _36419_ (
    .A1(_22271_),
    .A2(_02226_),
    .ZN(_02227_)
  );
  INV_X1 _36420_ (
    .A(_02227_),
    .ZN(_02228_)
  );
  AND2_X1 _36421_ (
    .A1(reg_op1[28]),
    .A2(_22285_),
    .ZN(_02229_)
  );
  INV_X1 _36422_ (
    .A(_02229_),
    .ZN(_02230_)
  );
  AND2_X1 _36423_ (
    .A1(_01623_),
    .A2(_02230_),
    .ZN(_02231_)
  );
  AND2_X1 _36424_ (
    .A1(_01620_),
    .A2(_02032_),
    .ZN(_02232_)
  );
  AND2_X1 _36425_ (
    .A1(_22572_),
    .A2(_02231_),
    .ZN(_02233_)
  );
  INV_X1 _36426_ (
    .A(_02233_),
    .ZN(_02234_)
  );
  AND2_X1 _36427_ (
    .A1(_22573_),
    .A2(_02232_),
    .ZN(_02235_)
  );
  INV_X1 _36428_ (
    .A(_02235_),
    .ZN(_02236_)
  );
  AND2_X1 _36429_ (
    .A1(_22295_),
    .A2(_02236_),
    .ZN(_02237_)
  );
  AND2_X1 _36430_ (
    .A1(_02234_),
    .A2(_02237_),
    .ZN(_02238_)
  );
  INV_X1 _36431_ (
    .A(_02238_),
    .ZN(_02239_)
  );
  AND2_X1 _36432_ (
    .A1(_22333_),
    .A2(_02228_),
    .ZN(_02240_)
  );
  AND2_X1 _36433_ (
    .A1(_02239_),
    .A2(_02240_),
    .ZN(_02241_)
  );
  AND2_X1 _36434_ (
    .A1(_02044_),
    .A2(_02056_),
    .ZN(_02242_)
  );
  INV_X1 _36435_ (
    .A(_02242_),
    .ZN(_02243_)
  );
  AND2_X1 _36436_ (
    .A1(reg_op1[29]),
    .A2(decoded_imm[29]),
    .ZN(_02244_)
  );
  INV_X1 _36437_ (
    .A(_02244_),
    .ZN(_02245_)
  );
  AND2_X1 _36438_ (
    .A1(_21196_),
    .A2(_21980_),
    .ZN(_02246_)
  );
  INV_X1 _36439_ (
    .A(_02246_),
    .ZN(_02247_)
  );
  AND2_X1 _36440_ (
    .A1(_02245_),
    .A2(_02247_),
    .ZN(_02248_)
  );
  INV_X1 _36441_ (
    .A(_02248_),
    .ZN(_02249_)
  );
  AND2_X1 _36442_ (
    .A1(_02243_),
    .A2(_02248_),
    .ZN(_02250_)
  );
  INV_X1 _36443_ (
    .A(_02250_),
    .ZN(_02251_)
  );
  AND2_X1 _36444_ (
    .A1(_02242_),
    .A2(_02249_),
    .ZN(_02252_)
  );
  INV_X1 _36445_ (
    .A(_02252_),
    .ZN(_02253_)
  );
  AND2_X1 _36446_ (
    .A1(_22559_),
    .A2(_02253_),
    .ZN(_02254_)
  );
  AND2_X1 _36447_ (
    .A1(_02251_),
    .A2(_02254_),
    .ZN(_02255_)
  );
  INV_X1 _36448_ (
    .A(_02255_),
    .ZN(_02256_)
  );
  AND2_X1 _36449_ (
    .A1(_02241_),
    .A2(_02256_),
    .ZN(_02257_)
  );
  INV_X1 _36450_ (
    .A(_02257_),
    .ZN(_02258_)
  );
  AND2_X1 _36451_ (
    .A1(_02065_),
    .A2(_02258_),
    .ZN(_00086_)
  );
  AND2_X1 _36452_ (
    .A1(_21197_),
    .A2(_22334_),
    .ZN(_02259_)
  );
  INV_X1 _36453_ (
    .A(_02259_),
    .ZN(_02260_)
  );
  AND2_X1 _36454_ (
    .A1(reg_pc[30]),
    .A2(_22335_),
    .ZN(_02261_)
  );
  INV_X1 _36455_ (
    .A(_02261_),
    .ZN(_02262_)
  );
  AND2_X1 _36456_ (
    .A1(_21566_),
    .A2(_22149_),
    .ZN(_02263_)
  );
  INV_X1 _36457_ (
    .A(_02263_),
    .ZN(_02264_)
  );
  AND2_X1 _36458_ (
    .A1(_21832_),
    .A2(_00008_[2]),
    .ZN(_02265_)
  );
  INV_X1 _36459_ (
    .A(_02265_),
    .ZN(_02266_)
  );
  AND2_X1 _36460_ (
    .A1(_02264_),
    .A2(_02266_),
    .ZN(_02267_)
  );
  AND2_X1 _36461_ (
    .A1(_22147_),
    .A2(_02267_),
    .ZN(_02268_)
  );
  INV_X1 _36462_ (
    .A(_02268_),
    .ZN(_02269_)
  );
  AND2_X1 _36463_ (
    .A1(_21803_),
    .A2(_00008_[2]),
    .ZN(_02270_)
  );
  INV_X1 _36464_ (
    .A(_02270_),
    .ZN(_02271_)
  );
  AND2_X1 _36465_ (
    .A1(_21511_),
    .A2(_22149_),
    .ZN(_02272_)
  );
  INV_X1 _36466_ (
    .A(_02272_),
    .ZN(_02273_)
  );
  AND2_X1 _36467_ (
    .A1(_00008_[0]),
    .A2(_02273_),
    .ZN(_02274_)
  );
  AND2_X1 _36468_ (
    .A1(_02271_),
    .A2(_02274_),
    .ZN(_02275_)
  );
  INV_X1 _36469_ (
    .A(_02275_),
    .ZN(_02276_)
  );
  AND2_X1 _36470_ (
    .A1(_02269_),
    .A2(_02276_),
    .ZN(_02277_)
  );
  AND2_X1 _36471_ (
    .A1(_21756_),
    .A2(_00008_[2]),
    .ZN(_02278_)
  );
  INV_X1 _36472_ (
    .A(_02278_),
    .ZN(_02279_)
  );
  AND2_X1 _36473_ (
    .A1(_21536_),
    .A2(_22149_),
    .ZN(_02280_)
  );
  INV_X1 _36474_ (
    .A(_02280_),
    .ZN(_02281_)
  );
  AND2_X1 _36475_ (
    .A1(_00008_[0]),
    .A2(_02279_),
    .ZN(_02282_)
  );
  AND2_X1 _36476_ (
    .A1(_02281_),
    .A2(_02282_),
    .ZN(_02283_)
  );
  INV_X1 _36477_ (
    .A(_02283_),
    .ZN(_02284_)
  );
  AND2_X1 _36478_ (
    .A1(_21977_),
    .A2(_22149_),
    .ZN(_02285_)
  );
  INV_X1 _36479_ (
    .A(_02285_),
    .ZN(_02286_)
  );
  AND2_X1 _36480_ (
    .A1(_21693_),
    .A2(_00008_[2]),
    .ZN(_02287_)
  );
  INV_X1 _36481_ (
    .A(_02287_),
    .ZN(_02288_)
  );
  AND2_X1 _36482_ (
    .A1(_02286_),
    .A2(_02288_),
    .ZN(_02289_)
  );
  AND2_X1 _36483_ (
    .A1(_22147_),
    .A2(_02289_),
    .ZN(_02290_)
  );
  INV_X1 _36484_ (
    .A(_02290_),
    .ZN(_02291_)
  );
  AND2_X1 _36485_ (
    .A1(_02284_),
    .A2(_02291_),
    .ZN(_02292_)
  );
  AND2_X1 _36486_ (
    .A1(_00008_[1]),
    .A2(_02277_),
    .ZN(_02293_)
  );
  INV_X1 _36487_ (
    .A(_02293_),
    .ZN(_02294_)
  );
  AND2_X1 _36488_ (
    .A1(_22148_),
    .A2(_02292_),
    .ZN(_02295_)
  );
  INV_X1 _36489_ (
    .A(_02295_),
    .ZN(_02296_)
  );
  AND2_X1 _36490_ (
    .A1(_02294_),
    .A2(_02296_),
    .ZN(_02297_)
  );
  AND2_X1 _36491_ (
    .A1(_22151_),
    .A2(_02297_),
    .ZN(_02298_)
  );
  INV_X1 _36492_ (
    .A(_02298_),
    .ZN(_02299_)
  );
  AND2_X1 _36493_ (
    .A1(\cpuregs[23] [30]),
    .A2(_00008_[2]),
    .ZN(_02300_)
  );
  INV_X1 _36494_ (
    .A(_02300_),
    .ZN(_02301_)
  );
  AND2_X1 _36495_ (
    .A1(\cpuregs[19] [30]),
    .A2(_22149_),
    .ZN(_02302_)
  );
  INV_X1 _36496_ (
    .A(_02302_),
    .ZN(_02303_)
  );
  AND2_X1 _36497_ (
    .A1(_02301_),
    .A2(_02303_),
    .ZN(_02304_)
  );
  INV_X1 _36498_ (
    .A(_02304_),
    .ZN(_02305_)
  );
  AND2_X1 _36499_ (
    .A1(_00008_[0]),
    .A2(_02305_),
    .ZN(_02306_)
  );
  INV_X1 _36500_ (
    .A(_02306_),
    .ZN(_02307_)
  );
  AND2_X1 _36501_ (
    .A1(_21615_),
    .A2(_22149_),
    .ZN(_02308_)
  );
  INV_X1 _36502_ (
    .A(_02308_),
    .ZN(_02309_)
  );
  AND2_X1 _36503_ (
    .A1(_21435_),
    .A2(_00008_[2]),
    .ZN(_02310_)
  );
  INV_X1 _36504_ (
    .A(_02310_),
    .ZN(_02311_)
  );
  AND2_X1 _36505_ (
    .A1(_02309_),
    .A2(_02311_),
    .ZN(_02312_)
  );
  AND2_X1 _36506_ (
    .A1(_22147_),
    .A2(_02312_),
    .ZN(_02313_)
  );
  INV_X1 _36507_ (
    .A(_02313_),
    .ZN(_02314_)
  );
  AND2_X1 _36508_ (
    .A1(\cpuregs[21] [30]),
    .A2(_00008_[2]),
    .ZN(_02315_)
  );
  INV_X1 _36509_ (
    .A(_02315_),
    .ZN(_02316_)
  );
  AND2_X1 _36510_ (
    .A1(\cpuregs[17] [30]),
    .A2(_22149_),
    .ZN(_02317_)
  );
  INV_X1 _36511_ (
    .A(_02317_),
    .ZN(_02318_)
  );
  AND2_X1 _36512_ (
    .A1(_02316_),
    .A2(_02318_),
    .ZN(_02319_)
  );
  INV_X1 _36513_ (
    .A(_02319_),
    .ZN(_02320_)
  );
  AND2_X1 _36514_ (
    .A1(_00008_[0]),
    .A2(_02320_),
    .ZN(_02321_)
  );
  INV_X1 _36515_ (
    .A(_02321_),
    .ZN(_02322_)
  );
  AND2_X1 _36516_ (
    .A1(\cpuregs[20] [30]),
    .A2(_00008_[2]),
    .ZN(_02323_)
  );
  INV_X1 _36517_ (
    .A(_02323_),
    .ZN(_02324_)
  );
  AND2_X1 _36518_ (
    .A1(\cpuregs[16] [30]),
    .A2(_22149_),
    .ZN(_02325_)
  );
  INV_X1 _36519_ (
    .A(_02325_),
    .ZN(_02326_)
  );
  AND2_X1 _36520_ (
    .A1(_02324_),
    .A2(_02326_),
    .ZN(_02327_)
  );
  INV_X1 _36521_ (
    .A(_02327_),
    .ZN(_02328_)
  );
  AND2_X1 _36522_ (
    .A1(_22147_),
    .A2(_02328_),
    .ZN(_02329_)
  );
  INV_X1 _36523_ (
    .A(_02329_),
    .ZN(_02330_)
  );
  AND2_X1 _36524_ (
    .A1(_02322_),
    .A2(_02330_),
    .ZN(_02331_)
  );
  AND2_X1 _36525_ (
    .A1(_22148_),
    .A2(_02331_),
    .ZN(_02332_)
  );
  INV_X1 _36526_ (
    .A(_02332_),
    .ZN(_02333_)
  );
  AND2_X1 _36527_ (
    .A1(_00008_[1]),
    .A2(_02314_),
    .ZN(_02334_)
  );
  AND2_X1 _36528_ (
    .A1(_02307_),
    .A2(_02334_),
    .ZN(_02335_)
  );
  INV_X1 _36529_ (
    .A(_02335_),
    .ZN(_02336_)
  );
  AND2_X1 _36530_ (
    .A1(_00008_[4]),
    .A2(_02333_),
    .ZN(_02337_)
  );
  AND2_X1 _36531_ (
    .A1(_02336_),
    .A2(_02337_),
    .ZN(_02338_)
  );
  INV_X1 _36532_ (
    .A(_02338_),
    .ZN(_02339_)
  );
  AND2_X1 _36533_ (
    .A1(_22150_),
    .A2(_02299_),
    .ZN(_02340_)
  );
  AND2_X1 _36534_ (
    .A1(_02339_),
    .A2(_02340_),
    .ZN(_02341_)
  );
  INV_X1 _36535_ (
    .A(_02341_),
    .ZN(_02342_)
  );
  AND2_X1 _36536_ (
    .A1(_21589_),
    .A2(_22149_),
    .ZN(_02343_)
  );
  INV_X1 _36537_ (
    .A(_02343_),
    .ZN(_02344_)
  );
  AND2_X1 _36538_ (
    .A1(_21407_),
    .A2(_00008_[2]),
    .ZN(_02345_)
  );
  INV_X1 _36539_ (
    .A(_02345_),
    .ZN(_02346_)
  );
  AND2_X1 _36540_ (
    .A1(_21716_),
    .A2(_22149_),
    .ZN(_02347_)
  );
  INV_X1 _36541_ (
    .A(_02347_),
    .ZN(_02348_)
  );
  AND2_X1 _36542_ (
    .A1(_21400_),
    .A2(_00008_[2]),
    .ZN(_02349_)
  );
  INV_X1 _36543_ (
    .A(_02349_),
    .ZN(_02350_)
  );
  AND2_X1 _36544_ (
    .A1(_02348_),
    .A2(_02350_),
    .ZN(_02351_)
  );
  AND2_X1 _36545_ (
    .A1(_22147_),
    .A2(_02351_),
    .ZN(_02352_)
  );
  INV_X1 _36546_ (
    .A(_02352_),
    .ZN(_02353_)
  );
  AND2_X1 _36547_ (
    .A1(_00008_[0]),
    .A2(_02344_),
    .ZN(_02354_)
  );
  AND2_X1 _36548_ (
    .A1(_02346_),
    .A2(_02354_),
    .ZN(_02355_)
  );
  INV_X1 _36549_ (
    .A(_02355_),
    .ZN(_02356_)
  );
  AND2_X1 _36550_ (
    .A1(_02353_),
    .A2(_02356_),
    .ZN(_02357_)
  );
  AND2_X1 _36551_ (
    .A1(_00008_[1]),
    .A2(_02357_),
    .ZN(_02358_)
  );
  INV_X1 _36552_ (
    .A(_02358_),
    .ZN(_02359_)
  );
  AND2_X1 _36553_ (
    .A1(_21724_),
    .A2(_22149_),
    .ZN(_02360_)
  );
  INV_X1 _36554_ (
    .A(_02360_),
    .ZN(_02361_)
  );
  AND2_X1 _36555_ (
    .A1(_21646_),
    .A2(_00008_[2]),
    .ZN(_02362_)
  );
  INV_X1 _36556_ (
    .A(_02362_),
    .ZN(_02363_)
  );
  AND2_X1 _36557_ (
    .A1(_21731_),
    .A2(_22149_),
    .ZN(_02364_)
  );
  INV_X1 _36558_ (
    .A(_02364_),
    .ZN(_02365_)
  );
  AND2_X1 _36559_ (
    .A1(_21486_),
    .A2(_00008_[2]),
    .ZN(_02366_)
  );
  INV_X1 _36560_ (
    .A(_02366_),
    .ZN(_02367_)
  );
  AND2_X1 _36561_ (
    .A1(_02365_),
    .A2(_02367_),
    .ZN(_02368_)
  );
  AND2_X1 _36562_ (
    .A1(_00008_[0]),
    .A2(_02361_),
    .ZN(_02369_)
  );
  AND2_X1 _36563_ (
    .A1(_02363_),
    .A2(_02369_),
    .ZN(_02370_)
  );
  INV_X1 _36564_ (
    .A(_02370_),
    .ZN(_02371_)
  );
  AND2_X1 _36565_ (
    .A1(_22147_),
    .A2(_02368_),
    .ZN(_02372_)
  );
  INV_X1 _36566_ (
    .A(_02372_),
    .ZN(_02373_)
  );
  AND2_X1 _36567_ (
    .A1(_02371_),
    .A2(_02373_),
    .ZN(_02374_)
  );
  AND2_X1 _36568_ (
    .A1(_22148_),
    .A2(_02374_),
    .ZN(_02375_)
  );
  INV_X1 _36569_ (
    .A(_02375_),
    .ZN(_02376_)
  );
  AND2_X1 _36570_ (
    .A1(_02359_),
    .A2(_02376_),
    .ZN(_02377_)
  );
  INV_X1 _36571_ (
    .A(_02377_),
    .ZN(_02378_)
  );
  AND2_X1 _36572_ (
    .A1(_22151_),
    .A2(_02378_),
    .ZN(_02379_)
  );
  INV_X1 _36573_ (
    .A(_02379_),
    .ZN(_02380_)
  );
  AND2_X1 _36574_ (
    .A1(\cpuregs[25] [30]),
    .A2(_22148_),
    .ZN(_02381_)
  );
  INV_X1 _36575_ (
    .A(_02381_),
    .ZN(_02382_)
  );
  AND2_X1 _36576_ (
    .A1(\cpuregs[27] [30]),
    .A2(_00008_[1]),
    .ZN(_02383_)
  );
  INV_X1 _36577_ (
    .A(_02383_),
    .ZN(_02384_)
  );
  AND2_X1 _36578_ (
    .A1(_22149_),
    .A2(_02384_),
    .ZN(_02385_)
  );
  AND2_X1 _36579_ (
    .A1(_02382_),
    .A2(_02385_),
    .ZN(_02386_)
  );
  INV_X1 _36580_ (
    .A(_02386_),
    .ZN(_02387_)
  );
  AND2_X1 _36581_ (
    .A1(\cpuregs[29] [30]),
    .A2(_22148_),
    .ZN(_02388_)
  );
  INV_X1 _36582_ (
    .A(_02388_),
    .ZN(_02389_)
  );
  AND2_X1 _36583_ (
    .A1(\cpuregs[31] [30]),
    .A2(_00008_[1]),
    .ZN(_02390_)
  );
  INV_X1 _36584_ (
    .A(_02390_),
    .ZN(_02391_)
  );
  AND2_X1 _36585_ (
    .A1(_00008_[2]),
    .A2(_02391_),
    .ZN(_02392_)
  );
  AND2_X1 _36586_ (
    .A1(_02389_),
    .A2(_02392_),
    .ZN(_02393_)
  );
  INV_X1 _36587_ (
    .A(_02393_),
    .ZN(_02394_)
  );
  AND2_X1 _36588_ (
    .A1(_02387_),
    .A2(_02394_),
    .ZN(_02395_)
  );
  INV_X1 _36589_ (
    .A(_02395_),
    .ZN(_02396_)
  );
  AND2_X1 _36590_ (
    .A1(_00008_[0]),
    .A2(_02396_),
    .ZN(_02397_)
  );
  INV_X1 _36591_ (
    .A(_02397_),
    .ZN(_02398_)
  );
  AND2_X1 _36592_ (
    .A1(\cpuregs[24] [30]),
    .A2(_22148_),
    .ZN(_02399_)
  );
  INV_X1 _36593_ (
    .A(_02399_),
    .ZN(_02400_)
  );
  AND2_X1 _36594_ (
    .A1(\cpuregs[26] [30]),
    .A2(_00008_[1]),
    .ZN(_02401_)
  );
  INV_X1 _36595_ (
    .A(_02401_),
    .ZN(_02402_)
  );
  AND2_X1 _36596_ (
    .A1(_22149_),
    .A2(_02402_),
    .ZN(_02403_)
  );
  AND2_X1 _36597_ (
    .A1(_02400_),
    .A2(_02403_),
    .ZN(_02404_)
  );
  INV_X1 _36598_ (
    .A(_02404_),
    .ZN(_02405_)
  );
  AND2_X1 _36599_ (
    .A1(\cpuregs[28] [30]),
    .A2(_22148_),
    .ZN(_02406_)
  );
  INV_X1 _36600_ (
    .A(_02406_),
    .ZN(_02407_)
  );
  AND2_X1 _36601_ (
    .A1(\cpuregs[30] [30]),
    .A2(_00008_[1]),
    .ZN(_02408_)
  );
  INV_X1 _36602_ (
    .A(_02408_),
    .ZN(_02409_)
  );
  AND2_X1 _36603_ (
    .A1(_00008_[2]),
    .A2(_02409_),
    .ZN(_02410_)
  );
  AND2_X1 _36604_ (
    .A1(_02407_),
    .A2(_02410_),
    .ZN(_02411_)
  );
  INV_X1 _36605_ (
    .A(_02411_),
    .ZN(_02412_)
  );
  AND2_X1 _36606_ (
    .A1(_02405_),
    .A2(_02412_),
    .ZN(_02413_)
  );
  INV_X1 _36607_ (
    .A(_02413_),
    .ZN(_02414_)
  );
  AND2_X1 _36608_ (
    .A1(_22147_),
    .A2(_02414_),
    .ZN(_02415_)
  );
  INV_X1 _36609_ (
    .A(_02415_),
    .ZN(_02416_)
  );
  AND2_X1 _36610_ (
    .A1(_02398_),
    .A2(_02416_),
    .ZN(_02417_)
  );
  INV_X1 _36611_ (
    .A(_02417_),
    .ZN(_02418_)
  );
  AND2_X1 _36612_ (
    .A1(_00008_[4]),
    .A2(_02418_),
    .ZN(_02419_)
  );
  INV_X1 _36613_ (
    .A(_02419_),
    .ZN(_02420_)
  );
  AND2_X1 _36614_ (
    .A1(_02380_),
    .A2(_02420_),
    .ZN(_02421_)
  );
  INV_X1 _36615_ (
    .A(_02421_),
    .ZN(_02422_)
  );
  AND2_X1 _36616_ (
    .A1(_00008_[3]),
    .A2(_02422_),
    .ZN(_02423_)
  );
  INV_X1 _36617_ (
    .A(_02423_),
    .ZN(_02424_)
  );
  AND2_X1 _36618_ (
    .A1(_22546_),
    .A2(_02342_),
    .ZN(_02425_)
  );
  AND2_X1 _36619_ (
    .A1(_02424_),
    .A2(_02425_),
    .ZN(_02426_)
  );
  INV_X1 _36620_ (
    .A(_02426_),
    .ZN(_02427_)
  );
  AND2_X1 _36621_ (
    .A1(_02262_),
    .A2(_02427_),
    .ZN(_02428_)
  );
  INV_X1 _36622_ (
    .A(_02428_),
    .ZN(_02429_)
  );
  AND2_X1 _36623_ (
    .A1(_22271_),
    .A2(_02429_),
    .ZN(_02430_)
  );
  INV_X1 _36624_ (
    .A(_02430_),
    .ZN(_02431_)
  );
  AND2_X1 _36625_ (
    .A1(reg_op1[29]),
    .A2(_22285_),
    .ZN(_02432_)
  );
  INV_X1 _36626_ (
    .A(_02432_),
    .ZN(_02433_)
  );
  AND2_X1 _36627_ (
    .A1(_01834_),
    .A2(_02433_),
    .ZN(_02434_)
  );
  AND2_X1 _36628_ (
    .A1(_01831_),
    .A2(_02032_),
    .ZN(_02435_)
  );
  AND2_X1 _36629_ (
    .A1(_22572_),
    .A2(_02434_),
    .ZN(_02436_)
  );
  INV_X1 _36630_ (
    .A(_02436_),
    .ZN(_02437_)
  );
  AND2_X1 _36631_ (
    .A1(_22573_),
    .A2(_02435_),
    .ZN(_02438_)
  );
  INV_X1 _36632_ (
    .A(_02438_),
    .ZN(_02439_)
  );
  AND2_X1 _36633_ (
    .A1(_22295_),
    .A2(_02439_),
    .ZN(_02440_)
  );
  AND2_X1 _36634_ (
    .A1(_02437_),
    .A2(_02440_),
    .ZN(_02441_)
  );
  INV_X1 _36635_ (
    .A(_02441_),
    .ZN(_02442_)
  );
  AND2_X1 _36636_ (
    .A1(_22333_),
    .A2(_02431_),
    .ZN(_02443_)
  );
  AND2_X1 _36637_ (
    .A1(_02442_),
    .A2(_02443_),
    .ZN(_02444_)
  );
  AND2_X1 _36638_ (
    .A1(_02245_),
    .A2(_02251_),
    .ZN(_02445_)
  );
  INV_X1 _36639_ (
    .A(_02445_),
    .ZN(_02446_)
  );
  AND2_X1 _36640_ (
    .A1(reg_op1[30]),
    .A2(decoded_imm[30]),
    .ZN(_02447_)
  );
  INV_X1 _36641_ (
    .A(_02447_),
    .ZN(_02448_)
  );
  AND2_X1 _36642_ (
    .A1(_21197_),
    .A2(_21979_),
    .ZN(_02449_)
  );
  INV_X1 _36643_ (
    .A(_02449_),
    .ZN(_02450_)
  );
  AND2_X1 _36644_ (
    .A1(_02448_),
    .A2(_02450_),
    .ZN(_02451_)
  );
  INV_X1 _36645_ (
    .A(_02451_),
    .ZN(_02452_)
  );
  AND2_X1 _36646_ (
    .A1(_02446_),
    .A2(_02451_),
    .ZN(_02453_)
  );
  INV_X1 _36647_ (
    .A(_02453_),
    .ZN(_02454_)
  );
  AND2_X1 _36648_ (
    .A1(_02445_),
    .A2(_02452_),
    .ZN(_02455_)
  );
  INV_X1 _36649_ (
    .A(_02455_),
    .ZN(_02456_)
  );
  AND2_X1 _36650_ (
    .A1(_22559_),
    .A2(_02456_),
    .ZN(_02457_)
  );
  AND2_X1 _36651_ (
    .A1(_02454_),
    .A2(_02457_),
    .ZN(_02458_)
  );
  INV_X1 _36652_ (
    .A(_02458_),
    .ZN(_02459_)
  );
  AND2_X1 _36653_ (
    .A1(_02444_),
    .A2(_02459_),
    .ZN(_02460_)
  );
  INV_X1 _36654_ (
    .A(_02460_),
    .ZN(_02461_)
  );
  AND2_X1 _36655_ (
    .A1(_02260_),
    .A2(_02461_),
    .ZN(_00087_)
  );
  AND2_X1 _36656_ (
    .A1(_22035_),
    .A2(_22059_),
    .ZN(_02462_)
  );
  AND2_X1 _36657_ (
    .A1(_22251_),
    .A2(_02462_),
    .ZN(_02463_)
  );
  AND2_X1 _36658_ (
    .A1(_22268_),
    .A2(_02463_),
    .ZN(_02464_)
  );
  INV_X1 _36659_ (
    .A(_02464_),
    .ZN(_02465_)
  );
  AND2_X1 _36660_ (
    .A1(decoder_trigger),
    .A2(_02464_),
    .ZN(_02466_)
  );
  AND2_X1 _36661_ (
    .A1(_21167_),
    .A2(_02466_),
    .ZN(_02467_)
  );
  INV_X1 _36662_ (
    .A(_02467_),
    .ZN(_02468_)
  );
  AND2_X1 _36663_ (
    .A1(resetn),
    .A2(_02466_),
    .ZN(_02469_)
  );
  INV_X1 _36664_ (
    .A(_02469_),
    .ZN(_02470_)
  );
  AND2_X1 _36665_ (
    .A1(count_instr[0]),
    .A2(resetn),
    .ZN(_02471_)
  );
  INV_X1 _36666_ (
    .A(_02471_),
    .ZN(_02472_)
  );
  AND2_X1 _36667_ (
    .A1(_02470_),
    .A2(_02472_),
    .ZN(_02473_)
  );
  INV_X1 _36668_ (
    .A(_02473_),
    .ZN(_02474_)
  );
  AND2_X1 _36669_ (
    .A1(_02468_),
    .A2(_02474_),
    .ZN(_00088_)
  );
  AND2_X1 _36670_ (
    .A1(count_instr[0]),
    .A2(_02466_),
    .ZN(_02475_)
  );
  INV_X1 _36671_ (
    .A(_02475_),
    .ZN(_02476_)
  );
  AND2_X1 _36672_ (
    .A1(count_instr[1]),
    .A2(count_instr[0]),
    .ZN(_02477_)
  );
  AND2_X1 _36673_ (
    .A1(_02466_),
    .A2(_02477_),
    .ZN(_02478_)
  );
  INV_X1 _36674_ (
    .A(_02478_),
    .ZN(_02479_)
  );
  AND2_X1 _36675_ (
    .A1(_21166_),
    .A2(_02476_),
    .ZN(_02480_)
  );
  INV_X1 _36676_ (
    .A(_02480_),
    .ZN(_02481_)
  );
  AND2_X1 _36677_ (
    .A1(resetn),
    .A2(_02481_),
    .ZN(_02482_)
  );
  AND2_X1 _36678_ (
    .A1(_02479_),
    .A2(_02482_),
    .ZN(_00089_)
  );
  AND2_X1 _36679_ (
    .A1(count_instr[2]),
    .A2(_02478_),
    .ZN(_02483_)
  );
  INV_X1 _36680_ (
    .A(_02483_),
    .ZN(_02484_)
  );
  AND2_X1 _36681_ (
    .A1(_21165_),
    .A2(_02479_),
    .ZN(_02485_)
  );
  INV_X1 _36682_ (
    .A(_02485_),
    .ZN(_02486_)
  );
  AND2_X1 _36683_ (
    .A1(resetn),
    .A2(_02486_),
    .ZN(_02487_)
  );
  AND2_X1 _36684_ (
    .A1(_02484_),
    .A2(_02487_),
    .ZN(_00090_)
  );
  AND2_X1 _36685_ (
    .A1(_21164_),
    .A2(_02484_),
    .ZN(_02488_)
  );
  INV_X1 _36686_ (
    .A(_02488_),
    .ZN(_02489_)
  );
  AND2_X1 _36687_ (
    .A1(count_instr[3]),
    .A2(count_instr[2]),
    .ZN(_02490_)
  );
  AND2_X1 _36688_ (
    .A1(_02477_),
    .A2(_02490_),
    .ZN(_02491_)
  );
  AND2_X1 _36689_ (
    .A1(_02466_),
    .A2(_02491_),
    .ZN(_02492_)
  );
  INV_X1 _36690_ (
    .A(_02492_),
    .ZN(_02493_)
  );
  AND2_X1 _36691_ (
    .A1(resetn),
    .A2(_02493_),
    .ZN(_02494_)
  );
  AND2_X1 _36692_ (
    .A1(_02489_),
    .A2(_02494_),
    .ZN(_00091_)
  );
  AND2_X1 _36693_ (
    .A1(count_instr[4]),
    .A2(_02492_),
    .ZN(_02495_)
  );
  INV_X1 _36694_ (
    .A(_02495_),
    .ZN(_02496_)
  );
  AND2_X1 _36695_ (
    .A1(_21163_),
    .A2(_02493_),
    .ZN(_02497_)
  );
  INV_X1 _36696_ (
    .A(_02497_),
    .ZN(_02498_)
  );
  AND2_X1 _36697_ (
    .A1(resetn),
    .A2(_02498_),
    .ZN(_02499_)
  );
  AND2_X1 _36698_ (
    .A1(_02496_),
    .A2(_02499_),
    .ZN(_00092_)
  );
  AND2_X1 _36699_ (
    .A1(_21162_),
    .A2(_02496_),
    .ZN(_02500_)
  );
  INV_X1 _36700_ (
    .A(_02500_),
    .ZN(_02501_)
  );
  AND2_X1 _36701_ (
    .A1(count_instr[5]),
    .A2(count_instr[4]),
    .ZN(_02502_)
  );
  AND2_X1 _36702_ (
    .A1(_02492_),
    .A2(_02502_),
    .ZN(_02503_)
  );
  INV_X1 _36703_ (
    .A(_02503_),
    .ZN(_02504_)
  );
  AND2_X1 _36704_ (
    .A1(resetn),
    .A2(_02504_),
    .ZN(_02505_)
  );
  AND2_X1 _36705_ (
    .A1(_02501_),
    .A2(_02505_),
    .ZN(_00093_)
  );
  AND2_X1 _36706_ (
    .A1(_21161_),
    .A2(_02504_),
    .ZN(_02506_)
  );
  INV_X1 _36707_ (
    .A(_02506_),
    .ZN(_02507_)
  );
  AND2_X1 _36708_ (
    .A1(resetn),
    .A2(_02507_),
    .ZN(_02508_)
  );
  AND2_X1 _36709_ (
    .A1(count_instr[6]),
    .A2(_02503_),
    .ZN(_02509_)
  );
  INV_X1 _36710_ (
    .A(_02509_),
    .ZN(_02510_)
  );
  AND2_X1 _36711_ (
    .A1(_02508_),
    .A2(_02510_),
    .ZN(_00094_)
  );
  AND2_X1 _36712_ (
    .A1(_21160_),
    .A2(_02510_),
    .ZN(_02511_)
  );
  INV_X1 _36713_ (
    .A(_02511_),
    .ZN(_02512_)
  );
  AND2_X1 _36714_ (
    .A1(count_instr[7]),
    .A2(count_instr[6]),
    .ZN(_02513_)
  );
  AND2_X1 _36715_ (
    .A1(_02503_),
    .A2(_02513_),
    .ZN(_02514_)
  );
  AND2_X1 _36716_ (
    .A1(resetn),
    .A2(_02512_),
    .ZN(_02515_)
  );
  AND2_X1 _36717_ (
    .A1(count_instr[7]),
    .A2(_02502_),
    .ZN(_02516_)
  );
  AND2_X1 _36718_ (
    .A1(count_instr[6]),
    .A2(_02516_),
    .ZN(_02517_)
  );
  AND2_X1 _36719_ (
    .A1(_02491_),
    .A2(_02517_),
    .ZN(_02518_)
  );
  AND2_X1 _36720_ (
    .A1(_02466_),
    .A2(_02518_),
    .ZN(_02519_)
  );
  AND2_X1 _36721_ (
    .A1(_02492_),
    .A2(_02517_),
    .ZN(_02520_)
  );
  INV_X1 _36722_ (
    .A(_02520_),
    .ZN(_02521_)
  );
  AND2_X1 _36723_ (
    .A1(_02515_),
    .A2(_02521_),
    .ZN(_00095_)
  );
  AND2_X1 _36724_ (
    .A1(_21159_),
    .A2(_02521_),
    .ZN(_02522_)
  );
  INV_X1 _36725_ (
    .A(_02522_),
    .ZN(_02523_)
  );
  AND2_X1 _36726_ (
    .A1(resetn),
    .A2(_02523_),
    .ZN(_02524_)
  );
  AND2_X1 _36727_ (
    .A1(count_instr[8]),
    .A2(_02519_),
    .ZN(_02525_)
  );
  INV_X1 _36728_ (
    .A(_02525_),
    .ZN(_02526_)
  );
  AND2_X1 _36729_ (
    .A1(_02524_),
    .A2(_02526_),
    .ZN(_00096_)
  );
  AND2_X1 _36730_ (
    .A1(_21158_),
    .A2(_02526_),
    .ZN(_02527_)
  );
  INV_X1 _36731_ (
    .A(_02527_),
    .ZN(_02528_)
  );
  AND2_X1 _36732_ (
    .A1(count_instr[9]),
    .A2(count_instr[8]),
    .ZN(_02529_)
  );
  AND2_X1 _36733_ (
    .A1(_02514_),
    .A2(_02529_),
    .ZN(_02530_)
  );
  INV_X1 _36734_ (
    .A(_02530_),
    .ZN(_02531_)
  );
  AND2_X1 _36735_ (
    .A1(resetn),
    .A2(_02531_),
    .ZN(_02532_)
  );
  AND2_X1 _36736_ (
    .A1(_02528_),
    .A2(_02532_),
    .ZN(_00097_)
  );
  AND2_X1 _36737_ (
    .A1(_21157_),
    .A2(_02531_),
    .ZN(_02533_)
  );
  INV_X1 _36738_ (
    .A(_02533_),
    .ZN(_02534_)
  );
  AND2_X1 _36739_ (
    .A1(resetn),
    .A2(_02534_),
    .ZN(_02535_)
  );
  AND2_X1 _36740_ (
    .A1(count_instr[10]),
    .A2(_02530_),
    .ZN(_02536_)
  );
  INV_X1 _36741_ (
    .A(_02536_),
    .ZN(_02537_)
  );
  AND2_X1 _36742_ (
    .A1(_02535_),
    .A2(_02537_),
    .ZN(_00098_)
  );
  AND2_X1 _36743_ (
    .A1(_21156_),
    .A2(_02537_),
    .ZN(_02538_)
  );
  INV_X1 _36744_ (
    .A(_02538_),
    .ZN(_02539_)
  );
  AND2_X1 _36745_ (
    .A1(resetn),
    .A2(_02539_),
    .ZN(_02540_)
  );
  AND2_X1 _36746_ (
    .A1(count_instr[11]),
    .A2(_02536_),
    .ZN(_02541_)
  );
  INV_X1 _36747_ (
    .A(_02541_),
    .ZN(_02542_)
  );
  AND2_X1 _36748_ (
    .A1(count_instr[11]),
    .A2(count_instr[10]),
    .ZN(_02543_)
  );
  AND2_X1 _36749_ (
    .A1(_02540_),
    .A2(_02542_),
    .ZN(_00099_)
  );
  AND2_X1 _36750_ (
    .A1(_21155_),
    .A2(_02542_),
    .ZN(_02544_)
  );
  INV_X1 _36751_ (
    .A(_02544_),
    .ZN(_02545_)
  );
  AND2_X1 _36752_ (
    .A1(resetn),
    .A2(_02545_),
    .ZN(_02546_)
  );
  AND2_X1 _36753_ (
    .A1(count_instr[12]),
    .A2(_02541_),
    .ZN(_02547_)
  );
  INV_X1 _36754_ (
    .A(_02547_),
    .ZN(_02548_)
  );
  AND2_X1 _36755_ (
    .A1(_02546_),
    .A2(_02548_),
    .ZN(_00100_)
  );
  AND2_X1 _36756_ (
    .A1(_21154_),
    .A2(_02548_),
    .ZN(_02549_)
  );
  INV_X1 _36757_ (
    .A(_02549_),
    .ZN(_02550_)
  );
  AND2_X1 _36758_ (
    .A1(count_instr[13]),
    .A2(count_instr[12]),
    .ZN(_02551_)
  );
  AND2_X1 _36759_ (
    .A1(_02543_),
    .A2(_02551_),
    .ZN(_02552_)
  );
  AND2_X1 _36760_ (
    .A1(_02530_),
    .A2(_02552_),
    .ZN(_02553_)
  );
  INV_X1 _36761_ (
    .A(_02553_),
    .ZN(_02554_)
  );
  AND2_X1 _36762_ (
    .A1(resetn),
    .A2(_02554_),
    .ZN(_02555_)
  );
  AND2_X1 _36763_ (
    .A1(_02550_),
    .A2(_02555_),
    .ZN(_00101_)
  );
  AND2_X1 _36764_ (
    .A1(_02529_),
    .A2(_02552_),
    .ZN(_02556_)
  );
  AND2_X1 _36765_ (
    .A1(_02519_),
    .A2(_02556_),
    .ZN(_02557_)
  );
  AND2_X1 _36766_ (
    .A1(count_instr[13]),
    .A2(_02517_),
    .ZN(_02558_)
  );
  AND2_X1 _36767_ (
    .A1(_02529_),
    .A2(_02543_),
    .ZN(_02559_)
  );
  AND2_X1 _36768_ (
    .A1(_02491_),
    .A2(_02559_),
    .ZN(_02560_)
  );
  AND2_X1 _36769_ (
    .A1(count_instr[12]),
    .A2(_02560_),
    .ZN(_02561_)
  );
  AND2_X1 _36770_ (
    .A1(_02558_),
    .A2(_02561_),
    .ZN(_02562_)
  );
  AND2_X1 _36771_ (
    .A1(_02466_),
    .A2(_02562_),
    .ZN(_02563_)
  );
  AND2_X1 _36772_ (
    .A1(_21153_),
    .A2(_02554_),
    .ZN(_02564_)
  );
  INV_X1 _36773_ (
    .A(_02564_),
    .ZN(_02565_)
  );
  AND2_X1 _36774_ (
    .A1(resetn),
    .A2(_02565_),
    .ZN(_02566_)
  );
  AND2_X1 _36775_ (
    .A1(count_instr[14]),
    .A2(_02553_),
    .ZN(_02567_)
  );
  INV_X1 _36776_ (
    .A(_02567_),
    .ZN(_02568_)
  );
  AND2_X1 _36777_ (
    .A1(count_instr[14]),
    .A2(_02557_),
    .ZN(_02569_)
  );
  AND2_X1 _36778_ (
    .A1(_02566_),
    .A2(_02568_),
    .ZN(_00102_)
  );
  AND2_X1 _36779_ (
    .A1(_21152_),
    .A2(_02568_),
    .ZN(_02570_)
  );
  INV_X1 _36780_ (
    .A(_02570_),
    .ZN(_02571_)
  );
  AND2_X1 _36781_ (
    .A1(count_instr[15]),
    .A2(count_instr[14]),
    .ZN(_02572_)
  );
  AND2_X1 _36782_ (
    .A1(resetn),
    .A2(_02571_),
    .ZN(_02573_)
  );
  AND2_X1 _36783_ (
    .A1(count_instr[15]),
    .A2(_02569_),
    .ZN(_02574_)
  );
  INV_X1 _36784_ (
    .A(_02574_),
    .ZN(_02575_)
  );
  AND2_X1 _36785_ (
    .A1(_02573_),
    .A2(_02575_),
    .ZN(_00103_)
  );
  AND2_X1 _36786_ (
    .A1(_21151_),
    .A2(_02575_),
    .ZN(_02576_)
  );
  INV_X1 _36787_ (
    .A(_02576_),
    .ZN(_02577_)
  );
  AND2_X1 _36788_ (
    .A1(resetn),
    .A2(_02577_),
    .ZN(_02578_)
  );
  AND2_X1 _36789_ (
    .A1(count_instr[16]),
    .A2(_02574_),
    .ZN(_02579_)
  );
  INV_X1 _36790_ (
    .A(_02579_),
    .ZN(_02580_)
  );
  AND2_X1 _36791_ (
    .A1(count_instr[16]),
    .A2(_02572_),
    .ZN(_02581_)
  );
  AND2_X1 _36792_ (
    .A1(_02578_),
    .A2(_02580_),
    .ZN(_00104_)
  );
  AND2_X1 _36793_ (
    .A1(_21150_),
    .A2(_02580_),
    .ZN(_02582_)
  );
  INV_X1 _36794_ (
    .A(_02582_),
    .ZN(_02583_)
  );
  AND2_X1 _36795_ (
    .A1(resetn),
    .A2(_02583_),
    .ZN(_02584_)
  );
  AND2_X1 _36796_ (
    .A1(count_instr[17]),
    .A2(_02579_),
    .ZN(_02585_)
  );
  INV_X1 _36797_ (
    .A(_02585_),
    .ZN(_02586_)
  );
  AND2_X1 _36798_ (
    .A1(_02584_),
    .A2(_02586_),
    .ZN(_00105_)
  );
  AND2_X1 _36799_ (
    .A1(_21149_),
    .A2(_02586_),
    .ZN(_02587_)
  );
  INV_X1 _36800_ (
    .A(_02587_),
    .ZN(_02588_)
  );
  AND2_X1 _36801_ (
    .A1(resetn),
    .A2(_02588_),
    .ZN(_02589_)
  );
  AND2_X1 _36802_ (
    .A1(count_instr[18]),
    .A2(_02585_),
    .ZN(_02590_)
  );
  INV_X1 _36803_ (
    .A(_02590_),
    .ZN(_02591_)
  );
  AND2_X1 _36804_ (
    .A1(_02589_),
    .A2(_02591_),
    .ZN(_00106_)
  );
  AND2_X1 _36805_ (
    .A1(_21148_),
    .A2(_02591_),
    .ZN(_02592_)
  );
  INV_X1 _36806_ (
    .A(_02592_),
    .ZN(_02593_)
  );
  AND2_X1 _36807_ (
    .A1(count_instr[18]),
    .A2(count_instr[17]),
    .ZN(_02594_)
  );
  AND2_X1 _36808_ (
    .A1(count_instr[19]),
    .A2(_02594_),
    .ZN(_02595_)
  );
  AND2_X1 _36809_ (
    .A1(_02581_),
    .A2(_02595_),
    .ZN(_02596_)
  );
  AND2_X1 _36810_ (
    .A1(_02553_),
    .A2(_02596_),
    .ZN(_02597_)
  );
  AND2_X1 _36811_ (
    .A1(resetn),
    .A2(_02593_),
    .ZN(_02598_)
  );
  AND2_X1 _36812_ (
    .A1(count_instr[19]),
    .A2(_02590_),
    .ZN(_02599_)
  );
  INV_X1 _36813_ (
    .A(_02599_),
    .ZN(_02600_)
  );
  AND2_X1 _36814_ (
    .A1(_02598_),
    .A2(_02600_),
    .ZN(_00107_)
  );
  AND2_X1 _36815_ (
    .A1(_21147_),
    .A2(_02600_),
    .ZN(_02601_)
  );
  INV_X1 _36816_ (
    .A(_02601_),
    .ZN(_02602_)
  );
  AND2_X1 _36817_ (
    .A1(resetn),
    .A2(_02602_),
    .ZN(_02603_)
  );
  AND2_X1 _36818_ (
    .A1(count_instr[20]),
    .A2(_02597_),
    .ZN(_02604_)
  );
  INV_X1 _36819_ (
    .A(_02604_),
    .ZN(_02605_)
  );
  AND2_X1 _36820_ (
    .A1(_02603_),
    .A2(_02605_),
    .ZN(_00108_)
  );
  AND2_X1 _36821_ (
    .A1(_21146_),
    .A2(_02605_),
    .ZN(_02606_)
  );
  INV_X1 _36822_ (
    .A(_02606_),
    .ZN(_02607_)
  );
  AND2_X1 _36823_ (
    .A1(resetn),
    .A2(_02607_),
    .ZN(_02608_)
  );
  AND2_X1 _36824_ (
    .A1(count_instr[21]),
    .A2(_02604_),
    .ZN(_02609_)
  );
  INV_X1 _36825_ (
    .A(_02609_),
    .ZN(_02610_)
  );
  AND2_X1 _36826_ (
    .A1(count_instr[21]),
    .A2(count_instr[20]),
    .ZN(_02611_)
  );
  AND2_X1 _36827_ (
    .A1(_02608_),
    .A2(_02610_),
    .ZN(_00109_)
  );
  AND2_X1 _36828_ (
    .A1(_21145_),
    .A2(_02610_),
    .ZN(_02612_)
  );
  INV_X1 _36829_ (
    .A(_02612_),
    .ZN(_02613_)
  );
  AND2_X1 _36830_ (
    .A1(resetn),
    .A2(_02613_),
    .ZN(_02614_)
  );
  AND2_X1 _36831_ (
    .A1(count_instr[22]),
    .A2(_02609_),
    .ZN(_02615_)
  );
  INV_X1 _36832_ (
    .A(_02615_),
    .ZN(_02616_)
  );
  AND2_X1 _36833_ (
    .A1(_02614_),
    .A2(_02616_),
    .ZN(_00110_)
  );
  AND2_X1 _36834_ (
    .A1(_21144_),
    .A2(_02616_),
    .ZN(_02617_)
  );
  INV_X1 _36835_ (
    .A(_02617_),
    .ZN(_02618_)
  );
  AND2_X1 _36836_ (
    .A1(count_instr[23]),
    .A2(count_instr[22]),
    .ZN(_02619_)
  );
  AND2_X1 _36837_ (
    .A1(count_instr[21]),
    .A2(_02619_),
    .ZN(_02620_)
  );
  AND2_X1 _36838_ (
    .A1(_02604_),
    .A2(_02620_),
    .ZN(_02621_)
  );
  INV_X1 _36839_ (
    .A(_02621_),
    .ZN(_02622_)
  );
  AND2_X1 _36840_ (
    .A1(resetn),
    .A2(_02622_),
    .ZN(_02623_)
  );
  AND2_X1 _36841_ (
    .A1(count_instr[23]),
    .A2(_02611_),
    .ZN(_02624_)
  );
  AND2_X1 _36842_ (
    .A1(count_instr[22]),
    .A2(_02624_),
    .ZN(_02625_)
  );
  AND2_X1 _36843_ (
    .A1(_02618_),
    .A2(_02623_),
    .ZN(_00111_)
  );
  AND2_X1 _36844_ (
    .A1(_02596_),
    .A2(_02625_),
    .ZN(_02626_)
  );
  AND2_X1 _36845_ (
    .A1(_02557_),
    .A2(_02626_),
    .ZN(_02627_)
  );
  AND2_X1 _36846_ (
    .A1(count_instr[22]),
    .A2(_02595_),
    .ZN(_02628_)
  );
  AND2_X1 _36847_ (
    .A1(_02581_),
    .A2(_02624_),
    .ZN(_02629_)
  );
  AND2_X1 _36848_ (
    .A1(_02628_),
    .A2(_02629_),
    .ZN(_02630_)
  );
  AND2_X1 _36849_ (
    .A1(_21143_),
    .A2(_02622_),
    .ZN(_02631_)
  );
  INV_X1 _36850_ (
    .A(_02631_),
    .ZN(_02632_)
  );
  AND2_X1 _36851_ (
    .A1(resetn),
    .A2(_02632_),
    .ZN(_02633_)
  );
  AND2_X1 _36852_ (
    .A1(count_instr[24]),
    .A2(_02621_),
    .ZN(_02634_)
  );
  INV_X1 _36853_ (
    .A(_02634_),
    .ZN(_02635_)
  );
  AND2_X1 _36854_ (
    .A1(_02633_),
    .A2(_02635_),
    .ZN(_00112_)
  );
  AND2_X1 _36855_ (
    .A1(_21142_),
    .A2(_02635_),
    .ZN(_02636_)
  );
  INV_X1 _36856_ (
    .A(_02636_),
    .ZN(_02637_)
  );
  AND2_X1 _36857_ (
    .A1(resetn),
    .A2(_02637_),
    .ZN(_02638_)
  );
  AND2_X1 _36858_ (
    .A1(count_instr[25]),
    .A2(_02634_),
    .ZN(_02639_)
  );
  INV_X1 _36859_ (
    .A(_02639_),
    .ZN(_02640_)
  );
  AND2_X1 _36860_ (
    .A1(count_instr[25]),
    .A2(count_instr[24]),
    .ZN(_02641_)
  );
  AND2_X1 _36861_ (
    .A1(_02627_),
    .A2(_02641_),
    .ZN(_02642_)
  );
  AND2_X1 _36862_ (
    .A1(_02638_),
    .A2(_02640_),
    .ZN(_00113_)
  );
  AND2_X1 _36863_ (
    .A1(_21141_),
    .A2(_02640_),
    .ZN(_02643_)
  );
  INV_X1 _36864_ (
    .A(_02643_),
    .ZN(_02644_)
  );
  AND2_X1 _36865_ (
    .A1(resetn),
    .A2(_02644_),
    .ZN(_02645_)
  );
  AND2_X1 _36866_ (
    .A1(count_instr[26]),
    .A2(_02639_),
    .ZN(_02646_)
  );
  INV_X1 _36867_ (
    .A(_02646_),
    .ZN(_02647_)
  );
  AND2_X1 _36868_ (
    .A1(count_instr[26]),
    .A2(_02642_),
    .ZN(_02648_)
  );
  AND2_X1 _36869_ (
    .A1(_02645_),
    .A2(_02647_),
    .ZN(_00114_)
  );
  AND2_X1 _36870_ (
    .A1(_21140_),
    .A2(_02647_),
    .ZN(_02649_)
  );
  INV_X1 _36871_ (
    .A(_02649_),
    .ZN(_02650_)
  );
  AND2_X1 _36872_ (
    .A1(count_instr[27]),
    .A2(count_instr[26]),
    .ZN(_02651_)
  );
  AND2_X1 _36873_ (
    .A1(_02639_),
    .A2(_02651_),
    .ZN(_02652_)
  );
  INV_X1 _36874_ (
    .A(_02652_),
    .ZN(_02653_)
  );
  AND2_X1 _36875_ (
    .A1(resetn),
    .A2(_02653_),
    .ZN(_02654_)
  );
  AND2_X1 _36876_ (
    .A1(count_instr[27]),
    .A2(_02648_),
    .ZN(_02655_)
  );
  AND2_X1 _36877_ (
    .A1(_02650_),
    .A2(_02654_),
    .ZN(_00115_)
  );
  AND2_X1 _36878_ (
    .A1(_21139_),
    .A2(_02653_),
    .ZN(_02656_)
  );
  INV_X1 _36879_ (
    .A(_02656_),
    .ZN(_02657_)
  );
  AND2_X1 _36880_ (
    .A1(resetn),
    .A2(_02657_),
    .ZN(_02658_)
  );
  AND2_X1 _36881_ (
    .A1(count_instr[28]),
    .A2(_02652_),
    .ZN(_02659_)
  );
  INV_X1 _36882_ (
    .A(_02659_),
    .ZN(_02660_)
  );
  AND2_X1 _36883_ (
    .A1(count_instr[28]),
    .A2(_02655_),
    .ZN(_02661_)
  );
  AND2_X1 _36884_ (
    .A1(_02658_),
    .A2(_02660_),
    .ZN(_00116_)
  );
  AND2_X1 _36885_ (
    .A1(_21138_),
    .A2(_02660_),
    .ZN(_02662_)
  );
  INV_X1 _36886_ (
    .A(_02662_),
    .ZN(_02663_)
  );
  AND2_X1 _36887_ (
    .A1(count_instr[29]),
    .A2(count_instr[28]),
    .ZN(_02664_)
  );
  AND2_X1 _36888_ (
    .A1(_02651_),
    .A2(_02664_),
    .ZN(_02665_)
  );
  AND2_X1 _36889_ (
    .A1(resetn),
    .A2(_02663_),
    .ZN(_02666_)
  );
  AND2_X1 _36890_ (
    .A1(count_instr[29]),
    .A2(_02661_),
    .ZN(_02667_)
  );
  INV_X1 _36891_ (
    .A(_02667_),
    .ZN(_02668_)
  );
  AND2_X1 _36892_ (
    .A1(_02666_),
    .A2(_02668_),
    .ZN(_00117_)
  );
  AND2_X1 _36893_ (
    .A1(_21137_),
    .A2(_02668_),
    .ZN(_02669_)
  );
  INV_X1 _36894_ (
    .A(_02669_),
    .ZN(_02670_)
  );
  AND2_X1 _36895_ (
    .A1(resetn),
    .A2(_02670_),
    .ZN(_02671_)
  );
  AND2_X1 _36896_ (
    .A1(count_instr[30]),
    .A2(_02667_),
    .ZN(_02672_)
  );
  INV_X1 _36897_ (
    .A(_02672_),
    .ZN(_02673_)
  );
  AND2_X1 _36898_ (
    .A1(_02671_),
    .A2(_02673_),
    .ZN(_00118_)
  );
  AND2_X1 _36899_ (
    .A1(_21136_),
    .A2(_02673_),
    .ZN(_02674_)
  );
  INV_X1 _36900_ (
    .A(_02674_),
    .ZN(_02675_)
  );
  AND2_X1 _36901_ (
    .A1(count_instr[31]),
    .A2(count_instr[30]),
    .ZN(_02676_)
  );
  AND2_X1 _36902_ (
    .A1(count_instr[25]),
    .A2(_02676_),
    .ZN(_02677_)
  );
  AND2_X1 _36903_ (
    .A1(_02665_),
    .A2(_02677_),
    .ZN(_02678_)
  );
  AND2_X1 _36904_ (
    .A1(_02634_),
    .A2(_02678_),
    .ZN(_02679_)
  );
  AND2_X1 _36905_ (
    .A1(resetn),
    .A2(_02675_),
    .ZN(_02680_)
  );
  AND2_X1 _36906_ (
    .A1(count_instr[31]),
    .A2(_02664_),
    .ZN(_02681_)
  );
  AND2_X1 _36907_ (
    .A1(count_instr[30]),
    .A2(_02681_),
    .ZN(_02682_)
  );
  AND2_X1 _36908_ (
    .A1(_02651_),
    .A2(_02682_),
    .ZN(_02683_)
  );
  AND2_X1 _36909_ (
    .A1(_02641_),
    .A2(_02683_),
    .ZN(_02684_)
  );
  AND2_X1 _36910_ (
    .A1(_02627_),
    .A2(_02684_),
    .ZN(_02685_)
  );
  INV_X1 _36911_ (
    .A(_02685_),
    .ZN(_02686_)
  );
  AND2_X1 _36912_ (
    .A1(_02630_),
    .A2(_02684_),
    .ZN(_02687_)
  );
  AND2_X1 _36913_ (
    .A1(_02563_),
    .A2(_02687_),
    .ZN(_02688_)
  );
  AND2_X1 _36914_ (
    .A1(_02680_),
    .A2(_02686_),
    .ZN(_00119_)
  );
  AND2_X1 _36915_ (
    .A1(_21135_),
    .A2(_02686_),
    .ZN(_02689_)
  );
  INV_X1 _36916_ (
    .A(_02689_),
    .ZN(_02690_)
  );
  AND2_X1 _36917_ (
    .A1(resetn),
    .A2(_02690_),
    .ZN(_02691_)
  );
  AND2_X1 _36918_ (
    .A1(count_instr[32]),
    .A2(_02685_),
    .ZN(_02692_)
  );
  INV_X1 _36919_ (
    .A(_02692_),
    .ZN(_02693_)
  );
  AND2_X1 _36920_ (
    .A1(count_instr[32]),
    .A2(_02688_),
    .ZN(_02694_)
  );
  AND2_X1 _36921_ (
    .A1(_02691_),
    .A2(_02693_),
    .ZN(_00120_)
  );
  AND2_X1 _36922_ (
    .A1(_21134_),
    .A2(_02693_),
    .ZN(_02695_)
  );
  INV_X1 _36923_ (
    .A(_02695_),
    .ZN(_02696_)
  );
  AND2_X1 _36924_ (
    .A1(count_instr[33]),
    .A2(count_instr[32]),
    .ZN(_02697_)
  );
  AND2_X1 _36925_ (
    .A1(resetn),
    .A2(_02696_),
    .ZN(_02698_)
  );
  AND2_X1 _36926_ (
    .A1(count_instr[33]),
    .A2(_02692_),
    .ZN(_02699_)
  );
  INV_X1 _36927_ (
    .A(_02699_),
    .ZN(_02700_)
  );
  AND2_X1 _36928_ (
    .A1(_02698_),
    .A2(_02700_),
    .ZN(_00121_)
  );
  AND2_X1 _36929_ (
    .A1(_21133_),
    .A2(_02700_),
    .ZN(_02701_)
  );
  INV_X1 _36930_ (
    .A(_02701_),
    .ZN(_02702_)
  );
  AND2_X1 _36931_ (
    .A1(resetn),
    .A2(_02702_),
    .ZN(_02703_)
  );
  AND2_X1 _36932_ (
    .A1(count_instr[34]),
    .A2(_02699_),
    .ZN(_02704_)
  );
  INV_X1 _36933_ (
    .A(_02704_),
    .ZN(_02705_)
  );
  AND2_X1 _36934_ (
    .A1(count_instr[34]),
    .A2(count_instr[33]),
    .ZN(_02706_)
  );
  AND2_X1 _36935_ (
    .A1(_02703_),
    .A2(_02705_),
    .ZN(_00122_)
  );
  AND2_X1 _36936_ (
    .A1(_21132_),
    .A2(_02705_),
    .ZN(_02707_)
  );
  INV_X1 _36937_ (
    .A(_02707_),
    .ZN(_02708_)
  );
  AND2_X1 _36938_ (
    .A1(count_instr[35]),
    .A2(count_instr[34]),
    .ZN(_02709_)
  );
  AND2_X1 _36939_ (
    .A1(_02697_),
    .A2(_02709_),
    .ZN(_02710_)
  );
  AND2_X1 _36940_ (
    .A1(_02679_),
    .A2(_02710_),
    .ZN(_02711_)
  );
  AND2_X1 _36941_ (
    .A1(resetn),
    .A2(_02708_),
    .ZN(_02712_)
  );
  AND2_X1 _36942_ (
    .A1(count_instr[35]),
    .A2(_02704_),
    .ZN(_02713_)
  );
  INV_X1 _36943_ (
    .A(_02713_),
    .ZN(_02714_)
  );
  AND2_X1 _36944_ (
    .A1(count_instr[35]),
    .A2(_02706_),
    .ZN(_02715_)
  );
  AND2_X1 _36945_ (
    .A1(_02694_),
    .A2(_02715_),
    .ZN(_02716_)
  );
  AND2_X1 _36946_ (
    .A1(_02712_),
    .A2(_02714_),
    .ZN(_00123_)
  );
  AND2_X1 _36947_ (
    .A1(_21131_),
    .A2(_02714_),
    .ZN(_02717_)
  );
  INV_X1 _36948_ (
    .A(_02717_),
    .ZN(_02718_)
  );
  AND2_X1 _36949_ (
    .A1(resetn),
    .A2(_02718_),
    .ZN(_02719_)
  );
  AND2_X1 _36950_ (
    .A1(count_instr[36]),
    .A2(_02711_),
    .ZN(_02720_)
  );
  AND2_X1 _36951_ (
    .A1(count_instr[36]),
    .A2(_02713_),
    .ZN(_02721_)
  );
  INV_X1 _36952_ (
    .A(_02721_),
    .ZN(_02722_)
  );
  AND2_X1 _36953_ (
    .A1(count_instr[36]),
    .A2(_02716_),
    .ZN(_02723_)
  );
  AND2_X1 _36954_ (
    .A1(_02719_),
    .A2(_02722_),
    .ZN(_00124_)
  );
  AND2_X1 _36955_ (
    .A1(_21130_),
    .A2(_02722_),
    .ZN(_02724_)
  );
  INV_X1 _36956_ (
    .A(_02724_),
    .ZN(_02725_)
  );
  AND2_X1 _36957_ (
    .A1(resetn),
    .A2(_02725_),
    .ZN(_02726_)
  );
  AND2_X1 _36958_ (
    .A1(count_instr[37]),
    .A2(count_instr[36]),
    .ZN(_02727_)
  );
  AND2_X1 _36959_ (
    .A1(count_instr[37]),
    .A2(_02723_),
    .ZN(_02728_)
  );
  INV_X1 _36960_ (
    .A(_02728_),
    .ZN(_02729_)
  );
  AND2_X1 _36961_ (
    .A1(_02726_),
    .A2(_02729_),
    .ZN(_00125_)
  );
  AND2_X1 _36962_ (
    .A1(_21129_),
    .A2(_02729_),
    .ZN(_02730_)
  );
  INV_X1 _36963_ (
    .A(_02730_),
    .ZN(_02731_)
  );
  AND2_X1 _36964_ (
    .A1(resetn),
    .A2(_02731_),
    .ZN(_02732_)
  );
  AND2_X1 _36965_ (
    .A1(count_instr[38]),
    .A2(_02728_),
    .ZN(_02733_)
  );
  INV_X1 _36966_ (
    .A(_02733_),
    .ZN(_02734_)
  );
  AND2_X1 _36967_ (
    .A1(_02732_),
    .A2(_02734_),
    .ZN(_00126_)
  );
  AND2_X1 _36968_ (
    .A1(_21128_),
    .A2(_02734_),
    .ZN(_02735_)
  );
  INV_X1 _36969_ (
    .A(_02735_),
    .ZN(_02736_)
  );
  AND2_X1 _36970_ (
    .A1(resetn),
    .A2(_02736_),
    .ZN(_02737_)
  );
  AND2_X1 _36971_ (
    .A1(count_instr[39]),
    .A2(_02733_),
    .ZN(_02738_)
  );
  INV_X1 _36972_ (
    .A(_02738_),
    .ZN(_02739_)
  );
  AND2_X1 _36973_ (
    .A1(_02737_),
    .A2(_02739_),
    .ZN(_00127_)
  );
  AND2_X1 _36974_ (
    .A1(count_instr[39]),
    .A2(count_instr[38]),
    .ZN(_02740_)
  );
  AND2_X1 _36975_ (
    .A1(count_instr[37]),
    .A2(_02740_),
    .ZN(_02741_)
  );
  AND2_X1 _36976_ (
    .A1(_02720_),
    .A2(_02741_),
    .ZN(_02742_)
  );
  AND2_X1 _36977_ (
    .A1(_02727_),
    .A2(_02740_),
    .ZN(_02743_)
  );
  AND2_X1 _36978_ (
    .A1(count_instr[32]),
    .A2(_02743_),
    .ZN(_02744_)
  );
  AND2_X1 _36979_ (
    .A1(_02715_),
    .A2(_02744_),
    .ZN(_02745_)
  );
  AND2_X1 _36980_ (
    .A1(_02685_),
    .A2(_02745_),
    .ZN(_02746_)
  );
  AND2_X1 _36981_ (
    .A1(count_instr[38]),
    .A2(_02687_),
    .ZN(_02747_)
  );
  AND2_X1 _36982_ (
    .A1(count_instr[39]),
    .A2(count_instr[32]),
    .ZN(_02748_)
  );
  AND2_X1 _36983_ (
    .A1(_02715_),
    .A2(_02748_),
    .ZN(_02749_)
  );
  AND2_X1 _36984_ (
    .A1(count_instr[37]),
    .A2(_02749_),
    .ZN(_02750_)
  );
  AND2_X1 _36985_ (
    .A1(count_instr[36]),
    .A2(_02750_),
    .ZN(_02751_)
  );
  AND2_X1 _36986_ (
    .A1(_02562_),
    .A2(_02751_),
    .ZN(_02752_)
  );
  AND2_X1 _36987_ (
    .A1(_02747_),
    .A2(_02752_),
    .ZN(_02753_)
  );
  AND2_X1 _36988_ (
    .A1(_02466_),
    .A2(_02753_),
    .ZN(_02754_)
  );
  INV_X1 _36989_ (
    .A(_02754_),
    .ZN(_02755_)
  );
  AND2_X1 _36990_ (
    .A1(_21127_),
    .A2(_02755_),
    .ZN(_02756_)
  );
  INV_X1 _36991_ (
    .A(_02756_),
    .ZN(_02757_)
  );
  AND2_X1 _36992_ (
    .A1(resetn),
    .A2(_02757_),
    .ZN(_02758_)
  );
  AND2_X1 _36993_ (
    .A1(count_instr[40]),
    .A2(_02742_),
    .ZN(_02759_)
  );
  INV_X1 _36994_ (
    .A(_02759_),
    .ZN(_02760_)
  );
  AND2_X1 _36995_ (
    .A1(_02758_),
    .A2(_02760_),
    .ZN(_00128_)
  );
  AND2_X1 _36996_ (
    .A1(_21126_),
    .A2(_02760_),
    .ZN(_02761_)
  );
  INV_X1 _36997_ (
    .A(_02761_),
    .ZN(_02762_)
  );
  AND2_X1 _36998_ (
    .A1(count_instr[41]),
    .A2(count_instr[40]),
    .ZN(_02763_)
  );
  AND2_X1 _36999_ (
    .A1(_02742_),
    .A2(_02763_),
    .ZN(_02764_)
  );
  INV_X1 _37000_ (
    .A(_02764_),
    .ZN(_02765_)
  );
  AND2_X1 _37001_ (
    .A1(resetn),
    .A2(_02765_),
    .ZN(_02766_)
  );
  AND2_X1 _37002_ (
    .A1(_02754_),
    .A2(_02763_),
    .ZN(_02767_)
  );
  AND2_X1 _37003_ (
    .A1(_02762_),
    .A2(_02766_),
    .ZN(_00129_)
  );
  AND2_X1 _37004_ (
    .A1(_21125_),
    .A2(_02765_),
    .ZN(_02768_)
  );
  INV_X1 _37005_ (
    .A(_02768_),
    .ZN(_02769_)
  );
  AND2_X1 _37006_ (
    .A1(resetn),
    .A2(_02769_),
    .ZN(_02770_)
  );
  AND2_X1 _37007_ (
    .A1(count_instr[42]),
    .A2(_02764_),
    .ZN(_02771_)
  );
  INV_X1 _37008_ (
    .A(_02771_),
    .ZN(_02772_)
  );
  AND2_X1 _37009_ (
    .A1(count_instr[42]),
    .A2(_02767_),
    .ZN(_02773_)
  );
  AND2_X1 _37010_ (
    .A1(_02770_),
    .A2(_02772_),
    .ZN(_00130_)
  );
  AND2_X1 _37011_ (
    .A1(_21124_),
    .A2(_02772_),
    .ZN(_02774_)
  );
  INV_X1 _37012_ (
    .A(_02774_),
    .ZN(_02775_)
  );
  AND2_X1 _37013_ (
    .A1(resetn),
    .A2(_02775_),
    .ZN(_02776_)
  );
  AND2_X1 _37014_ (
    .A1(count_instr[43]),
    .A2(_02771_),
    .ZN(_02777_)
  );
  INV_X1 _37015_ (
    .A(_02777_),
    .ZN(_02778_)
  );
  AND2_X1 _37016_ (
    .A1(count_instr[43]),
    .A2(count_instr[42]),
    .ZN(_02779_)
  );
  AND2_X1 _37017_ (
    .A1(count_instr[43]),
    .A2(_02773_),
    .ZN(_02780_)
  );
  AND2_X1 _37018_ (
    .A1(_02776_),
    .A2(_02778_),
    .ZN(_00131_)
  );
  AND2_X1 _37019_ (
    .A1(_21123_),
    .A2(_02778_),
    .ZN(_02781_)
  );
  INV_X1 _37020_ (
    .A(_02781_),
    .ZN(_02782_)
  );
  AND2_X1 _37021_ (
    .A1(resetn),
    .A2(_02782_),
    .ZN(_02783_)
  );
  AND2_X1 _37022_ (
    .A1(count_instr[44]),
    .A2(_02777_),
    .ZN(_02784_)
  );
  INV_X1 _37023_ (
    .A(_02784_),
    .ZN(_02785_)
  );
  AND2_X1 _37024_ (
    .A1(count_instr[44]),
    .A2(_02780_),
    .ZN(_02786_)
  );
  AND2_X1 _37025_ (
    .A1(_02783_),
    .A2(_02785_),
    .ZN(_00132_)
  );
  AND2_X1 _37026_ (
    .A1(_21122_),
    .A2(_02785_),
    .ZN(_02787_)
  );
  INV_X1 _37027_ (
    .A(_02787_),
    .ZN(_02788_)
  );
  AND2_X1 _37028_ (
    .A1(count_instr[45]),
    .A2(count_instr[44]),
    .ZN(_02789_)
  );
  AND2_X1 _37029_ (
    .A1(_02779_),
    .A2(_02789_),
    .ZN(_02790_)
  );
  AND2_X1 _37030_ (
    .A1(_02764_),
    .A2(_02790_),
    .ZN(_02791_)
  );
  INV_X1 _37031_ (
    .A(_02791_),
    .ZN(_02792_)
  );
  AND2_X1 _37032_ (
    .A1(resetn),
    .A2(_02792_),
    .ZN(_02793_)
  );
  AND2_X1 _37033_ (
    .A1(count_instr[45]),
    .A2(_02786_),
    .ZN(_02794_)
  );
  AND2_X1 _37034_ (
    .A1(_02788_),
    .A2(_02793_),
    .ZN(_00133_)
  );
  AND2_X1 _37035_ (
    .A1(_21121_),
    .A2(_02792_),
    .ZN(_02795_)
  );
  INV_X1 _37036_ (
    .A(_02795_),
    .ZN(_02796_)
  );
  AND2_X1 _37037_ (
    .A1(resetn),
    .A2(_02796_),
    .ZN(_02797_)
  );
  AND2_X1 _37038_ (
    .A1(count_instr[46]),
    .A2(_02794_),
    .ZN(_02798_)
  );
  INV_X1 _37039_ (
    .A(_02798_),
    .ZN(_02799_)
  );
  AND2_X1 _37040_ (
    .A1(_02797_),
    .A2(_02799_),
    .ZN(_00134_)
  );
  AND2_X1 _37041_ (
    .A1(_21120_),
    .A2(_02799_),
    .ZN(_02800_)
  );
  INV_X1 _37042_ (
    .A(_02800_),
    .ZN(_02801_)
  );
  AND2_X1 _37043_ (
    .A1(resetn),
    .A2(_02801_),
    .ZN(_02802_)
  );
  AND2_X1 _37044_ (
    .A1(count_instr[47]),
    .A2(_02798_),
    .ZN(_02803_)
  );
  INV_X1 _37045_ (
    .A(_02803_),
    .ZN(_02804_)
  );
  AND2_X1 _37046_ (
    .A1(_02802_),
    .A2(_02804_),
    .ZN(_00135_)
  );
  AND2_X1 _37047_ (
    .A1(count_instr[47]),
    .A2(count_instr[46]),
    .ZN(_02805_)
  );
  AND2_X1 _37048_ (
    .A1(_02763_),
    .A2(_02805_),
    .ZN(_02806_)
  );
  AND2_X1 _37049_ (
    .A1(_02790_),
    .A2(_02806_),
    .ZN(_02807_)
  );
  AND2_X1 _37050_ (
    .A1(_02742_),
    .A2(_02807_),
    .ZN(_02808_)
  );
  AND2_X1 _37051_ (
    .A1(_02746_),
    .A2(_02807_),
    .ZN(_02809_)
  );
  INV_X1 _37052_ (
    .A(_02809_),
    .ZN(_02810_)
  );
  AND2_X1 _37053_ (
    .A1(_21119_),
    .A2(_02810_),
    .ZN(_02811_)
  );
  INV_X1 _37054_ (
    .A(_02811_),
    .ZN(_02812_)
  );
  AND2_X1 _37055_ (
    .A1(resetn),
    .A2(_02812_),
    .ZN(_02813_)
  );
  AND2_X1 _37056_ (
    .A1(count_instr[48]),
    .A2(_02808_),
    .ZN(_02814_)
  );
  INV_X1 _37057_ (
    .A(_02814_),
    .ZN(_02815_)
  );
  AND2_X1 _37058_ (
    .A1(_02813_),
    .A2(_02815_),
    .ZN(_00136_)
  );
  AND2_X1 _37059_ (
    .A1(_21118_),
    .A2(_02815_),
    .ZN(_02816_)
  );
  INV_X1 _37060_ (
    .A(_02816_),
    .ZN(_02817_)
  );
  AND2_X1 _37061_ (
    .A1(resetn),
    .A2(_02817_),
    .ZN(_02818_)
  );
  AND2_X1 _37062_ (
    .A1(count_instr[49]),
    .A2(_02814_),
    .ZN(_02819_)
  );
  INV_X1 _37063_ (
    .A(_02819_),
    .ZN(_02820_)
  );
  AND2_X1 _37064_ (
    .A1(count_instr[49]),
    .A2(count_instr[48]),
    .ZN(_02821_)
  );
  AND2_X1 _37065_ (
    .A1(_02809_),
    .A2(_02821_),
    .ZN(_02822_)
  );
  AND2_X1 _37066_ (
    .A1(_02818_),
    .A2(_02820_),
    .ZN(_00137_)
  );
  AND2_X1 _37067_ (
    .A1(_21117_),
    .A2(_02820_),
    .ZN(_02823_)
  );
  INV_X1 _37068_ (
    .A(_02823_),
    .ZN(_02824_)
  );
  AND2_X1 _37069_ (
    .A1(resetn),
    .A2(_02824_),
    .ZN(_02825_)
  );
  AND2_X1 _37070_ (
    .A1(count_instr[50]),
    .A2(_02822_),
    .ZN(_02826_)
  );
  INV_X1 _37071_ (
    .A(_02826_),
    .ZN(_02827_)
  );
  AND2_X1 _37072_ (
    .A1(_02825_),
    .A2(_02827_),
    .ZN(_00138_)
  );
  AND2_X1 _37073_ (
    .A1(_21116_),
    .A2(_02827_),
    .ZN(_02828_)
  );
  INV_X1 _37074_ (
    .A(_02828_),
    .ZN(_02829_)
  );
  AND2_X1 _37075_ (
    .A1(resetn),
    .A2(_02829_),
    .ZN(_02830_)
  );
  AND2_X1 _37076_ (
    .A1(count_instr[51]),
    .A2(_02826_),
    .ZN(_02831_)
  );
  INV_X1 _37077_ (
    .A(_02831_),
    .ZN(_02832_)
  );
  AND2_X1 _37078_ (
    .A1(_02830_),
    .A2(_02832_),
    .ZN(_00139_)
  );
  AND2_X1 _37079_ (
    .A1(count_instr[51]),
    .A2(_02821_),
    .ZN(_02833_)
  );
  AND2_X1 _37080_ (
    .A1(_21115_),
    .A2(_02832_),
    .ZN(_02834_)
  );
  INV_X1 _37081_ (
    .A(_02834_),
    .ZN(_02835_)
  );
  AND2_X1 _37082_ (
    .A1(resetn),
    .A2(_02835_),
    .ZN(_02836_)
  );
  AND2_X1 _37083_ (
    .A1(count_instr[52]),
    .A2(_02831_),
    .ZN(_02837_)
  );
  INV_X1 _37084_ (
    .A(_02837_),
    .ZN(_02838_)
  );
  AND2_X1 _37085_ (
    .A1(_02836_),
    .A2(_02838_),
    .ZN(_00140_)
  );
  AND2_X1 _37086_ (
    .A1(_21114_),
    .A2(_02838_),
    .ZN(_02839_)
  );
  INV_X1 _37087_ (
    .A(_02839_),
    .ZN(_02840_)
  );
  AND2_X1 _37088_ (
    .A1(count_instr[53]),
    .A2(count_instr[52]),
    .ZN(_02841_)
  );
  AND2_X1 _37089_ (
    .A1(count_instr[50]),
    .A2(_02841_),
    .ZN(_02842_)
  );
  AND2_X1 _37090_ (
    .A1(_02833_),
    .A2(_02842_),
    .ZN(_02843_)
  );
  AND2_X1 _37091_ (
    .A1(_02808_),
    .A2(_02843_),
    .ZN(_02844_)
  );
  AND2_X1 _37092_ (
    .A1(resetn),
    .A2(_02840_),
    .ZN(_02845_)
  );
  AND2_X1 _37093_ (
    .A1(_02809_),
    .A2(_02843_),
    .ZN(_02846_)
  );
  INV_X1 _37094_ (
    .A(_02846_),
    .ZN(_02847_)
  );
  AND2_X1 _37095_ (
    .A1(_02845_),
    .A2(_02847_),
    .ZN(_00141_)
  );
  AND2_X1 _37096_ (
    .A1(_21113_),
    .A2(_02847_),
    .ZN(_02848_)
  );
  INV_X1 _37097_ (
    .A(_02848_),
    .ZN(_02849_)
  );
  AND2_X1 _37098_ (
    .A1(resetn),
    .A2(_02849_),
    .ZN(_02850_)
  );
  AND2_X1 _37099_ (
    .A1(count_instr[54]),
    .A2(_02844_),
    .ZN(_02851_)
  );
  AND2_X1 _37100_ (
    .A1(count_instr[54]),
    .A2(_02846_),
    .ZN(_02852_)
  );
  INV_X1 _37101_ (
    .A(_02852_),
    .ZN(_02853_)
  );
  AND2_X1 _37102_ (
    .A1(_02850_),
    .A2(_02853_),
    .ZN(_00142_)
  );
  AND2_X1 _37103_ (
    .A1(_21112_),
    .A2(_02853_),
    .ZN(_02854_)
  );
  INV_X1 _37104_ (
    .A(_02854_),
    .ZN(_02855_)
  );
  AND2_X1 _37105_ (
    .A1(resetn),
    .A2(_02855_),
    .ZN(_02856_)
  );
  AND2_X1 _37106_ (
    .A1(count_instr[55]),
    .A2(_02851_),
    .ZN(_02857_)
  );
  INV_X1 _37107_ (
    .A(_02857_),
    .ZN(_02858_)
  );
  AND2_X1 _37108_ (
    .A1(_02856_),
    .A2(_02858_),
    .ZN(_00143_)
  );
  AND2_X1 _37109_ (
    .A1(_21111_),
    .A2(_02858_),
    .ZN(_02859_)
  );
  INV_X1 _37110_ (
    .A(_02859_),
    .ZN(_02860_)
  );
  AND2_X1 _37111_ (
    .A1(resetn),
    .A2(_02860_),
    .ZN(_02861_)
  );
  AND2_X1 _37112_ (
    .A1(count_instr[56]),
    .A2(_02857_),
    .ZN(_02862_)
  );
  INV_X1 _37113_ (
    .A(_02862_),
    .ZN(_02863_)
  );
  AND2_X1 _37114_ (
    .A1(_02861_),
    .A2(_02863_),
    .ZN(_00144_)
  );
  AND2_X1 _37115_ (
    .A1(_21110_),
    .A2(_02863_),
    .ZN(_02864_)
  );
  INV_X1 _37116_ (
    .A(_02864_),
    .ZN(_02865_)
  );
  AND2_X1 _37117_ (
    .A1(resetn),
    .A2(_02865_),
    .ZN(_02866_)
  );
  AND2_X1 _37118_ (
    .A1(count_instr[57]),
    .A2(_02862_),
    .ZN(_02867_)
  );
  INV_X1 _37119_ (
    .A(_02867_),
    .ZN(_02868_)
  );
  AND2_X1 _37120_ (
    .A1(_02866_),
    .A2(_02868_),
    .ZN(_00145_)
  );
  AND2_X1 _37121_ (
    .A1(_21109_),
    .A2(_02868_),
    .ZN(_02869_)
  );
  INV_X1 _37122_ (
    .A(_02869_),
    .ZN(_02870_)
  );
  AND2_X1 _37123_ (
    .A1(resetn),
    .A2(_02870_),
    .ZN(_02871_)
  );
  AND2_X1 _37124_ (
    .A1(count_instr[58]),
    .A2(_02867_),
    .ZN(_02872_)
  );
  INV_X1 _37125_ (
    .A(_02872_),
    .ZN(_02873_)
  );
  AND2_X1 _37126_ (
    .A1(_02871_),
    .A2(_02873_),
    .ZN(_00146_)
  );
  AND2_X1 _37127_ (
    .A1(_21108_),
    .A2(_02873_),
    .ZN(_02874_)
  );
  INV_X1 _37128_ (
    .A(_02874_),
    .ZN(_02875_)
  );
  AND2_X1 _37129_ (
    .A1(resetn),
    .A2(_02875_),
    .ZN(_02876_)
  );
  AND2_X1 _37130_ (
    .A1(count_instr[59]),
    .A2(_02872_),
    .ZN(_02877_)
  );
  INV_X1 _37131_ (
    .A(_02877_),
    .ZN(_02878_)
  );
  AND2_X1 _37132_ (
    .A1(_02876_),
    .A2(_02878_),
    .ZN(_00147_)
  );
  AND2_X1 _37133_ (
    .A1(_21107_),
    .A2(_02878_),
    .ZN(_02879_)
  );
  INV_X1 _37134_ (
    .A(_02879_),
    .ZN(_02880_)
  );
  AND2_X1 _37135_ (
    .A1(resetn),
    .A2(_02880_),
    .ZN(_02881_)
  );
  AND2_X1 _37136_ (
    .A1(count_instr[60]),
    .A2(_02877_),
    .ZN(_02882_)
  );
  INV_X1 _37137_ (
    .A(_02882_),
    .ZN(_02883_)
  );
  AND2_X1 _37138_ (
    .A1(_02881_),
    .A2(_02883_),
    .ZN(_00148_)
  );
  AND2_X1 _37139_ (
    .A1(_21106_),
    .A2(_02883_),
    .ZN(_02884_)
  );
  INV_X1 _37140_ (
    .A(_02884_),
    .ZN(_02885_)
  );
  AND2_X1 _37141_ (
    .A1(resetn),
    .A2(_02885_),
    .ZN(_02886_)
  );
  AND2_X1 _37142_ (
    .A1(count_instr[61]),
    .A2(_02882_),
    .ZN(_02887_)
  );
  INV_X1 _37143_ (
    .A(_02887_),
    .ZN(_02888_)
  );
  AND2_X1 _37144_ (
    .A1(_02886_),
    .A2(_02888_),
    .ZN(_00149_)
  );
  AND2_X1 _37145_ (
    .A1(_21105_),
    .A2(_02888_),
    .ZN(_02889_)
  );
  INV_X1 _37146_ (
    .A(_02889_),
    .ZN(_02890_)
  );
  AND2_X1 _37147_ (
    .A1(resetn),
    .A2(_02890_),
    .ZN(_02891_)
  );
  AND2_X1 _37148_ (
    .A1(count_instr[62]),
    .A2(_02887_),
    .ZN(_02892_)
  );
  INV_X1 _37149_ (
    .A(_02892_),
    .ZN(_02893_)
  );
  AND2_X1 _37150_ (
    .A1(_02891_),
    .A2(_02893_),
    .ZN(_00150_)
  );
  AND2_X1 _37151_ (
    .A1(count_instr[63]),
    .A2(_02893_),
    .ZN(_02894_)
  );
  INV_X1 _37152_ (
    .A(_02894_),
    .ZN(_02895_)
  );
  AND2_X1 _37153_ (
    .A1(_21104_),
    .A2(_02892_),
    .ZN(_02896_)
  );
  INV_X1 _37154_ (
    .A(_02896_),
    .ZN(_02897_)
  );
  AND2_X1 _37155_ (
    .A1(_02895_),
    .A2(_02897_),
    .ZN(_02898_)
  );
  INV_X1 _37156_ (
    .A(_02898_),
    .ZN(_02899_)
  );
  AND2_X1 _37157_ (
    .A1(resetn),
    .A2(_02899_),
    .ZN(_00151_)
  );
  AND2_X1 _37158_ (
    .A1(eoi[30]),
    .A2(resetn),
    .ZN(_00152_)
  );
  AND2_X1 _37159_ (
    .A1(decoder_trigger),
    .A2(_00017_),
    .ZN(_02900_)
  );
  INV_X1 _37160_ (
    .A(_02900_),
    .ZN(_02901_)
  );
  AND2_X1 _37161_ (
    .A1(instr_sw),
    .A2(_02901_),
    .ZN(_02902_)
  );
  INV_X1 _37162_ (
    .A(_02902_),
    .ZN(_02903_)
  );
  AND2_X1 _37163_ (
    .A1(_21232_),
    .A2(_22052_),
    .ZN(_02904_)
  );
  AND2_X1 _37164_ (
    .A1(_21234_),
    .A2(_02904_),
    .ZN(_02905_)
  );
  INV_X1 _37165_ (
    .A(_02905_),
    .ZN(_02906_)
  );
  AND2_X1 _37166_ (
    .A1(is_sb_sh_sw),
    .A2(_02900_),
    .ZN(_02907_)
  );
  AND2_X1 _37167_ (
    .A1(_02905_),
    .A2(_02907_),
    .ZN(_02908_)
  );
  INV_X1 _37168_ (
    .A(_02908_),
    .ZN(_02909_)
  );
  AND2_X1 _37169_ (
    .A1(_02903_),
    .A2(_02909_),
    .ZN(_02910_)
  );
  INV_X1 _37170_ (
    .A(_02910_),
    .ZN(_00153_)
  );
  AND2_X1 _37171_ (
    .A1(resetn),
    .A2(_02464_),
    .ZN(_02911_)
  );
  INV_X1 _37172_ (
    .A(_02911_),
    .ZN(_02912_)
  );
  AND2_X1 _37173_ (
    .A1(latched_branch),
    .A2(latched_store),
    .ZN(_02913_)
  );
  INV_X1 _37174_ (
    .A(_02913_),
    .ZN(_02914_)
  );
  AND2_X1 _37175_ (
    .A1(reg_next_pc[1]),
    .A2(_02914_),
    .ZN(_02915_)
  );
  INV_X1 _37176_ (
    .A(_02915_),
    .ZN(_02916_)
  );
  AND2_X1 _37177_ (
    .A1(_21067_),
    .A2(_22112_),
    .ZN(_02917_)
  );
  INV_X1 _37178_ (
    .A(_02917_),
    .ZN(_02918_)
  );
  AND2_X1 _37179_ (
    .A1(latched_stalu),
    .A2(_22113_),
    .ZN(_02919_)
  );
  INV_X1 _37180_ (
    .A(_02919_),
    .ZN(_02920_)
  );
  AND2_X1 _37181_ (
    .A1(_02918_),
    .A2(_02920_),
    .ZN(_02921_)
  );
  AND2_X1 _37182_ (
    .A1(_02913_),
    .A2(_02921_),
    .ZN(_02922_)
  );
  INV_X1 _37183_ (
    .A(_02922_),
    .ZN(_02923_)
  );
  AND2_X1 _37184_ (
    .A1(_02916_),
    .A2(_02923_),
    .ZN(_02924_)
  );
  INV_X1 _37185_ (
    .A(_02924_),
    .ZN(_02925_)
  );
  AND2_X1 _37186_ (
    .A1(_02911_),
    .A2(_02925_),
    .ZN(_02926_)
  );
  INV_X1 _37187_ (
    .A(_02926_),
    .ZN(_02927_)
  );
  AND2_X1 _37188_ (
    .A1(resetn),
    .A2(_02465_),
    .ZN(_02928_)
  );
  AND2_X1 _37189_ (
    .A1(reg_pc[1]),
    .A2(_02928_),
    .ZN(_02929_)
  );
  INV_X1 _37190_ (
    .A(_02929_),
    .ZN(_02930_)
  );
  AND2_X1 _37191_ (
    .A1(_02927_),
    .A2(_02930_),
    .ZN(_02931_)
  );
  INV_X1 _37192_ (
    .A(_02931_),
    .ZN(_00154_)
  );
  AND2_X1 _37193_ (
    .A1(reg_next_pc[2]),
    .A2(_02914_),
    .ZN(_02932_)
  );
  INV_X1 _37194_ (
    .A(_02932_),
    .ZN(_02933_)
  );
  AND2_X1 _37195_ (
    .A1(_21067_),
    .A2(_22079_),
    .ZN(_02934_)
  );
  INV_X1 _37196_ (
    .A(_02934_),
    .ZN(_02935_)
  );
  AND2_X1 _37197_ (
    .A1(latched_stalu),
    .A2(_22114_),
    .ZN(_02936_)
  );
  INV_X1 _37198_ (
    .A(_02936_),
    .ZN(_02937_)
  );
  AND2_X1 _37199_ (
    .A1(_02935_),
    .A2(_02937_),
    .ZN(_02938_)
  );
  AND2_X1 _37200_ (
    .A1(_02913_),
    .A2(_02938_),
    .ZN(_02939_)
  );
  INV_X1 _37201_ (
    .A(_02939_),
    .ZN(_02940_)
  );
  AND2_X1 _37202_ (
    .A1(_02933_),
    .A2(_02940_),
    .ZN(_02941_)
  );
  INV_X1 _37203_ (
    .A(_02941_),
    .ZN(_02942_)
  );
  AND2_X1 _37204_ (
    .A1(_02911_),
    .A2(_02942_),
    .ZN(_02943_)
  );
  INV_X1 _37205_ (
    .A(_02943_),
    .ZN(_02944_)
  );
  AND2_X1 _37206_ (
    .A1(reg_pc[2]),
    .A2(_02928_),
    .ZN(_02945_)
  );
  INV_X1 _37207_ (
    .A(_02945_),
    .ZN(_02946_)
  );
  AND2_X1 _37208_ (
    .A1(_02944_),
    .A2(_02946_),
    .ZN(_02947_)
  );
  INV_X1 _37209_ (
    .A(_02947_),
    .ZN(_00155_)
  );
  AND2_X1 _37210_ (
    .A1(reg_next_pc[3]),
    .A2(_02914_),
    .ZN(_02948_)
  );
  INV_X1 _37211_ (
    .A(_02948_),
    .ZN(_02949_)
  );
  AND2_X1 _37212_ (
    .A1(_21067_),
    .A2(_22080_),
    .ZN(_02950_)
  );
  INV_X1 _37213_ (
    .A(_02950_),
    .ZN(_02951_)
  );
  AND2_X1 _37214_ (
    .A1(latched_stalu),
    .A2(_22115_),
    .ZN(_02952_)
  );
  INV_X1 _37215_ (
    .A(_02952_),
    .ZN(_02953_)
  );
  AND2_X1 _37216_ (
    .A1(_02951_),
    .A2(_02953_),
    .ZN(_02954_)
  );
  AND2_X1 _37217_ (
    .A1(_02913_),
    .A2(_02954_),
    .ZN(_02955_)
  );
  INV_X1 _37218_ (
    .A(_02955_),
    .ZN(_02956_)
  );
  AND2_X1 _37219_ (
    .A1(_02949_),
    .A2(_02956_),
    .ZN(_02957_)
  );
  INV_X1 _37220_ (
    .A(_02957_),
    .ZN(_02958_)
  );
  AND2_X1 _37221_ (
    .A1(_02911_),
    .A2(_02958_),
    .ZN(_02959_)
  );
  INV_X1 _37222_ (
    .A(_02959_),
    .ZN(_02960_)
  );
  AND2_X1 _37223_ (
    .A1(reg_pc[3]),
    .A2(_02928_),
    .ZN(_02961_)
  );
  INV_X1 _37224_ (
    .A(_02961_),
    .ZN(_02962_)
  );
  AND2_X1 _37225_ (
    .A1(_02960_),
    .A2(_02962_),
    .ZN(_02963_)
  );
  INV_X1 _37226_ (
    .A(_02963_),
    .ZN(_00156_)
  );
  AND2_X1 _37227_ (
    .A1(reg_next_pc[4]),
    .A2(_02914_),
    .ZN(_02964_)
  );
  INV_X1 _37228_ (
    .A(_02964_),
    .ZN(_02965_)
  );
  AND2_X1 _37229_ (
    .A1(_21067_),
    .A2(_22081_),
    .ZN(_02966_)
  );
  INV_X1 _37230_ (
    .A(_02966_),
    .ZN(_02967_)
  );
  AND2_X1 _37231_ (
    .A1(latched_stalu),
    .A2(_22116_),
    .ZN(_02968_)
  );
  INV_X1 _37232_ (
    .A(_02968_),
    .ZN(_02969_)
  );
  AND2_X1 _37233_ (
    .A1(_02967_),
    .A2(_02969_),
    .ZN(_02970_)
  );
  AND2_X1 _37234_ (
    .A1(_02913_),
    .A2(_02970_),
    .ZN(_02971_)
  );
  INV_X1 _37235_ (
    .A(_02971_),
    .ZN(_02972_)
  );
  AND2_X1 _37236_ (
    .A1(_02965_),
    .A2(_02972_),
    .ZN(_02973_)
  );
  INV_X1 _37237_ (
    .A(_02973_),
    .ZN(_02974_)
  );
  AND2_X1 _37238_ (
    .A1(_02911_),
    .A2(_02974_),
    .ZN(_02975_)
  );
  INV_X1 _37239_ (
    .A(_02975_),
    .ZN(_02976_)
  );
  AND2_X1 _37240_ (
    .A1(reg_pc[4]),
    .A2(_02928_),
    .ZN(_02977_)
  );
  INV_X1 _37241_ (
    .A(_02977_),
    .ZN(_02978_)
  );
  AND2_X1 _37242_ (
    .A1(_02976_),
    .A2(_02978_),
    .ZN(_02979_)
  );
  INV_X1 _37243_ (
    .A(_02979_),
    .ZN(_00157_)
  );
  AND2_X1 _37244_ (
    .A1(reg_next_pc[5]),
    .A2(_02914_),
    .ZN(_02980_)
  );
  INV_X1 _37245_ (
    .A(_02980_),
    .ZN(_02981_)
  );
  AND2_X1 _37246_ (
    .A1(_21067_),
    .A2(_22082_),
    .ZN(_02982_)
  );
  INV_X1 _37247_ (
    .A(_02982_),
    .ZN(_02983_)
  );
  AND2_X1 _37248_ (
    .A1(latched_stalu),
    .A2(_22117_),
    .ZN(_02984_)
  );
  INV_X1 _37249_ (
    .A(_02984_),
    .ZN(_02985_)
  );
  AND2_X1 _37250_ (
    .A1(_02983_),
    .A2(_02985_),
    .ZN(_02986_)
  );
  AND2_X1 _37251_ (
    .A1(_02913_),
    .A2(_02986_),
    .ZN(_02987_)
  );
  INV_X1 _37252_ (
    .A(_02987_),
    .ZN(_02988_)
  );
  AND2_X1 _37253_ (
    .A1(_02981_),
    .A2(_02988_),
    .ZN(_02989_)
  );
  INV_X1 _37254_ (
    .A(_02989_),
    .ZN(_02990_)
  );
  AND2_X1 _37255_ (
    .A1(_02911_),
    .A2(_02990_),
    .ZN(_02991_)
  );
  INV_X1 _37256_ (
    .A(_02991_),
    .ZN(_02992_)
  );
  AND2_X1 _37257_ (
    .A1(reg_pc[5]),
    .A2(_02928_),
    .ZN(_02993_)
  );
  INV_X1 _37258_ (
    .A(_02993_),
    .ZN(_02994_)
  );
  AND2_X1 _37259_ (
    .A1(_02992_),
    .A2(_02994_),
    .ZN(_02995_)
  );
  INV_X1 _37260_ (
    .A(_02995_),
    .ZN(_00158_)
  );
  AND2_X1 _37261_ (
    .A1(reg_next_pc[6]),
    .A2(_02914_),
    .ZN(_02996_)
  );
  INV_X1 _37262_ (
    .A(_02996_),
    .ZN(_02997_)
  );
  AND2_X1 _37263_ (
    .A1(_21067_),
    .A2(_22083_),
    .ZN(_02998_)
  );
  INV_X1 _37264_ (
    .A(_02998_),
    .ZN(_02999_)
  );
  AND2_X1 _37265_ (
    .A1(latched_stalu),
    .A2(_22118_),
    .ZN(_03000_)
  );
  INV_X1 _37266_ (
    .A(_03000_),
    .ZN(_03001_)
  );
  AND2_X1 _37267_ (
    .A1(_02999_),
    .A2(_03001_),
    .ZN(_03002_)
  );
  AND2_X1 _37268_ (
    .A1(_02913_),
    .A2(_03002_),
    .ZN(_03003_)
  );
  INV_X1 _37269_ (
    .A(_03003_),
    .ZN(_03004_)
  );
  AND2_X1 _37270_ (
    .A1(_02997_),
    .A2(_03004_),
    .ZN(_03005_)
  );
  INV_X1 _37271_ (
    .A(_03005_),
    .ZN(_03006_)
  );
  AND2_X1 _37272_ (
    .A1(_02911_),
    .A2(_03006_),
    .ZN(_03007_)
  );
  INV_X1 _37273_ (
    .A(_03007_),
    .ZN(_03008_)
  );
  AND2_X1 _37274_ (
    .A1(reg_pc[6]),
    .A2(_02928_),
    .ZN(_03009_)
  );
  INV_X1 _37275_ (
    .A(_03009_),
    .ZN(_03010_)
  );
  AND2_X1 _37276_ (
    .A1(_03008_),
    .A2(_03010_),
    .ZN(_03011_)
  );
  INV_X1 _37277_ (
    .A(_03011_),
    .ZN(_00159_)
  );
  AND2_X1 _37278_ (
    .A1(reg_next_pc[7]),
    .A2(_02914_),
    .ZN(_03012_)
  );
  INV_X1 _37279_ (
    .A(_03012_),
    .ZN(_03013_)
  );
  AND2_X1 _37280_ (
    .A1(_21067_),
    .A2(_22084_),
    .ZN(_03014_)
  );
  INV_X1 _37281_ (
    .A(_03014_),
    .ZN(_03015_)
  );
  AND2_X1 _37282_ (
    .A1(latched_stalu),
    .A2(_22119_),
    .ZN(_03016_)
  );
  INV_X1 _37283_ (
    .A(_03016_),
    .ZN(_03017_)
  );
  AND2_X1 _37284_ (
    .A1(_03015_),
    .A2(_03017_),
    .ZN(_03018_)
  );
  AND2_X1 _37285_ (
    .A1(_02913_),
    .A2(_03018_),
    .ZN(_03019_)
  );
  INV_X1 _37286_ (
    .A(_03019_),
    .ZN(_03020_)
  );
  AND2_X1 _37287_ (
    .A1(_03013_),
    .A2(_03020_),
    .ZN(_03021_)
  );
  INV_X1 _37288_ (
    .A(_03021_),
    .ZN(_03022_)
  );
  AND2_X1 _37289_ (
    .A1(_02911_),
    .A2(_03022_),
    .ZN(_03023_)
  );
  INV_X1 _37290_ (
    .A(_03023_),
    .ZN(_03024_)
  );
  AND2_X1 _37291_ (
    .A1(reg_pc[7]),
    .A2(_02928_),
    .ZN(_03025_)
  );
  INV_X1 _37292_ (
    .A(_03025_),
    .ZN(_03026_)
  );
  AND2_X1 _37293_ (
    .A1(_03024_),
    .A2(_03026_),
    .ZN(_03027_)
  );
  INV_X1 _37294_ (
    .A(_03027_),
    .ZN(_00160_)
  );
  AND2_X1 _37295_ (
    .A1(reg_next_pc[8]),
    .A2(_02914_),
    .ZN(_03028_)
  );
  INV_X1 _37296_ (
    .A(_03028_),
    .ZN(_03029_)
  );
  AND2_X1 _37297_ (
    .A1(_21067_),
    .A2(_22085_),
    .ZN(_03030_)
  );
  INV_X1 _37298_ (
    .A(_03030_),
    .ZN(_03031_)
  );
  AND2_X1 _37299_ (
    .A1(latched_stalu),
    .A2(_22120_),
    .ZN(_03032_)
  );
  INV_X1 _37300_ (
    .A(_03032_),
    .ZN(_03033_)
  );
  AND2_X1 _37301_ (
    .A1(_03031_),
    .A2(_03033_),
    .ZN(_03034_)
  );
  AND2_X1 _37302_ (
    .A1(_02913_),
    .A2(_03034_),
    .ZN(_03035_)
  );
  INV_X1 _37303_ (
    .A(_03035_),
    .ZN(_03036_)
  );
  AND2_X1 _37304_ (
    .A1(_03029_),
    .A2(_03036_),
    .ZN(_03037_)
  );
  INV_X1 _37305_ (
    .A(_03037_),
    .ZN(_03038_)
  );
  AND2_X1 _37306_ (
    .A1(_02911_),
    .A2(_03038_),
    .ZN(_03039_)
  );
  INV_X1 _37307_ (
    .A(_03039_),
    .ZN(_03040_)
  );
  AND2_X1 _37308_ (
    .A1(reg_pc[8]),
    .A2(_02928_),
    .ZN(_03041_)
  );
  INV_X1 _37309_ (
    .A(_03041_),
    .ZN(_03042_)
  );
  AND2_X1 _37310_ (
    .A1(_03040_),
    .A2(_03042_),
    .ZN(_03043_)
  );
  INV_X1 _37311_ (
    .A(_03043_),
    .ZN(_00161_)
  );
  AND2_X1 _37312_ (
    .A1(reg_next_pc[9]),
    .A2(_02914_),
    .ZN(_03044_)
  );
  INV_X1 _37313_ (
    .A(_03044_),
    .ZN(_03045_)
  );
  AND2_X1 _37314_ (
    .A1(_21067_),
    .A2(_22086_),
    .ZN(_03046_)
  );
  INV_X1 _37315_ (
    .A(_03046_),
    .ZN(_03047_)
  );
  AND2_X1 _37316_ (
    .A1(latched_stalu),
    .A2(_22121_),
    .ZN(_03048_)
  );
  INV_X1 _37317_ (
    .A(_03048_),
    .ZN(_03049_)
  );
  AND2_X1 _37318_ (
    .A1(_03047_),
    .A2(_03049_),
    .ZN(_03050_)
  );
  AND2_X1 _37319_ (
    .A1(_02913_),
    .A2(_03050_),
    .ZN(_03051_)
  );
  INV_X1 _37320_ (
    .A(_03051_),
    .ZN(_03052_)
  );
  AND2_X1 _37321_ (
    .A1(_03045_),
    .A2(_03052_),
    .ZN(_03053_)
  );
  INV_X1 _37322_ (
    .A(_03053_),
    .ZN(_03054_)
  );
  AND2_X1 _37323_ (
    .A1(_02911_),
    .A2(_03054_),
    .ZN(_03055_)
  );
  INV_X1 _37324_ (
    .A(_03055_),
    .ZN(_03056_)
  );
  AND2_X1 _37325_ (
    .A1(reg_pc[9]),
    .A2(_02928_),
    .ZN(_03057_)
  );
  INV_X1 _37326_ (
    .A(_03057_),
    .ZN(_03058_)
  );
  AND2_X1 _37327_ (
    .A1(_03056_),
    .A2(_03058_),
    .ZN(_03059_)
  );
  INV_X1 _37328_ (
    .A(_03059_),
    .ZN(_00162_)
  );
  AND2_X1 _37329_ (
    .A1(reg_next_pc[10]),
    .A2(_02914_),
    .ZN(_03060_)
  );
  INV_X1 _37330_ (
    .A(_03060_),
    .ZN(_03061_)
  );
  AND2_X1 _37331_ (
    .A1(_21067_),
    .A2(_22087_),
    .ZN(_03062_)
  );
  INV_X1 _37332_ (
    .A(_03062_),
    .ZN(_03063_)
  );
  AND2_X1 _37333_ (
    .A1(latched_stalu),
    .A2(_22122_),
    .ZN(_03064_)
  );
  INV_X1 _37334_ (
    .A(_03064_),
    .ZN(_03065_)
  );
  AND2_X1 _37335_ (
    .A1(_03063_),
    .A2(_03065_),
    .ZN(_03066_)
  );
  AND2_X1 _37336_ (
    .A1(_02913_),
    .A2(_03066_),
    .ZN(_03067_)
  );
  INV_X1 _37337_ (
    .A(_03067_),
    .ZN(_03068_)
  );
  AND2_X1 _37338_ (
    .A1(_03061_),
    .A2(_03068_),
    .ZN(_03069_)
  );
  INV_X1 _37339_ (
    .A(_03069_),
    .ZN(_03070_)
  );
  AND2_X1 _37340_ (
    .A1(_02911_),
    .A2(_03070_),
    .ZN(_03071_)
  );
  INV_X1 _37341_ (
    .A(_03071_),
    .ZN(_03072_)
  );
  AND2_X1 _37342_ (
    .A1(reg_pc[10]),
    .A2(_02928_),
    .ZN(_03073_)
  );
  INV_X1 _37343_ (
    .A(_03073_),
    .ZN(_03074_)
  );
  AND2_X1 _37344_ (
    .A1(_03072_),
    .A2(_03074_),
    .ZN(_03075_)
  );
  INV_X1 _37345_ (
    .A(_03075_),
    .ZN(_00163_)
  );
  AND2_X1 _37346_ (
    .A1(reg_next_pc[11]),
    .A2(_02914_),
    .ZN(_03076_)
  );
  INV_X1 _37347_ (
    .A(_03076_),
    .ZN(_03077_)
  );
  AND2_X1 _37348_ (
    .A1(_21067_),
    .A2(_22088_),
    .ZN(_03078_)
  );
  INV_X1 _37349_ (
    .A(_03078_),
    .ZN(_03079_)
  );
  AND2_X1 _37350_ (
    .A1(latched_stalu),
    .A2(_22123_),
    .ZN(_03080_)
  );
  INV_X1 _37351_ (
    .A(_03080_),
    .ZN(_03081_)
  );
  AND2_X1 _37352_ (
    .A1(_03079_),
    .A2(_03081_),
    .ZN(_03082_)
  );
  AND2_X1 _37353_ (
    .A1(_02913_),
    .A2(_03082_),
    .ZN(_03083_)
  );
  INV_X1 _37354_ (
    .A(_03083_),
    .ZN(_03084_)
  );
  AND2_X1 _37355_ (
    .A1(_03077_),
    .A2(_03084_),
    .ZN(_03085_)
  );
  INV_X1 _37356_ (
    .A(_03085_),
    .ZN(_03086_)
  );
  AND2_X1 _37357_ (
    .A1(_02911_),
    .A2(_03086_),
    .ZN(_03087_)
  );
  INV_X1 _37358_ (
    .A(_03087_),
    .ZN(_03088_)
  );
  AND2_X1 _37359_ (
    .A1(reg_pc[11]),
    .A2(_02928_),
    .ZN(_03089_)
  );
  INV_X1 _37360_ (
    .A(_03089_),
    .ZN(_03090_)
  );
  AND2_X1 _37361_ (
    .A1(_03088_),
    .A2(_03090_),
    .ZN(_03091_)
  );
  INV_X1 _37362_ (
    .A(_03091_),
    .ZN(_00164_)
  );
  AND2_X1 _37363_ (
    .A1(reg_next_pc[12]),
    .A2(_02914_),
    .ZN(_03092_)
  );
  INV_X1 _37364_ (
    .A(_03092_),
    .ZN(_03093_)
  );
  AND2_X1 _37365_ (
    .A1(_21067_),
    .A2(_22089_),
    .ZN(_03094_)
  );
  INV_X1 _37366_ (
    .A(_03094_),
    .ZN(_03095_)
  );
  AND2_X1 _37367_ (
    .A1(latched_stalu),
    .A2(_22124_),
    .ZN(_03096_)
  );
  INV_X1 _37368_ (
    .A(_03096_),
    .ZN(_03097_)
  );
  AND2_X1 _37369_ (
    .A1(_03095_),
    .A2(_03097_),
    .ZN(_03098_)
  );
  AND2_X1 _37370_ (
    .A1(_02913_),
    .A2(_03098_),
    .ZN(_03099_)
  );
  INV_X1 _37371_ (
    .A(_03099_),
    .ZN(_03100_)
  );
  AND2_X1 _37372_ (
    .A1(_03093_),
    .A2(_03100_),
    .ZN(_03101_)
  );
  INV_X1 _37373_ (
    .A(_03101_),
    .ZN(_03102_)
  );
  AND2_X1 _37374_ (
    .A1(_02911_),
    .A2(_03102_),
    .ZN(_03103_)
  );
  INV_X1 _37375_ (
    .A(_03103_),
    .ZN(_03104_)
  );
  AND2_X1 _37376_ (
    .A1(reg_pc[12]),
    .A2(_02928_),
    .ZN(_03105_)
  );
  INV_X1 _37377_ (
    .A(_03105_),
    .ZN(_03106_)
  );
  AND2_X1 _37378_ (
    .A1(_03104_),
    .A2(_03106_),
    .ZN(_03107_)
  );
  INV_X1 _37379_ (
    .A(_03107_),
    .ZN(_00165_)
  );
  AND2_X1 _37380_ (
    .A1(reg_next_pc[13]),
    .A2(_02914_),
    .ZN(_03108_)
  );
  INV_X1 _37381_ (
    .A(_03108_),
    .ZN(_03109_)
  );
  AND2_X1 _37382_ (
    .A1(_21067_),
    .A2(_22090_),
    .ZN(_03110_)
  );
  INV_X1 _37383_ (
    .A(_03110_),
    .ZN(_03111_)
  );
  AND2_X1 _37384_ (
    .A1(latched_stalu),
    .A2(_22125_),
    .ZN(_03112_)
  );
  INV_X1 _37385_ (
    .A(_03112_),
    .ZN(_03113_)
  );
  AND2_X1 _37386_ (
    .A1(_03111_),
    .A2(_03113_),
    .ZN(_03114_)
  );
  AND2_X1 _37387_ (
    .A1(_02913_),
    .A2(_03114_),
    .ZN(_03115_)
  );
  INV_X1 _37388_ (
    .A(_03115_),
    .ZN(_03116_)
  );
  AND2_X1 _37389_ (
    .A1(_03109_),
    .A2(_03116_),
    .ZN(_03117_)
  );
  INV_X1 _37390_ (
    .A(_03117_),
    .ZN(_03118_)
  );
  AND2_X1 _37391_ (
    .A1(_02911_),
    .A2(_03118_),
    .ZN(_03119_)
  );
  INV_X1 _37392_ (
    .A(_03119_),
    .ZN(_03120_)
  );
  AND2_X1 _37393_ (
    .A1(reg_pc[13]),
    .A2(_02928_),
    .ZN(_03121_)
  );
  INV_X1 _37394_ (
    .A(_03121_),
    .ZN(_03122_)
  );
  AND2_X1 _37395_ (
    .A1(_03120_),
    .A2(_03122_),
    .ZN(_03123_)
  );
  INV_X1 _37396_ (
    .A(_03123_),
    .ZN(_00166_)
  );
  AND2_X1 _37397_ (
    .A1(reg_next_pc[14]),
    .A2(_02914_),
    .ZN(_03124_)
  );
  INV_X1 _37398_ (
    .A(_03124_),
    .ZN(_03125_)
  );
  AND2_X1 _37399_ (
    .A1(_21067_),
    .A2(_22091_),
    .ZN(_03126_)
  );
  INV_X1 _37400_ (
    .A(_03126_),
    .ZN(_03127_)
  );
  AND2_X1 _37401_ (
    .A1(latched_stalu),
    .A2(_22126_),
    .ZN(_03128_)
  );
  INV_X1 _37402_ (
    .A(_03128_),
    .ZN(_03129_)
  );
  AND2_X1 _37403_ (
    .A1(_03127_),
    .A2(_03129_),
    .ZN(_03130_)
  );
  AND2_X1 _37404_ (
    .A1(_02913_),
    .A2(_03130_),
    .ZN(_03131_)
  );
  INV_X1 _37405_ (
    .A(_03131_),
    .ZN(_03132_)
  );
  AND2_X1 _37406_ (
    .A1(_03125_),
    .A2(_03132_),
    .ZN(_03133_)
  );
  INV_X1 _37407_ (
    .A(_03133_),
    .ZN(_03134_)
  );
  AND2_X1 _37408_ (
    .A1(_02911_),
    .A2(_03134_),
    .ZN(_03135_)
  );
  INV_X1 _37409_ (
    .A(_03135_),
    .ZN(_03136_)
  );
  AND2_X1 _37410_ (
    .A1(reg_pc[14]),
    .A2(_02928_),
    .ZN(_03137_)
  );
  INV_X1 _37411_ (
    .A(_03137_),
    .ZN(_03138_)
  );
  AND2_X1 _37412_ (
    .A1(_03136_),
    .A2(_03138_),
    .ZN(_03139_)
  );
  INV_X1 _37413_ (
    .A(_03139_),
    .ZN(_00167_)
  );
  AND2_X1 _37414_ (
    .A1(reg_next_pc[15]),
    .A2(_02914_),
    .ZN(_03140_)
  );
  INV_X1 _37415_ (
    .A(_03140_),
    .ZN(_03141_)
  );
  AND2_X1 _37416_ (
    .A1(_21067_),
    .A2(_22092_),
    .ZN(_03142_)
  );
  INV_X1 _37417_ (
    .A(_03142_),
    .ZN(_03143_)
  );
  AND2_X1 _37418_ (
    .A1(latched_stalu),
    .A2(_22127_),
    .ZN(_03144_)
  );
  INV_X1 _37419_ (
    .A(_03144_),
    .ZN(_03145_)
  );
  AND2_X1 _37420_ (
    .A1(_03143_),
    .A2(_03145_),
    .ZN(_03146_)
  );
  AND2_X1 _37421_ (
    .A1(_02913_),
    .A2(_03146_),
    .ZN(_03147_)
  );
  INV_X1 _37422_ (
    .A(_03147_),
    .ZN(_03148_)
  );
  AND2_X1 _37423_ (
    .A1(_03141_),
    .A2(_03148_),
    .ZN(_03149_)
  );
  INV_X1 _37424_ (
    .A(_03149_),
    .ZN(_03150_)
  );
  AND2_X1 _37425_ (
    .A1(_02911_),
    .A2(_03150_),
    .ZN(_03151_)
  );
  INV_X1 _37426_ (
    .A(_03151_),
    .ZN(_03152_)
  );
  AND2_X1 _37427_ (
    .A1(reg_pc[15]),
    .A2(_02928_),
    .ZN(_03153_)
  );
  INV_X1 _37428_ (
    .A(_03153_),
    .ZN(_03154_)
  );
  AND2_X1 _37429_ (
    .A1(_03152_),
    .A2(_03154_),
    .ZN(_03155_)
  );
  INV_X1 _37430_ (
    .A(_03155_),
    .ZN(_00168_)
  );
  AND2_X1 _37431_ (
    .A1(reg_next_pc[16]),
    .A2(_02914_),
    .ZN(_03156_)
  );
  INV_X1 _37432_ (
    .A(_03156_),
    .ZN(_03157_)
  );
  AND2_X1 _37433_ (
    .A1(_21067_),
    .A2(_22093_),
    .ZN(_03158_)
  );
  INV_X1 _37434_ (
    .A(_03158_),
    .ZN(_03159_)
  );
  AND2_X1 _37435_ (
    .A1(latched_stalu),
    .A2(_22128_),
    .ZN(_03160_)
  );
  INV_X1 _37436_ (
    .A(_03160_),
    .ZN(_03161_)
  );
  AND2_X1 _37437_ (
    .A1(_03159_),
    .A2(_03161_),
    .ZN(_03162_)
  );
  AND2_X1 _37438_ (
    .A1(_02913_),
    .A2(_03162_),
    .ZN(_03163_)
  );
  INV_X1 _37439_ (
    .A(_03163_),
    .ZN(_03164_)
  );
  AND2_X1 _37440_ (
    .A1(_03157_),
    .A2(_03164_),
    .ZN(_03165_)
  );
  INV_X1 _37441_ (
    .A(_03165_),
    .ZN(_03166_)
  );
  AND2_X1 _37442_ (
    .A1(_02911_),
    .A2(_03166_),
    .ZN(_03167_)
  );
  INV_X1 _37443_ (
    .A(_03167_),
    .ZN(_03168_)
  );
  AND2_X1 _37444_ (
    .A1(reg_pc[16]),
    .A2(_02928_),
    .ZN(_03169_)
  );
  INV_X1 _37445_ (
    .A(_03169_),
    .ZN(_03170_)
  );
  AND2_X1 _37446_ (
    .A1(_03168_),
    .A2(_03170_),
    .ZN(_03171_)
  );
  INV_X1 _37447_ (
    .A(_03171_),
    .ZN(_00169_)
  );
  AND2_X1 _37448_ (
    .A1(reg_next_pc[17]),
    .A2(_02914_),
    .ZN(_03172_)
  );
  INV_X1 _37449_ (
    .A(_03172_),
    .ZN(_03173_)
  );
  AND2_X1 _37450_ (
    .A1(_21067_),
    .A2(_22094_),
    .ZN(_03174_)
  );
  INV_X1 _37451_ (
    .A(_03174_),
    .ZN(_03175_)
  );
  AND2_X1 _37452_ (
    .A1(latched_stalu),
    .A2(_22129_),
    .ZN(_03176_)
  );
  INV_X1 _37453_ (
    .A(_03176_),
    .ZN(_03177_)
  );
  AND2_X1 _37454_ (
    .A1(_03175_),
    .A2(_03177_),
    .ZN(_03178_)
  );
  AND2_X1 _37455_ (
    .A1(_02913_),
    .A2(_03178_),
    .ZN(_03179_)
  );
  INV_X1 _37456_ (
    .A(_03179_),
    .ZN(_03180_)
  );
  AND2_X1 _37457_ (
    .A1(_03173_),
    .A2(_03180_),
    .ZN(_03181_)
  );
  INV_X1 _37458_ (
    .A(_03181_),
    .ZN(_03182_)
  );
  AND2_X1 _37459_ (
    .A1(_02911_),
    .A2(_03182_),
    .ZN(_03183_)
  );
  INV_X1 _37460_ (
    .A(_03183_),
    .ZN(_03184_)
  );
  AND2_X1 _37461_ (
    .A1(reg_pc[17]),
    .A2(_02928_),
    .ZN(_03185_)
  );
  INV_X1 _37462_ (
    .A(_03185_),
    .ZN(_03186_)
  );
  AND2_X1 _37463_ (
    .A1(_03184_),
    .A2(_03186_),
    .ZN(_03187_)
  );
  INV_X1 _37464_ (
    .A(_03187_),
    .ZN(_00170_)
  );
  AND2_X1 _37465_ (
    .A1(reg_next_pc[18]),
    .A2(_02914_),
    .ZN(_03188_)
  );
  INV_X1 _37466_ (
    .A(_03188_),
    .ZN(_03189_)
  );
  AND2_X1 _37467_ (
    .A1(_21067_),
    .A2(_22095_),
    .ZN(_03190_)
  );
  INV_X1 _37468_ (
    .A(_03190_),
    .ZN(_03191_)
  );
  AND2_X1 _37469_ (
    .A1(latched_stalu),
    .A2(_22130_),
    .ZN(_03192_)
  );
  INV_X1 _37470_ (
    .A(_03192_),
    .ZN(_03193_)
  );
  AND2_X1 _37471_ (
    .A1(_03191_),
    .A2(_03193_),
    .ZN(_03194_)
  );
  AND2_X1 _37472_ (
    .A1(_02913_),
    .A2(_03194_),
    .ZN(_03195_)
  );
  INV_X1 _37473_ (
    .A(_03195_),
    .ZN(_03196_)
  );
  AND2_X1 _37474_ (
    .A1(_03189_),
    .A2(_03196_),
    .ZN(_03197_)
  );
  INV_X1 _37475_ (
    .A(_03197_),
    .ZN(_03198_)
  );
  AND2_X1 _37476_ (
    .A1(_02911_),
    .A2(_03198_),
    .ZN(_03199_)
  );
  INV_X1 _37477_ (
    .A(_03199_),
    .ZN(_03200_)
  );
  AND2_X1 _37478_ (
    .A1(reg_pc[18]),
    .A2(_02928_),
    .ZN(_03201_)
  );
  INV_X1 _37479_ (
    .A(_03201_),
    .ZN(_03202_)
  );
  AND2_X1 _37480_ (
    .A1(_03200_),
    .A2(_03202_),
    .ZN(_03203_)
  );
  INV_X1 _37481_ (
    .A(_03203_),
    .ZN(_00171_)
  );
  AND2_X1 _37482_ (
    .A1(reg_next_pc[19]),
    .A2(_02914_),
    .ZN(_03204_)
  );
  INV_X1 _37483_ (
    .A(_03204_),
    .ZN(_03205_)
  );
  AND2_X1 _37484_ (
    .A1(_21067_),
    .A2(_22096_),
    .ZN(_03206_)
  );
  INV_X1 _37485_ (
    .A(_03206_),
    .ZN(_03207_)
  );
  AND2_X1 _37486_ (
    .A1(latched_stalu),
    .A2(_22131_),
    .ZN(_03208_)
  );
  INV_X1 _37487_ (
    .A(_03208_),
    .ZN(_03209_)
  );
  AND2_X1 _37488_ (
    .A1(_03207_),
    .A2(_03209_),
    .ZN(_03210_)
  );
  AND2_X1 _37489_ (
    .A1(_02913_),
    .A2(_03210_),
    .ZN(_03211_)
  );
  INV_X1 _37490_ (
    .A(_03211_),
    .ZN(_03212_)
  );
  AND2_X1 _37491_ (
    .A1(_03205_),
    .A2(_03212_),
    .ZN(_03213_)
  );
  INV_X1 _37492_ (
    .A(_03213_),
    .ZN(_03214_)
  );
  AND2_X1 _37493_ (
    .A1(_02911_),
    .A2(_03214_),
    .ZN(_03215_)
  );
  INV_X1 _37494_ (
    .A(_03215_),
    .ZN(_03216_)
  );
  AND2_X1 _37495_ (
    .A1(reg_pc[19]),
    .A2(_02928_),
    .ZN(_03217_)
  );
  INV_X1 _37496_ (
    .A(_03217_),
    .ZN(_03218_)
  );
  AND2_X1 _37497_ (
    .A1(_03216_),
    .A2(_03218_),
    .ZN(_03219_)
  );
  INV_X1 _37498_ (
    .A(_03219_),
    .ZN(_00172_)
  );
  AND2_X1 _37499_ (
    .A1(reg_next_pc[20]),
    .A2(_02914_),
    .ZN(_03220_)
  );
  INV_X1 _37500_ (
    .A(_03220_),
    .ZN(_03221_)
  );
  AND2_X1 _37501_ (
    .A1(_21067_),
    .A2(_22097_),
    .ZN(_03222_)
  );
  INV_X1 _37502_ (
    .A(_03222_),
    .ZN(_03223_)
  );
  AND2_X1 _37503_ (
    .A1(latched_stalu),
    .A2(_22132_),
    .ZN(_03224_)
  );
  INV_X1 _37504_ (
    .A(_03224_),
    .ZN(_03225_)
  );
  AND2_X1 _37505_ (
    .A1(_03223_),
    .A2(_03225_),
    .ZN(_03226_)
  );
  AND2_X1 _37506_ (
    .A1(_02913_),
    .A2(_03226_),
    .ZN(_03227_)
  );
  INV_X1 _37507_ (
    .A(_03227_),
    .ZN(_03228_)
  );
  AND2_X1 _37508_ (
    .A1(_03221_),
    .A2(_03228_),
    .ZN(_03229_)
  );
  INV_X1 _37509_ (
    .A(_03229_),
    .ZN(_03230_)
  );
  AND2_X1 _37510_ (
    .A1(_02911_),
    .A2(_03230_),
    .ZN(_03231_)
  );
  INV_X1 _37511_ (
    .A(_03231_),
    .ZN(_03232_)
  );
  AND2_X1 _37512_ (
    .A1(reg_pc[20]),
    .A2(_02928_),
    .ZN(_03233_)
  );
  INV_X1 _37513_ (
    .A(_03233_),
    .ZN(_03234_)
  );
  AND2_X1 _37514_ (
    .A1(_03232_),
    .A2(_03234_),
    .ZN(_03235_)
  );
  INV_X1 _37515_ (
    .A(_03235_),
    .ZN(_00173_)
  );
  AND2_X1 _37516_ (
    .A1(reg_next_pc[21]),
    .A2(_02914_),
    .ZN(_03236_)
  );
  INV_X1 _37517_ (
    .A(_03236_),
    .ZN(_03237_)
  );
  AND2_X1 _37518_ (
    .A1(_21067_),
    .A2(_22098_),
    .ZN(_03238_)
  );
  INV_X1 _37519_ (
    .A(_03238_),
    .ZN(_03239_)
  );
  AND2_X1 _37520_ (
    .A1(latched_stalu),
    .A2(_22133_),
    .ZN(_03240_)
  );
  INV_X1 _37521_ (
    .A(_03240_),
    .ZN(_03241_)
  );
  AND2_X1 _37522_ (
    .A1(_03239_),
    .A2(_03241_),
    .ZN(_03242_)
  );
  AND2_X1 _37523_ (
    .A1(_02913_),
    .A2(_03242_),
    .ZN(_03243_)
  );
  INV_X1 _37524_ (
    .A(_03243_),
    .ZN(_03244_)
  );
  AND2_X1 _37525_ (
    .A1(_03237_),
    .A2(_03244_),
    .ZN(_03245_)
  );
  INV_X1 _37526_ (
    .A(_03245_),
    .ZN(_03246_)
  );
  AND2_X1 _37527_ (
    .A1(_02911_),
    .A2(_03246_),
    .ZN(_03247_)
  );
  INV_X1 _37528_ (
    .A(_03247_),
    .ZN(_03248_)
  );
  AND2_X1 _37529_ (
    .A1(reg_pc[21]),
    .A2(_02928_),
    .ZN(_03249_)
  );
  INV_X1 _37530_ (
    .A(_03249_),
    .ZN(_03250_)
  );
  AND2_X1 _37531_ (
    .A1(_03248_),
    .A2(_03250_),
    .ZN(_03251_)
  );
  INV_X1 _37532_ (
    .A(_03251_),
    .ZN(_00174_)
  );
  AND2_X1 _37533_ (
    .A1(reg_next_pc[22]),
    .A2(_02914_),
    .ZN(_03252_)
  );
  INV_X1 _37534_ (
    .A(_03252_),
    .ZN(_03253_)
  );
  AND2_X1 _37535_ (
    .A1(_21067_),
    .A2(_22099_),
    .ZN(_03254_)
  );
  INV_X1 _37536_ (
    .A(_03254_),
    .ZN(_03255_)
  );
  AND2_X1 _37537_ (
    .A1(latched_stalu),
    .A2(_22134_),
    .ZN(_03256_)
  );
  INV_X1 _37538_ (
    .A(_03256_),
    .ZN(_03257_)
  );
  AND2_X1 _37539_ (
    .A1(_03255_),
    .A2(_03257_),
    .ZN(_03258_)
  );
  AND2_X1 _37540_ (
    .A1(_02913_),
    .A2(_03258_),
    .ZN(_03259_)
  );
  INV_X1 _37541_ (
    .A(_03259_),
    .ZN(_03260_)
  );
  AND2_X1 _37542_ (
    .A1(_03253_),
    .A2(_03260_),
    .ZN(_03261_)
  );
  INV_X1 _37543_ (
    .A(_03261_),
    .ZN(_03262_)
  );
  AND2_X1 _37544_ (
    .A1(_02911_),
    .A2(_03262_),
    .ZN(_03263_)
  );
  INV_X1 _37545_ (
    .A(_03263_),
    .ZN(_03264_)
  );
  AND2_X1 _37546_ (
    .A1(reg_pc[22]),
    .A2(_02928_),
    .ZN(_03265_)
  );
  INV_X1 _37547_ (
    .A(_03265_),
    .ZN(_03266_)
  );
  AND2_X1 _37548_ (
    .A1(_03264_),
    .A2(_03266_),
    .ZN(_03267_)
  );
  INV_X1 _37549_ (
    .A(_03267_),
    .ZN(_00175_)
  );
  AND2_X1 _37550_ (
    .A1(reg_next_pc[23]),
    .A2(_02914_),
    .ZN(_03268_)
  );
  INV_X1 _37551_ (
    .A(_03268_),
    .ZN(_03269_)
  );
  AND2_X1 _37552_ (
    .A1(_21067_),
    .A2(_22100_),
    .ZN(_03270_)
  );
  INV_X1 _37553_ (
    .A(_03270_),
    .ZN(_03271_)
  );
  AND2_X1 _37554_ (
    .A1(latched_stalu),
    .A2(_22135_),
    .ZN(_03272_)
  );
  INV_X1 _37555_ (
    .A(_03272_),
    .ZN(_03273_)
  );
  AND2_X1 _37556_ (
    .A1(_03271_),
    .A2(_03273_),
    .ZN(_03274_)
  );
  AND2_X1 _37557_ (
    .A1(_02913_),
    .A2(_03274_),
    .ZN(_03275_)
  );
  INV_X1 _37558_ (
    .A(_03275_),
    .ZN(_03276_)
  );
  AND2_X1 _37559_ (
    .A1(_03269_),
    .A2(_03276_),
    .ZN(_03277_)
  );
  INV_X1 _37560_ (
    .A(_03277_),
    .ZN(_03278_)
  );
  AND2_X1 _37561_ (
    .A1(_02911_),
    .A2(_03278_),
    .ZN(_03279_)
  );
  INV_X1 _37562_ (
    .A(_03279_),
    .ZN(_03280_)
  );
  AND2_X1 _37563_ (
    .A1(reg_pc[23]),
    .A2(_02928_),
    .ZN(_03281_)
  );
  INV_X1 _37564_ (
    .A(_03281_),
    .ZN(_03282_)
  );
  AND2_X1 _37565_ (
    .A1(_03280_),
    .A2(_03282_),
    .ZN(_03283_)
  );
  INV_X1 _37566_ (
    .A(_03283_),
    .ZN(_00176_)
  );
  AND2_X1 _37567_ (
    .A1(reg_next_pc[24]),
    .A2(_02914_),
    .ZN(_03284_)
  );
  INV_X1 _37568_ (
    .A(_03284_),
    .ZN(_03285_)
  );
  AND2_X1 _37569_ (
    .A1(_21067_),
    .A2(_22101_),
    .ZN(_03286_)
  );
  INV_X1 _37570_ (
    .A(_03286_),
    .ZN(_03287_)
  );
  AND2_X1 _37571_ (
    .A1(latched_stalu),
    .A2(_22136_),
    .ZN(_03288_)
  );
  INV_X1 _37572_ (
    .A(_03288_),
    .ZN(_03289_)
  );
  AND2_X1 _37573_ (
    .A1(_03287_),
    .A2(_03289_),
    .ZN(_03290_)
  );
  AND2_X1 _37574_ (
    .A1(_02913_),
    .A2(_03290_),
    .ZN(_03291_)
  );
  INV_X1 _37575_ (
    .A(_03291_),
    .ZN(_03292_)
  );
  AND2_X1 _37576_ (
    .A1(_03285_),
    .A2(_03292_),
    .ZN(_03293_)
  );
  INV_X1 _37577_ (
    .A(_03293_),
    .ZN(_03294_)
  );
  AND2_X1 _37578_ (
    .A1(_02911_),
    .A2(_03294_),
    .ZN(_03295_)
  );
  INV_X1 _37579_ (
    .A(_03295_),
    .ZN(_03296_)
  );
  AND2_X1 _37580_ (
    .A1(reg_pc[24]),
    .A2(_02928_),
    .ZN(_03297_)
  );
  INV_X1 _37581_ (
    .A(_03297_),
    .ZN(_03298_)
  );
  AND2_X1 _37582_ (
    .A1(_03296_),
    .A2(_03298_),
    .ZN(_03299_)
  );
  INV_X1 _37583_ (
    .A(_03299_),
    .ZN(_00177_)
  );
  AND2_X1 _37584_ (
    .A1(reg_next_pc[25]),
    .A2(_02914_),
    .ZN(_03300_)
  );
  INV_X1 _37585_ (
    .A(_03300_),
    .ZN(_03301_)
  );
  AND2_X1 _37586_ (
    .A1(_21067_),
    .A2(_22102_),
    .ZN(_03302_)
  );
  INV_X1 _37587_ (
    .A(_03302_),
    .ZN(_03303_)
  );
  AND2_X1 _37588_ (
    .A1(latched_stalu),
    .A2(_22137_),
    .ZN(_03304_)
  );
  INV_X1 _37589_ (
    .A(_03304_),
    .ZN(_03305_)
  );
  AND2_X1 _37590_ (
    .A1(_03303_),
    .A2(_03305_),
    .ZN(_03306_)
  );
  AND2_X1 _37591_ (
    .A1(_02913_),
    .A2(_03306_),
    .ZN(_03307_)
  );
  INV_X1 _37592_ (
    .A(_03307_),
    .ZN(_03308_)
  );
  AND2_X1 _37593_ (
    .A1(_03301_),
    .A2(_03308_),
    .ZN(_03309_)
  );
  INV_X1 _37594_ (
    .A(_03309_),
    .ZN(_03310_)
  );
  AND2_X1 _37595_ (
    .A1(_02911_),
    .A2(_03310_),
    .ZN(_03311_)
  );
  INV_X1 _37596_ (
    .A(_03311_),
    .ZN(_03312_)
  );
  AND2_X1 _37597_ (
    .A1(reg_pc[25]),
    .A2(_02928_),
    .ZN(_03313_)
  );
  INV_X1 _37598_ (
    .A(_03313_),
    .ZN(_03314_)
  );
  AND2_X1 _37599_ (
    .A1(_03312_),
    .A2(_03314_),
    .ZN(_03315_)
  );
  INV_X1 _37600_ (
    .A(_03315_),
    .ZN(_00178_)
  );
  AND2_X1 _37601_ (
    .A1(reg_next_pc[26]),
    .A2(_02914_),
    .ZN(_03316_)
  );
  INV_X1 _37602_ (
    .A(_03316_),
    .ZN(_03317_)
  );
  AND2_X1 _37603_ (
    .A1(_21067_),
    .A2(_22103_),
    .ZN(_03318_)
  );
  INV_X1 _37604_ (
    .A(_03318_),
    .ZN(_03319_)
  );
  AND2_X1 _37605_ (
    .A1(latched_stalu),
    .A2(_22138_),
    .ZN(_03320_)
  );
  INV_X1 _37606_ (
    .A(_03320_),
    .ZN(_03321_)
  );
  AND2_X1 _37607_ (
    .A1(_03319_),
    .A2(_03321_),
    .ZN(_03322_)
  );
  AND2_X1 _37608_ (
    .A1(_02913_),
    .A2(_03322_),
    .ZN(_03323_)
  );
  INV_X1 _37609_ (
    .A(_03323_),
    .ZN(_03324_)
  );
  AND2_X1 _37610_ (
    .A1(_03317_),
    .A2(_03324_),
    .ZN(_03325_)
  );
  INV_X1 _37611_ (
    .A(_03325_),
    .ZN(_03326_)
  );
  AND2_X1 _37612_ (
    .A1(_02911_),
    .A2(_03326_),
    .ZN(_03327_)
  );
  INV_X1 _37613_ (
    .A(_03327_),
    .ZN(_03328_)
  );
  AND2_X1 _37614_ (
    .A1(reg_pc[26]),
    .A2(_02928_),
    .ZN(_03329_)
  );
  INV_X1 _37615_ (
    .A(_03329_),
    .ZN(_03330_)
  );
  AND2_X1 _37616_ (
    .A1(_03328_),
    .A2(_03330_),
    .ZN(_03331_)
  );
  INV_X1 _37617_ (
    .A(_03331_),
    .ZN(_00179_)
  );
  AND2_X1 _37618_ (
    .A1(reg_next_pc[27]),
    .A2(_02914_),
    .ZN(_03332_)
  );
  INV_X1 _37619_ (
    .A(_03332_),
    .ZN(_03333_)
  );
  AND2_X1 _37620_ (
    .A1(_21067_),
    .A2(_22104_),
    .ZN(_03334_)
  );
  INV_X1 _37621_ (
    .A(_03334_),
    .ZN(_03335_)
  );
  AND2_X1 _37622_ (
    .A1(latched_stalu),
    .A2(_22139_),
    .ZN(_03336_)
  );
  INV_X1 _37623_ (
    .A(_03336_),
    .ZN(_03337_)
  );
  AND2_X1 _37624_ (
    .A1(_03335_),
    .A2(_03337_),
    .ZN(_03338_)
  );
  AND2_X1 _37625_ (
    .A1(_02913_),
    .A2(_03338_),
    .ZN(_03339_)
  );
  INV_X1 _37626_ (
    .A(_03339_),
    .ZN(_03340_)
  );
  AND2_X1 _37627_ (
    .A1(_03333_),
    .A2(_03340_),
    .ZN(_03341_)
  );
  INV_X1 _37628_ (
    .A(_03341_),
    .ZN(_03342_)
  );
  AND2_X1 _37629_ (
    .A1(_02911_),
    .A2(_03342_),
    .ZN(_03343_)
  );
  INV_X1 _37630_ (
    .A(_03343_),
    .ZN(_03344_)
  );
  AND2_X1 _37631_ (
    .A1(reg_pc[27]),
    .A2(_02928_),
    .ZN(_03345_)
  );
  INV_X1 _37632_ (
    .A(_03345_),
    .ZN(_03346_)
  );
  AND2_X1 _37633_ (
    .A1(_03344_),
    .A2(_03346_),
    .ZN(_03347_)
  );
  INV_X1 _37634_ (
    .A(_03347_),
    .ZN(_00180_)
  );
  AND2_X1 _37635_ (
    .A1(reg_next_pc[28]),
    .A2(_02914_),
    .ZN(_03348_)
  );
  INV_X1 _37636_ (
    .A(_03348_),
    .ZN(_03349_)
  );
  AND2_X1 _37637_ (
    .A1(_21067_),
    .A2(_22105_),
    .ZN(_03350_)
  );
  INV_X1 _37638_ (
    .A(_03350_),
    .ZN(_03351_)
  );
  AND2_X1 _37639_ (
    .A1(latched_stalu),
    .A2(_22140_),
    .ZN(_03352_)
  );
  INV_X1 _37640_ (
    .A(_03352_),
    .ZN(_03353_)
  );
  AND2_X1 _37641_ (
    .A1(_03351_),
    .A2(_03353_),
    .ZN(_03354_)
  );
  AND2_X1 _37642_ (
    .A1(_02913_),
    .A2(_03354_),
    .ZN(_03355_)
  );
  INV_X1 _37643_ (
    .A(_03355_),
    .ZN(_03356_)
  );
  AND2_X1 _37644_ (
    .A1(_03349_),
    .A2(_03356_),
    .ZN(_03357_)
  );
  INV_X1 _37645_ (
    .A(_03357_),
    .ZN(_03358_)
  );
  AND2_X1 _37646_ (
    .A1(_02911_),
    .A2(_03358_),
    .ZN(_03359_)
  );
  INV_X1 _37647_ (
    .A(_03359_),
    .ZN(_03360_)
  );
  AND2_X1 _37648_ (
    .A1(reg_pc[28]),
    .A2(_02928_),
    .ZN(_03361_)
  );
  INV_X1 _37649_ (
    .A(_03361_),
    .ZN(_03362_)
  );
  AND2_X1 _37650_ (
    .A1(_03360_),
    .A2(_03362_),
    .ZN(_03363_)
  );
  INV_X1 _37651_ (
    .A(_03363_),
    .ZN(_00181_)
  );
  AND2_X1 _37652_ (
    .A1(reg_next_pc[29]),
    .A2(_02914_),
    .ZN(_03364_)
  );
  INV_X1 _37653_ (
    .A(_03364_),
    .ZN(_03365_)
  );
  AND2_X1 _37654_ (
    .A1(_21067_),
    .A2(_22106_),
    .ZN(_03366_)
  );
  INV_X1 _37655_ (
    .A(_03366_),
    .ZN(_03367_)
  );
  AND2_X1 _37656_ (
    .A1(latched_stalu),
    .A2(_22141_),
    .ZN(_03368_)
  );
  INV_X1 _37657_ (
    .A(_03368_),
    .ZN(_03369_)
  );
  AND2_X1 _37658_ (
    .A1(_03367_),
    .A2(_03369_),
    .ZN(_03370_)
  );
  AND2_X1 _37659_ (
    .A1(_02913_),
    .A2(_03370_),
    .ZN(_03371_)
  );
  INV_X1 _37660_ (
    .A(_03371_),
    .ZN(_03372_)
  );
  AND2_X1 _37661_ (
    .A1(_03365_),
    .A2(_03372_),
    .ZN(_03373_)
  );
  INV_X1 _37662_ (
    .A(_03373_),
    .ZN(_03374_)
  );
  AND2_X1 _37663_ (
    .A1(_02911_),
    .A2(_03374_),
    .ZN(_03375_)
  );
  INV_X1 _37664_ (
    .A(_03375_),
    .ZN(_03376_)
  );
  AND2_X1 _37665_ (
    .A1(reg_pc[29]),
    .A2(_02928_),
    .ZN(_03377_)
  );
  INV_X1 _37666_ (
    .A(_03377_),
    .ZN(_03378_)
  );
  AND2_X1 _37667_ (
    .A1(_03376_),
    .A2(_03378_),
    .ZN(_03379_)
  );
  INV_X1 _37668_ (
    .A(_03379_),
    .ZN(_00182_)
  );
  AND2_X1 _37669_ (
    .A1(reg_next_pc[30]),
    .A2(_02914_),
    .ZN(_03380_)
  );
  INV_X1 _37670_ (
    .A(_03380_),
    .ZN(_03381_)
  );
  AND2_X1 _37671_ (
    .A1(_21067_),
    .A2(_22107_),
    .ZN(_03382_)
  );
  INV_X1 _37672_ (
    .A(_03382_),
    .ZN(_03383_)
  );
  AND2_X1 _37673_ (
    .A1(latched_stalu),
    .A2(_22142_),
    .ZN(_03384_)
  );
  INV_X1 _37674_ (
    .A(_03384_),
    .ZN(_03385_)
  );
  AND2_X1 _37675_ (
    .A1(_03383_),
    .A2(_03385_),
    .ZN(_03386_)
  );
  AND2_X1 _37676_ (
    .A1(_02913_),
    .A2(_03386_),
    .ZN(_03387_)
  );
  INV_X1 _37677_ (
    .A(_03387_),
    .ZN(_03388_)
  );
  AND2_X1 _37678_ (
    .A1(_03381_),
    .A2(_03388_),
    .ZN(_03389_)
  );
  INV_X1 _37679_ (
    .A(_03389_),
    .ZN(_03390_)
  );
  AND2_X1 _37680_ (
    .A1(_02911_),
    .A2(_03390_),
    .ZN(_03391_)
  );
  INV_X1 _37681_ (
    .A(_03391_),
    .ZN(_03392_)
  );
  AND2_X1 _37682_ (
    .A1(reg_pc[30]),
    .A2(_02928_),
    .ZN(_03393_)
  );
  INV_X1 _37683_ (
    .A(_03393_),
    .ZN(_03394_)
  );
  AND2_X1 _37684_ (
    .A1(_03392_),
    .A2(_03394_),
    .ZN(_03395_)
  );
  INV_X1 _37685_ (
    .A(_03395_),
    .ZN(_00183_)
  );
  AND2_X1 _37686_ (
    .A1(reg_next_pc[31]),
    .A2(_02914_),
    .ZN(_03396_)
  );
  INV_X1 _37687_ (
    .A(_03396_),
    .ZN(_03397_)
  );
  AND2_X1 _37688_ (
    .A1(_21067_),
    .A2(_22108_),
    .ZN(_03398_)
  );
  INV_X1 _37689_ (
    .A(_03398_),
    .ZN(_03399_)
  );
  AND2_X1 _37690_ (
    .A1(latched_stalu),
    .A2(_22143_),
    .ZN(_03400_)
  );
  INV_X1 _37691_ (
    .A(_03400_),
    .ZN(_03401_)
  );
  AND2_X1 _37692_ (
    .A1(_03399_),
    .A2(_03401_),
    .ZN(_03402_)
  );
  AND2_X1 _37693_ (
    .A1(_02913_),
    .A2(_03402_),
    .ZN(_03403_)
  );
  INV_X1 _37694_ (
    .A(_03403_),
    .ZN(_03404_)
  );
  AND2_X1 _37695_ (
    .A1(_03397_),
    .A2(_03404_),
    .ZN(_03405_)
  );
  INV_X1 _37696_ (
    .A(_03405_),
    .ZN(_03406_)
  );
  AND2_X1 _37697_ (
    .A1(_02911_),
    .A2(_03406_),
    .ZN(_03407_)
  );
  INV_X1 _37698_ (
    .A(_03407_),
    .ZN(_03408_)
  );
  AND2_X1 _37699_ (
    .A1(reg_pc[31]),
    .A2(_02928_),
    .ZN(_03409_)
  );
  INV_X1 _37700_ (
    .A(_03409_),
    .ZN(_03410_)
  );
  AND2_X1 _37701_ (
    .A1(_03408_),
    .A2(_03410_),
    .ZN(_03411_)
  );
  INV_X1 _37702_ (
    .A(_03411_),
    .ZN(_00184_)
  );
  AND2_X1 _37703_ (
    .A1(instr_jal),
    .A2(decoded_rs2[1]),
    .ZN(_03412_)
  );
  INV_X1 _37704_ (
    .A(_03412_),
    .ZN(_03413_)
  );
  AND2_X1 _37705_ (
    .A1(decoder_trigger),
    .A2(_03412_),
    .ZN(_03414_)
  );
  INV_X1 _37706_ (
    .A(_03414_),
    .ZN(_03415_)
  );
  AND2_X1 _37707_ (
    .A1(reg_next_pc[1]),
    .A2(resetn),
    .ZN(_03416_)
  );
  INV_X1 _37708_ (
    .A(_03416_),
    .ZN(_03417_)
  );
  AND2_X1 _37709_ (
    .A1(_02912_),
    .A2(_03417_),
    .ZN(_03418_)
  );
  INV_X1 _37710_ (
    .A(_03418_),
    .ZN(_03419_)
  );
  AND2_X1 _37711_ (
    .A1(_02926_),
    .A2(_03415_),
    .ZN(_03420_)
  );
  INV_X1 _37712_ (
    .A(_03420_),
    .ZN(_03421_)
  );
  AND2_X1 _37713_ (
    .A1(_02927_),
    .A2(_03414_),
    .ZN(_03422_)
  );
  INV_X1 _37714_ (
    .A(_03422_),
    .ZN(_03423_)
  );
  AND2_X1 _37715_ (
    .A1(_03421_),
    .A2(_03423_),
    .ZN(_03424_)
  );
  AND2_X1 _37716_ (
    .A1(_02464_),
    .A2(_03424_),
    .ZN(_03425_)
  );
  INV_X1 _37717_ (
    .A(_03425_),
    .ZN(_03426_)
  );
  AND2_X1 _37718_ (
    .A1(_03419_),
    .A2(_03426_),
    .ZN(_00185_)
  );
  AND2_X1 _37719_ (
    .A1(decoded_rs2[1]),
    .A2(_02926_),
    .ZN(_03427_)
  );
  INV_X1 _37720_ (
    .A(_03427_),
    .ZN(_03428_)
  );
  AND2_X1 _37721_ (
    .A1(decoded_rs2[2]),
    .A2(_02943_),
    .ZN(_03429_)
  );
  INV_X1 _37722_ (
    .A(_03429_),
    .ZN(_03430_)
  );
  AND2_X1 _37723_ (
    .A1(_21284_),
    .A2(_02944_),
    .ZN(_03431_)
  );
  INV_X1 _37724_ (
    .A(_03431_),
    .ZN(_03432_)
  );
  AND2_X1 _37725_ (
    .A1(_03430_),
    .A2(_03432_),
    .ZN(_03433_)
  );
  INV_X1 _37726_ (
    .A(_03433_),
    .ZN(_03434_)
  );
  AND2_X1 _37727_ (
    .A1(_03427_),
    .A2(_03433_),
    .ZN(_03435_)
  );
  INV_X1 _37728_ (
    .A(_03435_),
    .ZN(_03436_)
  );
  AND2_X1 _37729_ (
    .A1(_03428_),
    .A2(_03434_),
    .ZN(_03437_)
  );
  INV_X1 _37730_ (
    .A(_03437_),
    .ZN(_03438_)
  );
  AND2_X1 _37731_ (
    .A1(_21261_),
    .A2(_02944_),
    .ZN(_03439_)
  );
  INV_X1 _37732_ (
    .A(_03439_),
    .ZN(_03440_)
  );
  AND2_X1 _37733_ (
    .A1(decoder_trigger),
    .A2(_03440_),
    .ZN(_03441_)
  );
  AND2_X1 _37734_ (
    .A1(instr_jal),
    .A2(_03436_),
    .ZN(_03442_)
  );
  AND2_X1 _37735_ (
    .A1(_03438_),
    .A2(_03442_),
    .ZN(_03443_)
  );
  INV_X1 _37736_ (
    .A(_03443_),
    .ZN(_03444_)
  );
  AND2_X1 _37737_ (
    .A1(_03441_),
    .A2(_03444_),
    .ZN(_03445_)
  );
  INV_X1 _37738_ (
    .A(_03445_),
    .ZN(_03446_)
  );
  AND2_X1 _37739_ (
    .A1(_02470_),
    .A2(_02944_),
    .ZN(_03447_)
  );
  INV_X1 _37740_ (
    .A(_03447_),
    .ZN(_03448_)
  );
  AND2_X1 _37741_ (
    .A1(_03446_),
    .A2(_03448_),
    .ZN(_03449_)
  );
  INV_X1 _37742_ (
    .A(_03449_),
    .ZN(_03450_)
  );
  AND2_X1 _37743_ (
    .A1(reg_next_pc[2]),
    .A2(_02928_),
    .ZN(_03451_)
  );
  INV_X1 _37744_ (
    .A(_03451_),
    .ZN(_03452_)
  );
  AND2_X1 _37745_ (
    .A1(_03450_),
    .A2(_03452_),
    .ZN(_03453_)
  );
  INV_X1 _37746_ (
    .A(_03453_),
    .ZN(_00186_)
  );
  AND2_X1 _37747_ (
    .A1(reg_next_pc[3]),
    .A2(_02928_),
    .ZN(_03454_)
  );
  INV_X1 _37748_ (
    .A(_03454_),
    .ZN(_03455_)
  );
  AND2_X1 _37749_ (
    .A1(_03430_),
    .A2(_03436_),
    .ZN(_03456_)
  );
  INV_X1 _37750_ (
    .A(_03456_),
    .ZN(_03457_)
  );
  AND2_X1 _37751_ (
    .A1(decoded_rs2[3]),
    .A2(_02959_),
    .ZN(_03458_)
  );
  INV_X1 _37752_ (
    .A(_03458_),
    .ZN(_03459_)
  );
  AND2_X1 _37753_ (
    .A1(_21285_),
    .A2(_02960_),
    .ZN(_03460_)
  );
  INV_X1 _37754_ (
    .A(_03460_),
    .ZN(_03461_)
  );
  AND2_X1 _37755_ (
    .A1(_03459_),
    .A2(_03461_),
    .ZN(_03462_)
  );
  INV_X1 _37756_ (
    .A(_03462_),
    .ZN(_03463_)
  );
  AND2_X1 _37757_ (
    .A1(_03457_),
    .A2(_03462_),
    .ZN(_03464_)
  );
  INV_X1 _37758_ (
    .A(_03464_),
    .ZN(_03465_)
  );
  AND2_X1 _37759_ (
    .A1(_03456_),
    .A2(_03463_),
    .ZN(_03466_)
  );
  INV_X1 _37760_ (
    .A(_03466_),
    .ZN(_03467_)
  );
  AND2_X1 _37761_ (
    .A1(instr_jal),
    .A2(_03467_),
    .ZN(_03468_)
  );
  AND2_X1 _37762_ (
    .A1(_03465_),
    .A2(_03468_),
    .ZN(_03469_)
  );
  INV_X1 _37763_ (
    .A(_03469_),
    .ZN(_03470_)
  );
  AND2_X1 _37764_ (
    .A1(_02944_),
    .A2(_02960_),
    .ZN(_03471_)
  );
  INV_X1 _37765_ (
    .A(_03471_),
    .ZN(_03472_)
  );
  AND2_X1 _37766_ (
    .A1(_02943_),
    .A2(_02958_),
    .ZN(_03473_)
  );
  INV_X1 _37767_ (
    .A(_03473_),
    .ZN(_03474_)
  );
  AND2_X1 _37768_ (
    .A1(_21261_),
    .A2(_03474_),
    .ZN(_03475_)
  );
  AND2_X1 _37769_ (
    .A1(_03472_),
    .A2(_03475_),
    .ZN(_03476_)
  );
  INV_X1 _37770_ (
    .A(_03476_),
    .ZN(_03477_)
  );
  AND2_X1 _37771_ (
    .A1(decoder_trigger),
    .A2(_03477_),
    .ZN(_03478_)
  );
  AND2_X1 _37772_ (
    .A1(_03470_),
    .A2(_03478_),
    .ZN(_03479_)
  );
  INV_X1 _37773_ (
    .A(_03479_),
    .ZN(_03480_)
  );
  AND2_X1 _37774_ (
    .A1(_02470_),
    .A2(_02960_),
    .ZN(_03481_)
  );
  INV_X1 _37775_ (
    .A(_03481_),
    .ZN(_03482_)
  );
  AND2_X1 _37776_ (
    .A1(_03480_),
    .A2(_03482_),
    .ZN(_03483_)
  );
  INV_X1 _37777_ (
    .A(_03483_),
    .ZN(_03484_)
  );
  AND2_X1 _37778_ (
    .A1(_03455_),
    .A2(_03484_),
    .ZN(_03485_)
  );
  INV_X1 _37779_ (
    .A(_03485_),
    .ZN(_00187_)
  );
  AND2_X1 _37780_ (
    .A1(reg_next_pc[4]),
    .A2(_02928_),
    .ZN(_03486_)
  );
  INV_X1 _37781_ (
    .A(_03486_),
    .ZN(_03487_)
  );
  AND2_X1 _37782_ (
    .A1(_03459_),
    .A2(_03465_),
    .ZN(_03488_)
  );
  INV_X1 _37783_ (
    .A(_03488_),
    .ZN(_03489_)
  );
  AND2_X1 _37784_ (
    .A1(decoded_imm_j[4]),
    .A2(_02975_),
    .ZN(_03490_)
  );
  INV_X1 _37785_ (
    .A(_03490_),
    .ZN(_03491_)
  );
  AND2_X1 _37786_ (
    .A1(_22015_),
    .A2(_02976_),
    .ZN(_03492_)
  );
  INV_X1 _37787_ (
    .A(_03492_),
    .ZN(_03493_)
  );
  AND2_X1 _37788_ (
    .A1(_03491_),
    .A2(_03493_),
    .ZN(_03494_)
  );
  INV_X1 _37789_ (
    .A(_03494_),
    .ZN(_03495_)
  );
  AND2_X1 _37790_ (
    .A1(_03488_),
    .A2(_03495_),
    .ZN(_03496_)
  );
  INV_X1 _37791_ (
    .A(_03496_),
    .ZN(_03497_)
  );
  AND2_X1 _37792_ (
    .A1(_03489_),
    .A2(_03494_),
    .ZN(_03498_)
  );
  INV_X1 _37793_ (
    .A(_03498_),
    .ZN(_03499_)
  );
  AND2_X1 _37794_ (
    .A1(_03497_),
    .A2(_03499_),
    .ZN(_03500_)
  );
  AND2_X1 _37795_ (
    .A1(instr_jal),
    .A2(_03500_),
    .ZN(_03501_)
  );
  INV_X1 _37796_ (
    .A(_03501_),
    .ZN(_03502_)
  );
  AND2_X1 _37797_ (
    .A1(_02974_),
    .A2(_03473_),
    .ZN(_03503_)
  );
  INV_X1 _37798_ (
    .A(_03503_),
    .ZN(_03504_)
  );
  AND2_X1 _37799_ (
    .A1(_02976_),
    .A2(_03474_),
    .ZN(_03505_)
  );
  INV_X1 _37800_ (
    .A(_03505_),
    .ZN(_03506_)
  );
  AND2_X1 _37801_ (
    .A1(_03504_),
    .A2(_03506_),
    .ZN(_03507_)
  );
  AND2_X1 _37802_ (
    .A1(_21261_),
    .A2(_03507_),
    .ZN(_03508_)
  );
  INV_X1 _37803_ (
    .A(_03508_),
    .ZN(_03509_)
  );
  AND2_X1 _37804_ (
    .A1(decoder_trigger),
    .A2(_03509_),
    .ZN(_03510_)
  );
  AND2_X1 _37805_ (
    .A1(_03502_),
    .A2(_03510_),
    .ZN(_03511_)
  );
  INV_X1 _37806_ (
    .A(_03511_),
    .ZN(_03512_)
  );
  AND2_X1 _37807_ (
    .A1(_02470_),
    .A2(_02976_),
    .ZN(_03513_)
  );
  INV_X1 _37808_ (
    .A(_03513_),
    .ZN(_03514_)
  );
  AND2_X1 _37809_ (
    .A1(_03512_),
    .A2(_03514_),
    .ZN(_03515_)
  );
  INV_X1 _37810_ (
    .A(_03515_),
    .ZN(_03516_)
  );
  AND2_X1 _37811_ (
    .A1(_03487_),
    .A2(_03516_),
    .ZN(_03517_)
  );
  INV_X1 _37812_ (
    .A(_03517_),
    .ZN(_00188_)
  );
  AND2_X1 _37813_ (
    .A1(reg_next_pc[5]),
    .A2(_02928_),
    .ZN(_03518_)
  );
  INV_X1 _37814_ (
    .A(_03518_),
    .ZN(_03519_)
  );
  AND2_X1 _37815_ (
    .A1(_03491_),
    .A2(_03499_),
    .ZN(_03520_)
  );
  INV_X1 _37816_ (
    .A(_03520_),
    .ZN(_03521_)
  );
  AND2_X1 _37817_ (
    .A1(decoded_imm_j[5]),
    .A2(_02991_),
    .ZN(_03522_)
  );
  INV_X1 _37818_ (
    .A(_03522_),
    .ZN(_03523_)
  );
  AND2_X1 _37819_ (
    .A1(_22011_),
    .A2(_02992_),
    .ZN(_03524_)
  );
  INV_X1 _37820_ (
    .A(_03524_),
    .ZN(_03525_)
  );
  AND2_X1 _37821_ (
    .A1(_03523_),
    .A2(_03525_),
    .ZN(_03526_)
  );
  INV_X1 _37822_ (
    .A(_03526_),
    .ZN(_03527_)
  );
  AND2_X1 _37823_ (
    .A1(_03521_),
    .A2(_03526_),
    .ZN(_03528_)
  );
  INV_X1 _37824_ (
    .A(_03528_),
    .ZN(_03529_)
  );
  AND2_X1 _37825_ (
    .A1(_03520_),
    .A2(_03527_),
    .ZN(_03530_)
  );
  INV_X1 _37826_ (
    .A(_03530_),
    .ZN(_03531_)
  );
  AND2_X1 _37827_ (
    .A1(_03529_),
    .A2(_03531_),
    .ZN(_03532_)
  );
  AND2_X1 _37828_ (
    .A1(_02991_),
    .A2(_03503_),
    .ZN(_03533_)
  );
  INV_X1 _37829_ (
    .A(_03533_),
    .ZN(_03534_)
  );
  AND2_X1 _37830_ (
    .A1(_02992_),
    .A2(_03504_),
    .ZN(_03535_)
  );
  INV_X1 _37831_ (
    .A(_03535_),
    .ZN(_03536_)
  );
  AND2_X1 _37832_ (
    .A1(_03534_),
    .A2(_03536_),
    .ZN(_03537_)
  );
  AND2_X1 _37833_ (
    .A1(_21261_),
    .A2(_03537_),
    .ZN(_03538_)
  );
  INV_X1 _37834_ (
    .A(_03538_),
    .ZN(_03539_)
  );
  AND2_X1 _37835_ (
    .A1(decoder_trigger),
    .A2(_03539_),
    .ZN(_03540_)
  );
  AND2_X1 _37836_ (
    .A1(instr_jal),
    .A2(_03532_),
    .ZN(_03541_)
  );
  INV_X1 _37837_ (
    .A(_03541_),
    .ZN(_03542_)
  );
  AND2_X1 _37838_ (
    .A1(_03540_),
    .A2(_03542_),
    .ZN(_03543_)
  );
  INV_X1 _37839_ (
    .A(_03543_),
    .ZN(_03544_)
  );
  AND2_X1 _37840_ (
    .A1(_02470_),
    .A2(_02992_),
    .ZN(_03545_)
  );
  INV_X1 _37841_ (
    .A(_03545_),
    .ZN(_03546_)
  );
  AND2_X1 _37842_ (
    .A1(_03544_),
    .A2(_03546_),
    .ZN(_03547_)
  );
  INV_X1 _37843_ (
    .A(_03547_),
    .ZN(_03548_)
  );
  AND2_X1 _37844_ (
    .A1(_03519_),
    .A2(_03548_),
    .ZN(_03549_)
  );
  INV_X1 _37845_ (
    .A(_03549_),
    .ZN(_00189_)
  );
  AND2_X1 _37846_ (
    .A1(reg_next_pc[6]),
    .A2(_02928_),
    .ZN(_03550_)
  );
  INV_X1 _37847_ (
    .A(_03550_),
    .ZN(_03551_)
  );
  AND2_X1 _37848_ (
    .A1(_03523_),
    .A2(_03529_),
    .ZN(_03552_)
  );
  INV_X1 _37849_ (
    .A(_03552_),
    .ZN(_03553_)
  );
  AND2_X1 _37850_ (
    .A1(decoded_imm_j[6]),
    .A2(_03007_),
    .ZN(_03554_)
  );
  INV_X1 _37851_ (
    .A(_03554_),
    .ZN(_03555_)
  );
  AND2_X1 _37852_ (
    .A1(_22010_),
    .A2(_03008_),
    .ZN(_03556_)
  );
  INV_X1 _37853_ (
    .A(_03556_),
    .ZN(_03557_)
  );
  AND2_X1 _37854_ (
    .A1(_03555_),
    .A2(_03557_),
    .ZN(_03558_)
  );
  INV_X1 _37855_ (
    .A(_03558_),
    .ZN(_03559_)
  );
  AND2_X1 _37856_ (
    .A1(_03552_),
    .A2(_03559_),
    .ZN(_03560_)
  );
  INV_X1 _37857_ (
    .A(_03560_),
    .ZN(_03561_)
  );
  AND2_X1 _37858_ (
    .A1(_03553_),
    .A2(_03558_),
    .ZN(_03562_)
  );
  INV_X1 _37859_ (
    .A(_03562_),
    .ZN(_03563_)
  );
  AND2_X1 _37860_ (
    .A1(_03561_),
    .A2(_03563_),
    .ZN(_03564_)
  );
  AND2_X1 _37861_ (
    .A1(instr_jal),
    .A2(_03564_),
    .ZN(_03565_)
  );
  INV_X1 _37862_ (
    .A(_03565_),
    .ZN(_03566_)
  );
  AND2_X1 _37863_ (
    .A1(_03006_),
    .A2(_03533_),
    .ZN(_03567_)
  );
  INV_X1 _37864_ (
    .A(_03567_),
    .ZN(_03568_)
  );
  AND2_X1 _37865_ (
    .A1(_03008_),
    .A2(_03534_),
    .ZN(_03569_)
  );
  INV_X1 _37866_ (
    .A(_03569_),
    .ZN(_03570_)
  );
  AND2_X1 _37867_ (
    .A1(_03568_),
    .A2(_03570_),
    .ZN(_03571_)
  );
  AND2_X1 _37868_ (
    .A1(_21261_),
    .A2(_03571_),
    .ZN(_03572_)
  );
  INV_X1 _37869_ (
    .A(_03572_),
    .ZN(_03573_)
  );
  AND2_X1 _37870_ (
    .A1(decoder_trigger),
    .A2(_03573_),
    .ZN(_03574_)
  );
  AND2_X1 _37871_ (
    .A1(_03566_),
    .A2(_03574_),
    .ZN(_03575_)
  );
  INV_X1 _37872_ (
    .A(_03575_),
    .ZN(_03576_)
  );
  AND2_X1 _37873_ (
    .A1(_02470_),
    .A2(_03008_),
    .ZN(_03577_)
  );
  INV_X1 _37874_ (
    .A(_03577_),
    .ZN(_03578_)
  );
  AND2_X1 _37875_ (
    .A1(_03576_),
    .A2(_03578_),
    .ZN(_03579_)
  );
  INV_X1 _37876_ (
    .A(_03579_),
    .ZN(_03580_)
  );
  AND2_X1 _37877_ (
    .A1(_03551_),
    .A2(_03580_),
    .ZN(_03581_)
  );
  INV_X1 _37878_ (
    .A(_03581_),
    .ZN(_00190_)
  );
  AND2_X1 _37879_ (
    .A1(reg_next_pc[7]),
    .A2(_02928_),
    .ZN(_03582_)
  );
  INV_X1 _37880_ (
    .A(_03582_),
    .ZN(_03583_)
  );
  AND2_X1 _37881_ (
    .A1(_03555_),
    .A2(_03563_),
    .ZN(_03584_)
  );
  INV_X1 _37882_ (
    .A(_03584_),
    .ZN(_03585_)
  );
  AND2_X1 _37883_ (
    .A1(decoded_imm_j[7]),
    .A2(_03023_),
    .ZN(_03586_)
  );
  INV_X1 _37884_ (
    .A(_03586_),
    .ZN(_03587_)
  );
  AND2_X1 _37885_ (
    .A1(_22009_),
    .A2(_03024_),
    .ZN(_03588_)
  );
  INV_X1 _37886_ (
    .A(_03588_),
    .ZN(_03589_)
  );
  AND2_X1 _37887_ (
    .A1(_03587_),
    .A2(_03589_),
    .ZN(_03590_)
  );
  INV_X1 _37888_ (
    .A(_03590_),
    .ZN(_03591_)
  );
  AND2_X1 _37889_ (
    .A1(_03585_),
    .A2(_03590_),
    .ZN(_03592_)
  );
  INV_X1 _37890_ (
    .A(_03592_),
    .ZN(_03593_)
  );
  AND2_X1 _37891_ (
    .A1(_03584_),
    .A2(_03591_),
    .ZN(_03594_)
  );
  INV_X1 _37892_ (
    .A(_03594_),
    .ZN(_03595_)
  );
  AND2_X1 _37893_ (
    .A1(instr_jal),
    .A2(_03595_),
    .ZN(_03596_)
  );
  AND2_X1 _37894_ (
    .A1(_03593_),
    .A2(_03596_),
    .ZN(_03597_)
  );
  INV_X1 _37895_ (
    .A(_03597_),
    .ZN(_03598_)
  );
  AND2_X1 _37896_ (
    .A1(_03023_),
    .A2(_03567_),
    .ZN(_03599_)
  );
  INV_X1 _37897_ (
    .A(_03599_),
    .ZN(_03600_)
  );
  AND2_X1 _37898_ (
    .A1(_03024_),
    .A2(_03568_),
    .ZN(_03601_)
  );
  INV_X1 _37899_ (
    .A(_03601_),
    .ZN(_03602_)
  );
  AND2_X1 _37900_ (
    .A1(_03600_),
    .A2(_03602_),
    .ZN(_03603_)
  );
  AND2_X1 _37901_ (
    .A1(_21261_),
    .A2(_03603_),
    .ZN(_03604_)
  );
  INV_X1 _37902_ (
    .A(_03604_),
    .ZN(_03605_)
  );
  AND2_X1 _37903_ (
    .A1(decoder_trigger),
    .A2(_03605_),
    .ZN(_03606_)
  );
  AND2_X1 _37904_ (
    .A1(_03598_),
    .A2(_03606_),
    .ZN(_03607_)
  );
  INV_X1 _37905_ (
    .A(_03607_),
    .ZN(_03608_)
  );
  AND2_X1 _37906_ (
    .A1(_02470_),
    .A2(_03024_),
    .ZN(_03609_)
  );
  INV_X1 _37907_ (
    .A(_03609_),
    .ZN(_03610_)
  );
  AND2_X1 _37908_ (
    .A1(_03608_),
    .A2(_03610_),
    .ZN(_03611_)
  );
  INV_X1 _37909_ (
    .A(_03611_),
    .ZN(_03612_)
  );
  AND2_X1 _37910_ (
    .A1(_03583_),
    .A2(_03612_),
    .ZN(_03613_)
  );
  INV_X1 _37911_ (
    .A(_03613_),
    .ZN(_00191_)
  );
  AND2_X1 _37912_ (
    .A1(reg_next_pc[8]),
    .A2(_02928_),
    .ZN(_03614_)
  );
  INV_X1 _37913_ (
    .A(_03614_),
    .ZN(_03615_)
  );
  AND2_X1 _37914_ (
    .A1(decoded_imm_j[8]),
    .A2(_03039_),
    .ZN(_03616_)
  );
  INV_X1 _37915_ (
    .A(_03616_),
    .ZN(_03617_)
  );
  AND2_X1 _37916_ (
    .A1(_22012_),
    .A2(_03040_),
    .ZN(_03618_)
  );
  INV_X1 _37917_ (
    .A(_03618_),
    .ZN(_03619_)
  );
  AND2_X1 _37918_ (
    .A1(_03617_),
    .A2(_03619_),
    .ZN(_03620_)
  );
  INV_X1 _37919_ (
    .A(_03620_),
    .ZN(_03621_)
  );
  AND2_X1 _37920_ (
    .A1(_03585_),
    .A2(_03589_),
    .ZN(_03622_)
  );
  INV_X1 _37921_ (
    .A(_03622_),
    .ZN(_03623_)
  );
  AND2_X1 _37922_ (
    .A1(_03584_),
    .A2(_03587_),
    .ZN(_03624_)
  );
  INV_X1 _37923_ (
    .A(_03624_),
    .ZN(_03625_)
  );
  AND2_X1 _37924_ (
    .A1(_03587_),
    .A2(_03623_),
    .ZN(_03626_)
  );
  AND2_X1 _37925_ (
    .A1(_03589_),
    .A2(_03625_),
    .ZN(_03627_)
  );
  AND2_X1 _37926_ (
    .A1(_03621_),
    .A2(_03626_),
    .ZN(_03628_)
  );
  INV_X1 _37927_ (
    .A(_03628_),
    .ZN(_03629_)
  );
  AND2_X1 _37928_ (
    .A1(_03620_),
    .A2(_03627_),
    .ZN(_03630_)
  );
  INV_X1 _37929_ (
    .A(_03630_),
    .ZN(_03631_)
  );
  AND2_X1 _37930_ (
    .A1(instr_jal),
    .A2(_03631_),
    .ZN(_03632_)
  );
  AND2_X1 _37931_ (
    .A1(_03629_),
    .A2(_03632_),
    .ZN(_03633_)
  );
  INV_X1 _37932_ (
    .A(_03633_),
    .ZN(_03634_)
  );
  AND2_X1 _37933_ (
    .A1(_03038_),
    .A2(_03599_),
    .ZN(_03635_)
  );
  INV_X1 _37934_ (
    .A(_03635_),
    .ZN(_03636_)
  );
  AND2_X1 _37935_ (
    .A1(_03040_),
    .A2(_03600_),
    .ZN(_03637_)
  );
  INV_X1 _37936_ (
    .A(_03637_),
    .ZN(_03638_)
  );
  AND2_X1 _37937_ (
    .A1(_03636_),
    .A2(_03638_),
    .ZN(_03639_)
  );
  AND2_X1 _37938_ (
    .A1(_21261_),
    .A2(_03639_),
    .ZN(_03640_)
  );
  INV_X1 _37939_ (
    .A(_03640_),
    .ZN(_03641_)
  );
  AND2_X1 _37940_ (
    .A1(decoder_trigger),
    .A2(_03641_),
    .ZN(_03642_)
  );
  AND2_X1 _37941_ (
    .A1(_03634_),
    .A2(_03642_),
    .ZN(_03643_)
  );
  INV_X1 _37942_ (
    .A(_03643_),
    .ZN(_03644_)
  );
  AND2_X1 _37943_ (
    .A1(_02470_),
    .A2(_03040_),
    .ZN(_03645_)
  );
  INV_X1 _37944_ (
    .A(_03645_),
    .ZN(_03646_)
  );
  AND2_X1 _37945_ (
    .A1(_03644_),
    .A2(_03646_),
    .ZN(_03647_)
  );
  INV_X1 _37946_ (
    .A(_03647_),
    .ZN(_03648_)
  );
  AND2_X1 _37947_ (
    .A1(_03615_),
    .A2(_03648_),
    .ZN(_03649_)
  );
  INV_X1 _37948_ (
    .A(_03649_),
    .ZN(_00192_)
  );
  AND2_X1 _37949_ (
    .A1(reg_next_pc[9]),
    .A2(_02928_),
    .ZN(_03650_)
  );
  INV_X1 _37950_ (
    .A(_03650_),
    .ZN(_03651_)
  );
  AND2_X1 _37951_ (
    .A1(_03617_),
    .A2(_03631_),
    .ZN(_03652_)
  );
  INV_X1 _37952_ (
    .A(_03652_),
    .ZN(_03653_)
  );
  AND2_X1 _37953_ (
    .A1(decoded_imm_j[9]),
    .A2(_03055_),
    .ZN(_03654_)
  );
  INV_X1 _37954_ (
    .A(_03654_),
    .ZN(_03655_)
  );
  AND2_X1 _37955_ (
    .A1(_22013_),
    .A2(_03056_),
    .ZN(_03656_)
  );
  INV_X1 _37956_ (
    .A(_03656_),
    .ZN(_03657_)
  );
  AND2_X1 _37957_ (
    .A1(_03655_),
    .A2(_03657_),
    .ZN(_03658_)
  );
  INV_X1 _37958_ (
    .A(_03658_),
    .ZN(_03659_)
  );
  AND2_X1 _37959_ (
    .A1(_03653_),
    .A2(_03658_),
    .ZN(_03660_)
  );
  INV_X1 _37960_ (
    .A(_03660_),
    .ZN(_03661_)
  );
  AND2_X1 _37961_ (
    .A1(_03652_),
    .A2(_03659_),
    .ZN(_03662_)
  );
  INV_X1 _37962_ (
    .A(_03662_),
    .ZN(_03663_)
  );
  AND2_X1 _37963_ (
    .A1(instr_jal),
    .A2(_03663_),
    .ZN(_03664_)
  );
  AND2_X1 _37964_ (
    .A1(_03661_),
    .A2(_03664_),
    .ZN(_03665_)
  );
  INV_X1 _37965_ (
    .A(_03665_),
    .ZN(_03666_)
  );
  AND2_X1 _37966_ (
    .A1(_03056_),
    .A2(_03636_),
    .ZN(_03667_)
  );
  INV_X1 _37967_ (
    .A(_03667_),
    .ZN(_03668_)
  );
  AND2_X1 _37968_ (
    .A1(_03055_),
    .A2(_03635_),
    .ZN(_03669_)
  );
  INV_X1 _37969_ (
    .A(_03669_),
    .ZN(_03670_)
  );
  AND2_X1 _37970_ (
    .A1(_21261_),
    .A2(_03670_),
    .ZN(_03671_)
  );
  AND2_X1 _37971_ (
    .A1(_03668_),
    .A2(_03671_),
    .ZN(_03672_)
  );
  INV_X1 _37972_ (
    .A(_03672_),
    .ZN(_03673_)
  );
  AND2_X1 _37973_ (
    .A1(decoder_trigger),
    .A2(_03673_),
    .ZN(_03674_)
  );
  AND2_X1 _37974_ (
    .A1(_03666_),
    .A2(_03674_),
    .ZN(_03675_)
  );
  INV_X1 _37975_ (
    .A(_03675_),
    .ZN(_03676_)
  );
  AND2_X1 _37976_ (
    .A1(_02470_),
    .A2(_03056_),
    .ZN(_03677_)
  );
  INV_X1 _37977_ (
    .A(_03677_),
    .ZN(_03678_)
  );
  AND2_X1 _37978_ (
    .A1(_03676_),
    .A2(_03678_),
    .ZN(_03679_)
  );
  INV_X1 _37979_ (
    .A(_03679_),
    .ZN(_03680_)
  );
  AND2_X1 _37980_ (
    .A1(_03651_),
    .A2(_03680_),
    .ZN(_03681_)
  );
  INV_X1 _37981_ (
    .A(_03681_),
    .ZN(_00193_)
  );
  AND2_X1 _37982_ (
    .A1(reg_next_pc[10]),
    .A2(_02928_),
    .ZN(_03682_)
  );
  INV_X1 _37983_ (
    .A(_03682_),
    .ZN(_03683_)
  );
  AND2_X1 _37984_ (
    .A1(decoded_imm_j[10]),
    .A2(_03071_),
    .ZN(_03684_)
  );
  INV_X1 _37985_ (
    .A(_03684_),
    .ZN(_03685_)
  );
  AND2_X1 _37986_ (
    .A1(_21287_),
    .A2(_03072_),
    .ZN(_03686_)
  );
  INV_X1 _37987_ (
    .A(_03686_),
    .ZN(_03687_)
  );
  AND2_X1 _37988_ (
    .A1(_03685_),
    .A2(_03687_),
    .ZN(_03688_)
  );
  INV_X1 _37989_ (
    .A(_03688_),
    .ZN(_03689_)
  );
  AND2_X1 _37990_ (
    .A1(_03652_),
    .A2(_03655_),
    .ZN(_03690_)
  );
  INV_X1 _37991_ (
    .A(_03690_),
    .ZN(_03691_)
  );
  AND2_X1 _37992_ (
    .A1(_03653_),
    .A2(_03657_),
    .ZN(_03692_)
  );
  INV_X1 _37993_ (
    .A(_03692_),
    .ZN(_03693_)
  );
  AND2_X1 _37994_ (
    .A1(_03657_),
    .A2(_03691_),
    .ZN(_03694_)
  );
  AND2_X1 _37995_ (
    .A1(_03655_),
    .A2(_03693_),
    .ZN(_03695_)
  );
  AND2_X1 _37996_ (
    .A1(_03689_),
    .A2(_03695_),
    .ZN(_03696_)
  );
  INV_X1 _37997_ (
    .A(_03696_),
    .ZN(_03697_)
  );
  AND2_X1 _37998_ (
    .A1(_03688_),
    .A2(_03694_),
    .ZN(_03698_)
  );
  INV_X1 _37999_ (
    .A(_03698_),
    .ZN(_03699_)
  );
  AND2_X1 _38000_ (
    .A1(instr_jal),
    .A2(_03699_),
    .ZN(_03700_)
  );
  AND2_X1 _38001_ (
    .A1(_03697_),
    .A2(_03700_),
    .ZN(_03701_)
  );
  INV_X1 _38002_ (
    .A(_03701_),
    .ZN(_03702_)
  );
  AND2_X1 _38003_ (
    .A1(_03070_),
    .A2(_03669_),
    .ZN(_03703_)
  );
  INV_X1 _38004_ (
    .A(_03703_),
    .ZN(_03704_)
  );
  AND2_X1 _38005_ (
    .A1(_03072_),
    .A2(_03670_),
    .ZN(_03705_)
  );
  INV_X1 _38006_ (
    .A(_03705_),
    .ZN(_03706_)
  );
  AND2_X1 _38007_ (
    .A1(_03704_),
    .A2(_03706_),
    .ZN(_03707_)
  );
  AND2_X1 _38008_ (
    .A1(_21261_),
    .A2(_03707_),
    .ZN(_03708_)
  );
  INV_X1 _38009_ (
    .A(_03708_),
    .ZN(_03709_)
  );
  AND2_X1 _38010_ (
    .A1(decoder_trigger),
    .A2(_03709_),
    .ZN(_03710_)
  );
  AND2_X1 _38011_ (
    .A1(_03702_),
    .A2(_03710_),
    .ZN(_03711_)
  );
  INV_X1 _38012_ (
    .A(_03711_),
    .ZN(_03712_)
  );
  AND2_X1 _38013_ (
    .A1(_02470_),
    .A2(_03072_),
    .ZN(_03713_)
  );
  INV_X1 _38014_ (
    .A(_03713_),
    .ZN(_03714_)
  );
  AND2_X1 _38015_ (
    .A1(_03712_),
    .A2(_03714_),
    .ZN(_03715_)
  );
  INV_X1 _38016_ (
    .A(_03715_),
    .ZN(_03716_)
  );
  AND2_X1 _38017_ (
    .A1(_03683_),
    .A2(_03716_),
    .ZN(_03717_)
  );
  INV_X1 _38018_ (
    .A(_03717_),
    .ZN(_00194_)
  );
  AND2_X1 _38019_ (
    .A1(reg_next_pc[11]),
    .A2(_02928_),
    .ZN(_03718_)
  );
  INV_X1 _38020_ (
    .A(_03718_),
    .ZN(_03719_)
  );
  AND2_X1 _38021_ (
    .A1(_03685_),
    .A2(_03699_),
    .ZN(_03720_)
  );
  INV_X1 _38022_ (
    .A(_03720_),
    .ZN(_03721_)
  );
  AND2_X1 _38023_ (
    .A1(decoded_rs2[0]),
    .A2(_03087_),
    .ZN(_03722_)
  );
  INV_X1 _38024_ (
    .A(_03722_),
    .ZN(_03723_)
  );
  AND2_X1 _38025_ (
    .A1(_21282_),
    .A2(_03088_),
    .ZN(_03724_)
  );
  INV_X1 _38026_ (
    .A(_03724_),
    .ZN(_03725_)
  );
  AND2_X1 _38027_ (
    .A1(_03723_),
    .A2(_03725_),
    .ZN(_03726_)
  );
  INV_X1 _38028_ (
    .A(_03726_),
    .ZN(_03727_)
  );
  AND2_X1 _38029_ (
    .A1(_03721_),
    .A2(_03726_),
    .ZN(_03728_)
  );
  INV_X1 _38030_ (
    .A(_03728_),
    .ZN(_03729_)
  );
  AND2_X1 _38031_ (
    .A1(_03720_),
    .A2(_03727_),
    .ZN(_03730_)
  );
  INV_X1 _38032_ (
    .A(_03730_),
    .ZN(_03731_)
  );
  AND2_X1 _38033_ (
    .A1(instr_jal),
    .A2(_03731_),
    .ZN(_03732_)
  );
  AND2_X1 _38034_ (
    .A1(_03729_),
    .A2(_03732_),
    .ZN(_03733_)
  );
  INV_X1 _38035_ (
    .A(_03733_),
    .ZN(_03734_)
  );
  AND2_X1 _38036_ (
    .A1(_03088_),
    .A2(_03704_),
    .ZN(_03735_)
  );
  INV_X1 _38037_ (
    .A(_03735_),
    .ZN(_03736_)
  );
  AND2_X1 _38038_ (
    .A1(_03087_),
    .A2(_03703_),
    .ZN(_03737_)
  );
  INV_X1 _38039_ (
    .A(_03737_),
    .ZN(_03738_)
  );
  AND2_X1 _38040_ (
    .A1(_21261_),
    .A2(_03738_),
    .ZN(_03739_)
  );
  AND2_X1 _38041_ (
    .A1(_03736_),
    .A2(_03739_),
    .ZN(_03740_)
  );
  INV_X1 _38042_ (
    .A(_03740_),
    .ZN(_03741_)
  );
  AND2_X1 _38043_ (
    .A1(decoder_trigger),
    .A2(_03741_),
    .ZN(_03742_)
  );
  AND2_X1 _38044_ (
    .A1(_03734_),
    .A2(_03742_),
    .ZN(_03743_)
  );
  INV_X1 _38045_ (
    .A(_03743_),
    .ZN(_03744_)
  );
  AND2_X1 _38046_ (
    .A1(_02470_),
    .A2(_03088_),
    .ZN(_03745_)
  );
  INV_X1 _38047_ (
    .A(_03745_),
    .ZN(_03746_)
  );
  AND2_X1 _38048_ (
    .A1(_03744_),
    .A2(_03746_),
    .ZN(_03747_)
  );
  INV_X1 _38049_ (
    .A(_03747_),
    .ZN(_03748_)
  );
  AND2_X1 _38050_ (
    .A1(_03719_),
    .A2(_03748_),
    .ZN(_03749_)
  );
  INV_X1 _38051_ (
    .A(_03749_),
    .ZN(_00195_)
  );
  AND2_X1 _38052_ (
    .A1(reg_next_pc[12]),
    .A2(_02928_),
    .ZN(_03750_)
  );
  INV_X1 _38053_ (
    .A(_03750_),
    .ZN(_03751_)
  );
  AND2_X1 _38054_ (
    .A1(decoded_imm_j[12]),
    .A2(_03103_),
    .ZN(_03752_)
  );
  INV_X1 _38055_ (
    .A(_03752_),
    .ZN(_03753_)
  );
  AND2_X1 _38056_ (
    .A1(_22016_),
    .A2(_03104_),
    .ZN(_03754_)
  );
  INV_X1 _38057_ (
    .A(_03754_),
    .ZN(_03755_)
  );
  AND2_X1 _38058_ (
    .A1(_03753_),
    .A2(_03755_),
    .ZN(_03756_)
  );
  INV_X1 _38059_ (
    .A(_03756_),
    .ZN(_03757_)
  );
  AND2_X1 _38060_ (
    .A1(_03720_),
    .A2(_03723_),
    .ZN(_03758_)
  );
  INV_X1 _38061_ (
    .A(_03758_),
    .ZN(_03759_)
  );
  AND2_X1 _38062_ (
    .A1(_03721_),
    .A2(_03725_),
    .ZN(_03760_)
  );
  INV_X1 _38063_ (
    .A(_03760_),
    .ZN(_03761_)
  );
  AND2_X1 _38064_ (
    .A1(_03725_),
    .A2(_03759_),
    .ZN(_03762_)
  );
  AND2_X1 _38065_ (
    .A1(_03723_),
    .A2(_03761_),
    .ZN(_03763_)
  );
  AND2_X1 _38066_ (
    .A1(_03757_),
    .A2(_03763_),
    .ZN(_03764_)
  );
  INV_X1 _38067_ (
    .A(_03764_),
    .ZN(_03765_)
  );
  AND2_X1 _38068_ (
    .A1(_03756_),
    .A2(_03762_),
    .ZN(_03766_)
  );
  INV_X1 _38069_ (
    .A(_03766_),
    .ZN(_03767_)
  );
  AND2_X1 _38070_ (
    .A1(instr_jal),
    .A2(_03767_),
    .ZN(_03768_)
  );
  AND2_X1 _38071_ (
    .A1(_03765_),
    .A2(_03768_),
    .ZN(_03769_)
  );
  INV_X1 _38072_ (
    .A(_03769_),
    .ZN(_03770_)
  );
  AND2_X1 _38073_ (
    .A1(_03102_),
    .A2(_03737_),
    .ZN(_03771_)
  );
  INV_X1 _38074_ (
    .A(_03771_),
    .ZN(_03772_)
  );
  AND2_X1 _38075_ (
    .A1(_03104_),
    .A2(_03738_),
    .ZN(_03773_)
  );
  INV_X1 _38076_ (
    .A(_03773_),
    .ZN(_03774_)
  );
  AND2_X1 _38077_ (
    .A1(_03772_),
    .A2(_03774_),
    .ZN(_03775_)
  );
  AND2_X1 _38078_ (
    .A1(_21261_),
    .A2(_03775_),
    .ZN(_03776_)
  );
  INV_X1 _38079_ (
    .A(_03776_),
    .ZN(_03777_)
  );
  AND2_X1 _38080_ (
    .A1(decoder_trigger),
    .A2(_03777_),
    .ZN(_03778_)
  );
  AND2_X1 _38081_ (
    .A1(_03770_),
    .A2(_03778_),
    .ZN(_03779_)
  );
  INV_X1 _38082_ (
    .A(_03779_),
    .ZN(_03780_)
  );
  AND2_X1 _38083_ (
    .A1(_02470_),
    .A2(_03104_),
    .ZN(_03781_)
  );
  INV_X1 _38084_ (
    .A(_03781_),
    .ZN(_03782_)
  );
  AND2_X1 _38085_ (
    .A1(_03780_),
    .A2(_03782_),
    .ZN(_03783_)
  );
  INV_X1 _38086_ (
    .A(_03783_),
    .ZN(_03784_)
  );
  AND2_X1 _38087_ (
    .A1(_03751_),
    .A2(_03784_),
    .ZN(_03785_)
  );
  INV_X1 _38088_ (
    .A(_03785_),
    .ZN(_00196_)
  );
  AND2_X1 _38089_ (
    .A1(reg_next_pc[13]),
    .A2(_02928_),
    .ZN(_03786_)
  );
  INV_X1 _38090_ (
    .A(_03786_),
    .ZN(_03787_)
  );
  AND2_X1 _38091_ (
    .A1(_03753_),
    .A2(_03767_),
    .ZN(_03788_)
  );
  INV_X1 _38092_ (
    .A(_03788_),
    .ZN(_03789_)
  );
  AND2_X1 _38093_ (
    .A1(decoded_imm_j[13]),
    .A2(_03119_),
    .ZN(_03790_)
  );
  INV_X1 _38094_ (
    .A(_03790_),
    .ZN(_03791_)
  );
  AND2_X1 _38095_ (
    .A1(_22017_),
    .A2(_03120_),
    .ZN(_03792_)
  );
  INV_X1 _38096_ (
    .A(_03792_),
    .ZN(_03793_)
  );
  AND2_X1 _38097_ (
    .A1(_03791_),
    .A2(_03793_),
    .ZN(_03794_)
  );
  INV_X1 _38098_ (
    .A(_03794_),
    .ZN(_03795_)
  );
  AND2_X1 _38099_ (
    .A1(_03789_),
    .A2(_03794_),
    .ZN(_03796_)
  );
  INV_X1 _38100_ (
    .A(_03796_),
    .ZN(_03797_)
  );
  AND2_X1 _38101_ (
    .A1(_03788_),
    .A2(_03795_),
    .ZN(_03798_)
  );
  INV_X1 _38102_ (
    .A(_03798_),
    .ZN(_03799_)
  );
  AND2_X1 _38103_ (
    .A1(instr_jal),
    .A2(_03799_),
    .ZN(_03800_)
  );
  AND2_X1 _38104_ (
    .A1(_03797_),
    .A2(_03800_),
    .ZN(_03801_)
  );
  INV_X1 _38105_ (
    .A(_03801_),
    .ZN(_03802_)
  );
  AND2_X1 _38106_ (
    .A1(_03120_),
    .A2(_03772_),
    .ZN(_03803_)
  );
  INV_X1 _38107_ (
    .A(_03803_),
    .ZN(_03804_)
  );
  AND2_X1 _38108_ (
    .A1(_03119_),
    .A2(_03771_),
    .ZN(_03805_)
  );
  INV_X1 _38109_ (
    .A(_03805_),
    .ZN(_03806_)
  );
  AND2_X1 _38110_ (
    .A1(_21261_),
    .A2(_03806_),
    .ZN(_03807_)
  );
  AND2_X1 _38111_ (
    .A1(_03804_),
    .A2(_03807_),
    .ZN(_03808_)
  );
  INV_X1 _38112_ (
    .A(_03808_),
    .ZN(_03809_)
  );
  AND2_X1 _38113_ (
    .A1(decoder_trigger),
    .A2(_03809_),
    .ZN(_03810_)
  );
  AND2_X1 _38114_ (
    .A1(_03802_),
    .A2(_03810_),
    .ZN(_03811_)
  );
  INV_X1 _38115_ (
    .A(_03811_),
    .ZN(_03812_)
  );
  AND2_X1 _38116_ (
    .A1(_02470_),
    .A2(_03120_),
    .ZN(_03813_)
  );
  INV_X1 _38117_ (
    .A(_03813_),
    .ZN(_03814_)
  );
  AND2_X1 _38118_ (
    .A1(_03812_),
    .A2(_03814_),
    .ZN(_03815_)
  );
  INV_X1 _38119_ (
    .A(_03815_),
    .ZN(_03816_)
  );
  AND2_X1 _38120_ (
    .A1(_03787_),
    .A2(_03816_),
    .ZN(_03817_)
  );
  INV_X1 _38121_ (
    .A(_03817_),
    .ZN(_00197_)
  );
  AND2_X1 _38122_ (
    .A1(reg_next_pc[14]),
    .A2(_02928_),
    .ZN(_03818_)
  );
  INV_X1 _38123_ (
    .A(_03818_),
    .ZN(_03819_)
  );
  AND2_X1 _38124_ (
    .A1(decoded_imm_j[14]),
    .A2(_03135_),
    .ZN(_03820_)
  );
  INV_X1 _38125_ (
    .A(_03820_),
    .ZN(_03821_)
  );
  AND2_X1 _38126_ (
    .A1(_22018_),
    .A2(_03136_),
    .ZN(_03822_)
  );
  INV_X1 _38127_ (
    .A(_03822_),
    .ZN(_03823_)
  );
  AND2_X1 _38128_ (
    .A1(_03821_),
    .A2(_03823_),
    .ZN(_03824_)
  );
  INV_X1 _38129_ (
    .A(_03824_),
    .ZN(_03825_)
  );
  AND2_X1 _38130_ (
    .A1(_03788_),
    .A2(_03791_),
    .ZN(_03826_)
  );
  INV_X1 _38131_ (
    .A(_03826_),
    .ZN(_03827_)
  );
  AND2_X1 _38132_ (
    .A1(_03789_),
    .A2(_03793_),
    .ZN(_03828_)
  );
  INV_X1 _38133_ (
    .A(_03828_),
    .ZN(_03829_)
  );
  AND2_X1 _38134_ (
    .A1(_03793_),
    .A2(_03827_),
    .ZN(_03830_)
  );
  AND2_X1 _38135_ (
    .A1(_03791_),
    .A2(_03829_),
    .ZN(_03831_)
  );
  AND2_X1 _38136_ (
    .A1(_03825_),
    .A2(_03831_),
    .ZN(_03832_)
  );
  INV_X1 _38137_ (
    .A(_03832_),
    .ZN(_03833_)
  );
  AND2_X1 _38138_ (
    .A1(_03824_),
    .A2(_03830_),
    .ZN(_03834_)
  );
  INV_X1 _38139_ (
    .A(_03834_),
    .ZN(_03835_)
  );
  AND2_X1 _38140_ (
    .A1(instr_jal),
    .A2(_03835_),
    .ZN(_03836_)
  );
  AND2_X1 _38141_ (
    .A1(_03833_),
    .A2(_03836_),
    .ZN(_03837_)
  );
  INV_X1 _38142_ (
    .A(_03837_),
    .ZN(_03838_)
  );
  AND2_X1 _38143_ (
    .A1(_03134_),
    .A2(_03805_),
    .ZN(_03839_)
  );
  INV_X1 _38144_ (
    .A(_03839_),
    .ZN(_03840_)
  );
  AND2_X1 _38145_ (
    .A1(_03136_),
    .A2(_03806_),
    .ZN(_03841_)
  );
  INV_X1 _38146_ (
    .A(_03841_),
    .ZN(_03842_)
  );
  AND2_X1 _38147_ (
    .A1(_03840_),
    .A2(_03842_),
    .ZN(_03843_)
  );
  AND2_X1 _38148_ (
    .A1(_21261_),
    .A2(_03843_),
    .ZN(_03844_)
  );
  INV_X1 _38149_ (
    .A(_03844_),
    .ZN(_03845_)
  );
  AND2_X1 _38150_ (
    .A1(decoder_trigger),
    .A2(_03845_),
    .ZN(_03846_)
  );
  AND2_X1 _38151_ (
    .A1(_03838_),
    .A2(_03846_),
    .ZN(_03847_)
  );
  INV_X1 _38152_ (
    .A(_03847_),
    .ZN(_03848_)
  );
  AND2_X1 _38153_ (
    .A1(_02470_),
    .A2(_03136_),
    .ZN(_03849_)
  );
  INV_X1 _38154_ (
    .A(_03849_),
    .ZN(_03850_)
  );
  AND2_X1 _38155_ (
    .A1(_03848_),
    .A2(_03850_),
    .ZN(_03851_)
  );
  INV_X1 _38156_ (
    .A(_03851_),
    .ZN(_03852_)
  );
  AND2_X1 _38157_ (
    .A1(_03819_),
    .A2(_03852_),
    .ZN(_03853_)
  );
  INV_X1 _38158_ (
    .A(_03853_),
    .ZN(_00198_)
  );
  AND2_X1 _38159_ (
    .A1(reg_next_pc[15]),
    .A2(_02928_),
    .ZN(_03854_)
  );
  INV_X1 _38160_ (
    .A(_03854_),
    .ZN(_03855_)
  );
  AND2_X1 _38161_ (
    .A1(_03821_),
    .A2(_03835_),
    .ZN(_03856_)
  );
  INV_X1 _38162_ (
    .A(_03856_),
    .ZN(_03857_)
  );
  AND2_X1 _38163_ (
    .A1(decoded_rs1[0]),
    .A2(_03151_),
    .ZN(_03858_)
  );
  INV_X1 _38164_ (
    .A(_03858_),
    .ZN(_03859_)
  );
  AND2_X1 _38165_ (
    .A1(_22021_),
    .A2(_03152_),
    .ZN(_03860_)
  );
  INV_X1 _38166_ (
    .A(_03860_),
    .ZN(_03861_)
  );
  AND2_X1 _38167_ (
    .A1(_03859_),
    .A2(_03861_),
    .ZN(_03862_)
  );
  INV_X1 _38168_ (
    .A(_03862_),
    .ZN(_03863_)
  );
  AND2_X1 _38169_ (
    .A1(_03857_),
    .A2(_03862_),
    .ZN(_03864_)
  );
  INV_X1 _38170_ (
    .A(_03864_),
    .ZN(_03865_)
  );
  AND2_X1 _38171_ (
    .A1(_03856_),
    .A2(_03863_),
    .ZN(_03866_)
  );
  INV_X1 _38172_ (
    .A(_03866_),
    .ZN(_03867_)
  );
  AND2_X1 _38173_ (
    .A1(instr_jal),
    .A2(_03867_),
    .ZN(_03868_)
  );
  AND2_X1 _38174_ (
    .A1(_03865_),
    .A2(_03868_),
    .ZN(_03869_)
  );
  INV_X1 _38175_ (
    .A(_03869_),
    .ZN(_03870_)
  );
  AND2_X1 _38176_ (
    .A1(_03152_),
    .A2(_03840_),
    .ZN(_03871_)
  );
  INV_X1 _38177_ (
    .A(_03871_),
    .ZN(_03872_)
  );
  AND2_X1 _38178_ (
    .A1(_03151_),
    .A2(_03839_),
    .ZN(_03873_)
  );
  INV_X1 _38179_ (
    .A(_03873_),
    .ZN(_03874_)
  );
  AND2_X1 _38180_ (
    .A1(_21261_),
    .A2(_03874_),
    .ZN(_03875_)
  );
  AND2_X1 _38181_ (
    .A1(_03872_),
    .A2(_03875_),
    .ZN(_03876_)
  );
  INV_X1 _38182_ (
    .A(_03876_),
    .ZN(_03877_)
  );
  AND2_X1 _38183_ (
    .A1(decoder_trigger),
    .A2(_03877_),
    .ZN(_03878_)
  );
  AND2_X1 _38184_ (
    .A1(_03870_),
    .A2(_03878_),
    .ZN(_03879_)
  );
  INV_X1 _38185_ (
    .A(_03879_),
    .ZN(_03880_)
  );
  AND2_X1 _38186_ (
    .A1(_02470_),
    .A2(_03152_),
    .ZN(_03881_)
  );
  INV_X1 _38187_ (
    .A(_03881_),
    .ZN(_03882_)
  );
  AND2_X1 _38188_ (
    .A1(_03880_),
    .A2(_03882_),
    .ZN(_03883_)
  );
  INV_X1 _38189_ (
    .A(_03883_),
    .ZN(_03884_)
  );
  AND2_X1 _38190_ (
    .A1(_03855_),
    .A2(_03884_),
    .ZN(_03885_)
  );
  INV_X1 _38191_ (
    .A(_03885_),
    .ZN(_00199_)
  );
  AND2_X1 _38192_ (
    .A1(reg_next_pc[16]),
    .A2(_02928_),
    .ZN(_03886_)
  );
  INV_X1 _38193_ (
    .A(_03886_),
    .ZN(_03887_)
  );
  AND2_X1 _38194_ (
    .A1(decoded_rs1[1]),
    .A2(_03167_),
    .ZN(_03888_)
  );
  INV_X1 _38195_ (
    .A(_03888_),
    .ZN(_03889_)
  );
  AND2_X1 _38196_ (
    .A1(_22022_),
    .A2(_03168_),
    .ZN(_03890_)
  );
  INV_X1 _38197_ (
    .A(_03890_),
    .ZN(_03891_)
  );
  AND2_X1 _38198_ (
    .A1(_03889_),
    .A2(_03891_),
    .ZN(_03892_)
  );
  INV_X1 _38199_ (
    .A(_03892_),
    .ZN(_03893_)
  );
  AND2_X1 _38200_ (
    .A1(_03856_),
    .A2(_03859_),
    .ZN(_03894_)
  );
  INV_X1 _38201_ (
    .A(_03894_),
    .ZN(_03895_)
  );
  AND2_X1 _38202_ (
    .A1(_03857_),
    .A2(_03861_),
    .ZN(_03896_)
  );
  INV_X1 _38203_ (
    .A(_03896_),
    .ZN(_03897_)
  );
  AND2_X1 _38204_ (
    .A1(_03861_),
    .A2(_03895_),
    .ZN(_03898_)
  );
  AND2_X1 _38205_ (
    .A1(_03859_),
    .A2(_03897_),
    .ZN(_03899_)
  );
  AND2_X1 _38206_ (
    .A1(_03893_),
    .A2(_03899_),
    .ZN(_03900_)
  );
  INV_X1 _38207_ (
    .A(_03900_),
    .ZN(_03901_)
  );
  AND2_X1 _38208_ (
    .A1(_03892_),
    .A2(_03898_),
    .ZN(_03902_)
  );
  INV_X1 _38209_ (
    .A(_03902_),
    .ZN(_03903_)
  );
  AND2_X1 _38210_ (
    .A1(instr_jal),
    .A2(_03903_),
    .ZN(_03904_)
  );
  AND2_X1 _38211_ (
    .A1(_03901_),
    .A2(_03904_),
    .ZN(_03905_)
  );
  INV_X1 _38212_ (
    .A(_03905_),
    .ZN(_03906_)
  );
  AND2_X1 _38213_ (
    .A1(_03166_),
    .A2(_03873_),
    .ZN(_03907_)
  );
  INV_X1 _38214_ (
    .A(_03907_),
    .ZN(_03908_)
  );
  AND2_X1 _38215_ (
    .A1(_03168_),
    .A2(_03874_),
    .ZN(_03909_)
  );
  INV_X1 _38216_ (
    .A(_03909_),
    .ZN(_03910_)
  );
  AND2_X1 _38217_ (
    .A1(_03908_),
    .A2(_03910_),
    .ZN(_03911_)
  );
  AND2_X1 _38218_ (
    .A1(_21261_),
    .A2(_03911_),
    .ZN(_03912_)
  );
  INV_X1 _38219_ (
    .A(_03912_),
    .ZN(_03913_)
  );
  AND2_X1 _38220_ (
    .A1(decoder_trigger),
    .A2(_03913_),
    .ZN(_03914_)
  );
  AND2_X1 _38221_ (
    .A1(_03906_),
    .A2(_03914_),
    .ZN(_03915_)
  );
  INV_X1 _38222_ (
    .A(_03915_),
    .ZN(_03916_)
  );
  AND2_X1 _38223_ (
    .A1(_02470_),
    .A2(_03168_),
    .ZN(_03917_)
  );
  INV_X1 _38224_ (
    .A(_03917_),
    .ZN(_03918_)
  );
  AND2_X1 _38225_ (
    .A1(_03916_),
    .A2(_03918_),
    .ZN(_03919_)
  );
  INV_X1 _38226_ (
    .A(_03919_),
    .ZN(_03920_)
  );
  AND2_X1 _38227_ (
    .A1(_03887_),
    .A2(_03920_),
    .ZN(_03921_)
  );
  INV_X1 _38228_ (
    .A(_03921_),
    .ZN(_00200_)
  );
  AND2_X1 _38229_ (
    .A1(reg_next_pc[17]),
    .A2(_02928_),
    .ZN(_03922_)
  );
  INV_X1 _38230_ (
    .A(_03922_),
    .ZN(_03923_)
  );
  AND2_X1 _38231_ (
    .A1(_03889_),
    .A2(_03903_),
    .ZN(_03924_)
  );
  INV_X1 _38232_ (
    .A(_03924_),
    .ZN(_03925_)
  );
  AND2_X1 _38233_ (
    .A1(decoded_rs1[2]),
    .A2(_03183_),
    .ZN(_03926_)
  );
  INV_X1 _38234_ (
    .A(_03926_),
    .ZN(_03927_)
  );
  AND2_X1 _38235_ (
    .A1(_22023_),
    .A2(_03184_),
    .ZN(_03928_)
  );
  INV_X1 _38236_ (
    .A(_03928_),
    .ZN(_03929_)
  );
  AND2_X1 _38237_ (
    .A1(_03927_),
    .A2(_03929_),
    .ZN(_03930_)
  );
  INV_X1 _38238_ (
    .A(_03930_),
    .ZN(_03931_)
  );
  AND2_X1 _38239_ (
    .A1(_03925_),
    .A2(_03930_),
    .ZN(_03932_)
  );
  INV_X1 _38240_ (
    .A(_03932_),
    .ZN(_03933_)
  );
  AND2_X1 _38241_ (
    .A1(_03924_),
    .A2(_03931_),
    .ZN(_03934_)
  );
  INV_X1 _38242_ (
    .A(_03934_),
    .ZN(_03935_)
  );
  AND2_X1 _38243_ (
    .A1(instr_jal),
    .A2(_03935_),
    .ZN(_03936_)
  );
  AND2_X1 _38244_ (
    .A1(_03933_),
    .A2(_03936_),
    .ZN(_03937_)
  );
  INV_X1 _38245_ (
    .A(_03937_),
    .ZN(_03938_)
  );
  AND2_X1 _38246_ (
    .A1(_03183_),
    .A2(_03907_),
    .ZN(_03939_)
  );
  INV_X1 _38247_ (
    .A(_03939_),
    .ZN(_03940_)
  );
  AND2_X1 _38248_ (
    .A1(_03184_),
    .A2(_03908_),
    .ZN(_03941_)
  );
  INV_X1 _38249_ (
    .A(_03941_),
    .ZN(_03942_)
  );
  AND2_X1 _38250_ (
    .A1(_03940_),
    .A2(_03942_),
    .ZN(_03943_)
  );
  AND2_X1 _38251_ (
    .A1(_21261_),
    .A2(_03943_),
    .ZN(_03944_)
  );
  INV_X1 _38252_ (
    .A(_03944_),
    .ZN(_03945_)
  );
  AND2_X1 _38253_ (
    .A1(decoder_trigger),
    .A2(_03945_),
    .ZN(_03946_)
  );
  AND2_X1 _38254_ (
    .A1(_03938_),
    .A2(_03946_),
    .ZN(_03947_)
  );
  INV_X1 _38255_ (
    .A(_03947_),
    .ZN(_03948_)
  );
  AND2_X1 _38256_ (
    .A1(_02470_),
    .A2(_03184_),
    .ZN(_03949_)
  );
  INV_X1 _38257_ (
    .A(_03949_),
    .ZN(_03950_)
  );
  AND2_X1 _38258_ (
    .A1(_03948_),
    .A2(_03950_),
    .ZN(_03951_)
  );
  INV_X1 _38259_ (
    .A(_03951_),
    .ZN(_03952_)
  );
  AND2_X1 _38260_ (
    .A1(_03923_),
    .A2(_03952_),
    .ZN(_03953_)
  );
  INV_X1 _38261_ (
    .A(_03953_),
    .ZN(_00201_)
  );
  AND2_X1 _38262_ (
    .A1(reg_next_pc[18]),
    .A2(_02928_),
    .ZN(_03954_)
  );
  INV_X1 _38263_ (
    .A(_03954_),
    .ZN(_03955_)
  );
  AND2_X1 _38264_ (
    .A1(decoded_imm_j[18]),
    .A2(_03199_),
    .ZN(_03956_)
  );
  INV_X1 _38265_ (
    .A(_03956_),
    .ZN(_03957_)
  );
  AND2_X1 _38266_ (
    .A1(_22019_),
    .A2(_03200_),
    .ZN(_03958_)
  );
  INV_X1 _38267_ (
    .A(_03958_),
    .ZN(_03959_)
  );
  AND2_X1 _38268_ (
    .A1(_03957_),
    .A2(_03959_),
    .ZN(_03960_)
  );
  INV_X1 _38269_ (
    .A(_03960_),
    .ZN(_03961_)
  );
  AND2_X1 _38270_ (
    .A1(_03924_),
    .A2(_03927_),
    .ZN(_03962_)
  );
  INV_X1 _38271_ (
    .A(_03962_),
    .ZN(_03963_)
  );
  AND2_X1 _38272_ (
    .A1(_03925_),
    .A2(_03929_),
    .ZN(_03964_)
  );
  INV_X1 _38273_ (
    .A(_03964_),
    .ZN(_03965_)
  );
  AND2_X1 _38274_ (
    .A1(_03929_),
    .A2(_03963_),
    .ZN(_03966_)
  );
  AND2_X1 _38275_ (
    .A1(_03927_),
    .A2(_03965_),
    .ZN(_03967_)
  );
  AND2_X1 _38276_ (
    .A1(_03961_),
    .A2(_03967_),
    .ZN(_03968_)
  );
  INV_X1 _38277_ (
    .A(_03968_),
    .ZN(_03969_)
  );
  AND2_X1 _38278_ (
    .A1(_03960_),
    .A2(_03966_),
    .ZN(_03970_)
  );
  INV_X1 _38279_ (
    .A(_03970_),
    .ZN(_03971_)
  );
  AND2_X1 _38280_ (
    .A1(instr_jal),
    .A2(_03971_),
    .ZN(_03972_)
  );
  AND2_X1 _38281_ (
    .A1(_03969_),
    .A2(_03972_),
    .ZN(_03973_)
  );
  INV_X1 _38282_ (
    .A(_03973_),
    .ZN(_03974_)
  );
  AND2_X1 _38283_ (
    .A1(_03198_),
    .A2(_03939_),
    .ZN(_03975_)
  );
  INV_X1 _38284_ (
    .A(_03975_),
    .ZN(_03976_)
  );
  AND2_X1 _38285_ (
    .A1(_03200_),
    .A2(_03940_),
    .ZN(_03977_)
  );
  INV_X1 _38286_ (
    .A(_03977_),
    .ZN(_03978_)
  );
  AND2_X1 _38287_ (
    .A1(_03976_),
    .A2(_03978_),
    .ZN(_03979_)
  );
  AND2_X1 _38288_ (
    .A1(_21261_),
    .A2(_03979_),
    .ZN(_03980_)
  );
  INV_X1 _38289_ (
    .A(_03980_),
    .ZN(_03981_)
  );
  AND2_X1 _38290_ (
    .A1(decoder_trigger),
    .A2(_03981_),
    .ZN(_03982_)
  );
  AND2_X1 _38291_ (
    .A1(_03974_),
    .A2(_03982_),
    .ZN(_03983_)
  );
  INV_X1 _38292_ (
    .A(_03983_),
    .ZN(_03984_)
  );
  AND2_X1 _38293_ (
    .A1(_02470_),
    .A2(_03200_),
    .ZN(_03985_)
  );
  INV_X1 _38294_ (
    .A(_03985_),
    .ZN(_03986_)
  );
  AND2_X1 _38295_ (
    .A1(_03984_),
    .A2(_03986_),
    .ZN(_03987_)
  );
  INV_X1 _38296_ (
    .A(_03987_),
    .ZN(_03988_)
  );
  AND2_X1 _38297_ (
    .A1(_03955_),
    .A2(_03988_),
    .ZN(_03989_)
  );
  INV_X1 _38298_ (
    .A(_03989_),
    .ZN(_00202_)
  );
  AND2_X1 _38299_ (
    .A1(reg_next_pc[19]),
    .A2(_02928_),
    .ZN(_03990_)
  );
  INV_X1 _38300_ (
    .A(_03990_),
    .ZN(_03991_)
  );
  AND2_X1 _38301_ (
    .A1(_03957_),
    .A2(_03971_),
    .ZN(_03992_)
  );
  INV_X1 _38302_ (
    .A(_03992_),
    .ZN(_03993_)
  );
  AND2_X1 _38303_ (
    .A1(decoded_imm_j[19]),
    .A2(_03215_),
    .ZN(_03994_)
  );
  INV_X1 _38304_ (
    .A(_03994_),
    .ZN(_03995_)
  );
  AND2_X1 _38305_ (
    .A1(_22020_),
    .A2(_03216_),
    .ZN(_03996_)
  );
  INV_X1 _38306_ (
    .A(_03996_),
    .ZN(_03997_)
  );
  AND2_X1 _38307_ (
    .A1(_03995_),
    .A2(_03997_),
    .ZN(_03998_)
  );
  INV_X1 _38308_ (
    .A(_03998_),
    .ZN(_03999_)
  );
  AND2_X1 _38309_ (
    .A1(_03993_),
    .A2(_03998_),
    .ZN(_04000_)
  );
  INV_X1 _38310_ (
    .A(_04000_),
    .ZN(_04001_)
  );
  AND2_X1 _38311_ (
    .A1(_03992_),
    .A2(_03999_),
    .ZN(_04002_)
  );
  INV_X1 _38312_ (
    .A(_04002_),
    .ZN(_04003_)
  );
  AND2_X1 _38313_ (
    .A1(instr_jal),
    .A2(_04003_),
    .ZN(_04004_)
  );
  AND2_X1 _38314_ (
    .A1(_04001_),
    .A2(_04004_),
    .ZN(_04005_)
  );
  INV_X1 _38315_ (
    .A(_04005_),
    .ZN(_04006_)
  );
  AND2_X1 _38316_ (
    .A1(_03215_),
    .A2(_03975_),
    .ZN(_04007_)
  );
  INV_X1 _38317_ (
    .A(_04007_),
    .ZN(_04008_)
  );
  AND2_X1 _38318_ (
    .A1(_03216_),
    .A2(_03976_),
    .ZN(_04009_)
  );
  INV_X1 _38319_ (
    .A(_04009_),
    .ZN(_04010_)
  );
  AND2_X1 _38320_ (
    .A1(_04008_),
    .A2(_04010_),
    .ZN(_04011_)
  );
  AND2_X1 _38321_ (
    .A1(_21261_),
    .A2(_04011_),
    .ZN(_04012_)
  );
  INV_X1 _38322_ (
    .A(_04012_),
    .ZN(_04013_)
  );
  AND2_X1 _38323_ (
    .A1(decoder_trigger),
    .A2(_04013_),
    .ZN(_04014_)
  );
  AND2_X1 _38324_ (
    .A1(_04006_),
    .A2(_04014_),
    .ZN(_04015_)
  );
  INV_X1 _38325_ (
    .A(_04015_),
    .ZN(_04016_)
  );
  AND2_X1 _38326_ (
    .A1(_02470_),
    .A2(_03216_),
    .ZN(_04017_)
  );
  INV_X1 _38327_ (
    .A(_04017_),
    .ZN(_04018_)
  );
  AND2_X1 _38328_ (
    .A1(_04016_),
    .A2(_04018_),
    .ZN(_04019_)
  );
  INV_X1 _38329_ (
    .A(_04019_),
    .ZN(_04020_)
  );
  AND2_X1 _38330_ (
    .A1(_03991_),
    .A2(_04020_),
    .ZN(_04021_)
  );
  INV_X1 _38331_ (
    .A(_04021_),
    .ZN(_00203_)
  );
  AND2_X1 _38332_ (
    .A1(reg_next_pc[20]),
    .A2(_02928_),
    .ZN(_04022_)
  );
  INV_X1 _38333_ (
    .A(_04022_),
    .ZN(_04023_)
  );
  AND2_X1 _38334_ (
    .A1(decoded_imm_j[30]),
    .A2(_03231_),
    .ZN(_04024_)
  );
  INV_X1 _38335_ (
    .A(_04024_),
    .ZN(_04025_)
  );
  AND2_X1 _38336_ (
    .A1(_22014_),
    .A2(_03232_),
    .ZN(_04026_)
  );
  INV_X1 _38337_ (
    .A(_04026_),
    .ZN(_04027_)
  );
  AND2_X1 _38338_ (
    .A1(_04025_),
    .A2(_04027_),
    .ZN(_04028_)
  );
  INV_X1 _38339_ (
    .A(_04028_),
    .ZN(_04029_)
  );
  AND2_X1 _38340_ (
    .A1(_03992_),
    .A2(_03995_),
    .ZN(_04030_)
  );
  INV_X1 _38341_ (
    .A(_04030_),
    .ZN(_04031_)
  );
  AND2_X1 _38342_ (
    .A1(_03993_),
    .A2(_03997_),
    .ZN(_04032_)
  );
  INV_X1 _38343_ (
    .A(_04032_),
    .ZN(_04033_)
  );
  AND2_X1 _38344_ (
    .A1(_03997_),
    .A2(_04031_),
    .ZN(_04034_)
  );
  AND2_X1 _38345_ (
    .A1(_03995_),
    .A2(_04033_),
    .ZN(_04035_)
  );
  AND2_X1 _38346_ (
    .A1(_04029_),
    .A2(_04035_),
    .ZN(_04036_)
  );
  INV_X1 _38347_ (
    .A(_04036_),
    .ZN(_04037_)
  );
  AND2_X1 _38348_ (
    .A1(_04028_),
    .A2(_04034_),
    .ZN(_04038_)
  );
  INV_X1 _38349_ (
    .A(_04038_),
    .ZN(_04039_)
  );
  AND2_X1 _38350_ (
    .A1(instr_jal),
    .A2(_04039_),
    .ZN(_04040_)
  );
  AND2_X1 _38351_ (
    .A1(_04037_),
    .A2(_04040_),
    .ZN(_04041_)
  );
  INV_X1 _38352_ (
    .A(_04041_),
    .ZN(_04042_)
  );
  AND2_X1 _38353_ (
    .A1(_03230_),
    .A2(_04007_),
    .ZN(_04043_)
  );
  INV_X1 _38354_ (
    .A(_04043_),
    .ZN(_04044_)
  );
  AND2_X1 _38355_ (
    .A1(_03232_),
    .A2(_04008_),
    .ZN(_04045_)
  );
  INV_X1 _38356_ (
    .A(_04045_),
    .ZN(_04046_)
  );
  AND2_X1 _38357_ (
    .A1(_04044_),
    .A2(_04046_),
    .ZN(_04047_)
  );
  AND2_X1 _38358_ (
    .A1(_21261_),
    .A2(_04047_),
    .ZN(_04048_)
  );
  INV_X1 _38359_ (
    .A(_04048_),
    .ZN(_04049_)
  );
  AND2_X1 _38360_ (
    .A1(decoder_trigger),
    .A2(_04049_),
    .ZN(_04050_)
  );
  AND2_X1 _38361_ (
    .A1(_04042_),
    .A2(_04050_),
    .ZN(_04051_)
  );
  INV_X1 _38362_ (
    .A(_04051_),
    .ZN(_04052_)
  );
  AND2_X1 _38363_ (
    .A1(_02470_),
    .A2(_03232_),
    .ZN(_04053_)
  );
  INV_X1 _38364_ (
    .A(_04053_),
    .ZN(_04054_)
  );
  AND2_X1 _38365_ (
    .A1(_04052_),
    .A2(_04054_),
    .ZN(_04055_)
  );
  INV_X1 _38366_ (
    .A(_04055_),
    .ZN(_04056_)
  );
  AND2_X1 _38367_ (
    .A1(_04023_),
    .A2(_04056_),
    .ZN(_04057_)
  );
  INV_X1 _38368_ (
    .A(_04057_),
    .ZN(_00204_)
  );
  AND2_X1 _38369_ (
    .A1(_04025_),
    .A2(_04039_),
    .ZN(_04058_)
  );
  INV_X1 _38370_ (
    .A(_04058_),
    .ZN(_04059_)
  );
  AND2_X1 _38371_ (
    .A1(decoded_imm_j[30]),
    .A2(_03247_),
    .ZN(_04060_)
  );
  INV_X1 _38372_ (
    .A(_04060_),
    .ZN(_04061_)
  );
  AND2_X1 _38373_ (
    .A1(_22014_),
    .A2(_03248_),
    .ZN(_04062_)
  );
  INV_X1 _38374_ (
    .A(_04062_),
    .ZN(_04063_)
  );
  AND2_X1 _38375_ (
    .A1(_04061_),
    .A2(_04063_),
    .ZN(_04064_)
  );
  INV_X1 _38376_ (
    .A(_04064_),
    .ZN(_04065_)
  );
  AND2_X1 _38377_ (
    .A1(_04059_),
    .A2(_04064_),
    .ZN(_04066_)
  );
  INV_X1 _38378_ (
    .A(_04066_),
    .ZN(_04067_)
  );
  AND2_X1 _38379_ (
    .A1(_04058_),
    .A2(_04065_),
    .ZN(_04068_)
  );
  INV_X1 _38380_ (
    .A(_04068_),
    .ZN(_04069_)
  );
  AND2_X1 _38381_ (
    .A1(instr_jal),
    .A2(_04069_),
    .ZN(_04070_)
  );
  AND2_X1 _38382_ (
    .A1(_04067_),
    .A2(_04070_),
    .ZN(_04071_)
  );
  INV_X1 _38383_ (
    .A(_04071_),
    .ZN(_04072_)
  );
  AND2_X1 _38384_ (
    .A1(_03248_),
    .A2(_04044_),
    .ZN(_04073_)
  );
  INV_X1 _38385_ (
    .A(_04073_),
    .ZN(_04074_)
  );
  AND2_X1 _38386_ (
    .A1(_03247_),
    .A2(_04043_),
    .ZN(_04075_)
  );
  INV_X1 _38387_ (
    .A(_04075_),
    .ZN(_04076_)
  );
  AND2_X1 _38388_ (
    .A1(_21261_),
    .A2(_04076_),
    .ZN(_04077_)
  );
  AND2_X1 _38389_ (
    .A1(_04074_),
    .A2(_04077_),
    .ZN(_04078_)
  );
  INV_X1 _38390_ (
    .A(_04078_),
    .ZN(_04079_)
  );
  AND2_X1 _38391_ (
    .A1(decoder_trigger),
    .A2(_04079_),
    .ZN(_04080_)
  );
  AND2_X1 _38392_ (
    .A1(_04072_),
    .A2(_04080_),
    .ZN(_04081_)
  );
  INV_X1 _38393_ (
    .A(_04081_),
    .ZN(_04082_)
  );
  AND2_X1 _38394_ (
    .A1(_02470_),
    .A2(_03248_),
    .ZN(_04083_)
  );
  INV_X1 _38395_ (
    .A(_04083_),
    .ZN(_04084_)
  );
  AND2_X1 _38396_ (
    .A1(_04082_),
    .A2(_04084_),
    .ZN(_04085_)
  );
  INV_X1 _38397_ (
    .A(_04085_),
    .ZN(_04086_)
  );
  AND2_X1 _38398_ (
    .A1(reg_next_pc[21]),
    .A2(_02928_),
    .ZN(_04087_)
  );
  INV_X1 _38399_ (
    .A(_04087_),
    .ZN(_04088_)
  );
  AND2_X1 _38400_ (
    .A1(_04086_),
    .A2(_04088_),
    .ZN(_04089_)
  );
  INV_X1 _38401_ (
    .A(_04089_),
    .ZN(_00205_)
  );
  AND2_X1 _38402_ (
    .A1(reg_next_pc[22]),
    .A2(_02928_),
    .ZN(_04090_)
  );
  INV_X1 _38403_ (
    .A(_04090_),
    .ZN(_04091_)
  );
  AND2_X1 _38404_ (
    .A1(_04038_),
    .A2(_04064_),
    .ZN(_04092_)
  );
  INV_X1 _38405_ (
    .A(_04092_),
    .ZN(_04093_)
  );
  AND2_X1 _38406_ (
    .A1(_04025_),
    .A2(_04061_),
    .ZN(_04094_)
  );
  AND2_X1 _38407_ (
    .A1(_04093_),
    .A2(_04094_),
    .ZN(_04095_)
  );
  INV_X1 _38408_ (
    .A(_04095_),
    .ZN(_04096_)
  );
  AND2_X1 _38409_ (
    .A1(decoded_imm_j[30]),
    .A2(_03263_),
    .ZN(_04097_)
  );
  INV_X1 _38410_ (
    .A(_04097_),
    .ZN(_04098_)
  );
  AND2_X1 _38411_ (
    .A1(_22014_),
    .A2(_03264_),
    .ZN(_04099_)
  );
  INV_X1 _38412_ (
    .A(_04099_),
    .ZN(_04100_)
  );
  AND2_X1 _38413_ (
    .A1(_04098_),
    .A2(_04100_),
    .ZN(_04101_)
  );
  INV_X1 _38414_ (
    .A(_04101_),
    .ZN(_04102_)
  );
  AND2_X1 _38415_ (
    .A1(_04095_),
    .A2(_04102_),
    .ZN(_04103_)
  );
  INV_X1 _38416_ (
    .A(_04103_),
    .ZN(_04104_)
  );
  AND2_X1 _38417_ (
    .A1(_04096_),
    .A2(_04101_),
    .ZN(_04105_)
  );
  INV_X1 _38418_ (
    .A(_04105_),
    .ZN(_04106_)
  );
  AND2_X1 _38419_ (
    .A1(instr_jal),
    .A2(_04104_),
    .ZN(_04107_)
  );
  AND2_X1 _38420_ (
    .A1(_04106_),
    .A2(_04107_),
    .ZN(_04108_)
  );
  INV_X1 _38421_ (
    .A(_04108_),
    .ZN(_04109_)
  );
  AND2_X1 _38422_ (
    .A1(_03262_),
    .A2(_04075_),
    .ZN(_04110_)
  );
  INV_X1 _38423_ (
    .A(_04110_),
    .ZN(_04111_)
  );
  AND2_X1 _38424_ (
    .A1(_03264_),
    .A2(_04076_),
    .ZN(_04112_)
  );
  INV_X1 _38425_ (
    .A(_04112_),
    .ZN(_04113_)
  );
  AND2_X1 _38426_ (
    .A1(_04111_),
    .A2(_04113_),
    .ZN(_04114_)
  );
  AND2_X1 _38427_ (
    .A1(_21261_),
    .A2(_04114_),
    .ZN(_04115_)
  );
  INV_X1 _38428_ (
    .A(_04115_),
    .ZN(_04116_)
  );
  AND2_X1 _38429_ (
    .A1(decoder_trigger),
    .A2(_04116_),
    .ZN(_04117_)
  );
  AND2_X1 _38430_ (
    .A1(_04109_),
    .A2(_04117_),
    .ZN(_04118_)
  );
  INV_X1 _38431_ (
    .A(_04118_),
    .ZN(_04119_)
  );
  AND2_X1 _38432_ (
    .A1(_02470_),
    .A2(_03264_),
    .ZN(_04120_)
  );
  INV_X1 _38433_ (
    .A(_04120_),
    .ZN(_04121_)
  );
  AND2_X1 _38434_ (
    .A1(_04119_),
    .A2(_04121_),
    .ZN(_04122_)
  );
  INV_X1 _38435_ (
    .A(_04122_),
    .ZN(_04123_)
  );
  AND2_X1 _38436_ (
    .A1(_04091_),
    .A2(_04123_),
    .ZN(_04124_)
  );
  INV_X1 _38437_ (
    .A(_04124_),
    .ZN(_00206_)
  );
  AND2_X1 _38438_ (
    .A1(_04098_),
    .A2(_04106_),
    .ZN(_04125_)
  );
  INV_X1 _38439_ (
    .A(_04125_),
    .ZN(_04126_)
  );
  AND2_X1 _38440_ (
    .A1(decoded_imm_j[30]),
    .A2(_03279_),
    .ZN(_04127_)
  );
  INV_X1 _38441_ (
    .A(_04127_),
    .ZN(_04128_)
  );
  AND2_X1 _38442_ (
    .A1(_22014_),
    .A2(_03280_),
    .ZN(_04129_)
  );
  INV_X1 _38443_ (
    .A(_04129_),
    .ZN(_04130_)
  );
  AND2_X1 _38444_ (
    .A1(_04128_),
    .A2(_04130_),
    .ZN(_04131_)
  );
  INV_X1 _38445_ (
    .A(_04131_),
    .ZN(_04132_)
  );
  AND2_X1 _38446_ (
    .A1(_04126_),
    .A2(_04131_),
    .ZN(_04133_)
  );
  INV_X1 _38447_ (
    .A(_04133_),
    .ZN(_04134_)
  );
  AND2_X1 _38448_ (
    .A1(_04125_),
    .A2(_04132_),
    .ZN(_04135_)
  );
  INV_X1 _38449_ (
    .A(_04135_),
    .ZN(_04136_)
  );
  AND2_X1 _38450_ (
    .A1(instr_jal),
    .A2(_04136_),
    .ZN(_04137_)
  );
  AND2_X1 _38451_ (
    .A1(_04134_),
    .A2(_04137_),
    .ZN(_04138_)
  );
  INV_X1 _38452_ (
    .A(_04138_),
    .ZN(_04139_)
  );
  AND2_X1 _38453_ (
    .A1(_03280_),
    .A2(_04111_),
    .ZN(_04140_)
  );
  INV_X1 _38454_ (
    .A(_04140_),
    .ZN(_04141_)
  );
  AND2_X1 _38455_ (
    .A1(_03279_),
    .A2(_04110_),
    .ZN(_04142_)
  );
  INV_X1 _38456_ (
    .A(_04142_),
    .ZN(_04143_)
  );
  AND2_X1 _38457_ (
    .A1(_21261_),
    .A2(_04143_),
    .ZN(_04144_)
  );
  AND2_X1 _38458_ (
    .A1(_04141_),
    .A2(_04144_),
    .ZN(_04145_)
  );
  INV_X1 _38459_ (
    .A(_04145_),
    .ZN(_04146_)
  );
  AND2_X1 _38460_ (
    .A1(decoder_trigger),
    .A2(_04146_),
    .ZN(_04147_)
  );
  AND2_X1 _38461_ (
    .A1(_04139_),
    .A2(_04147_),
    .ZN(_04148_)
  );
  INV_X1 _38462_ (
    .A(_04148_),
    .ZN(_04149_)
  );
  AND2_X1 _38463_ (
    .A1(_02470_),
    .A2(_03280_),
    .ZN(_04150_)
  );
  INV_X1 _38464_ (
    .A(_04150_),
    .ZN(_04151_)
  );
  AND2_X1 _38465_ (
    .A1(_04149_),
    .A2(_04151_),
    .ZN(_04152_)
  );
  INV_X1 _38466_ (
    .A(_04152_),
    .ZN(_04153_)
  );
  AND2_X1 _38467_ (
    .A1(reg_next_pc[23]),
    .A2(_02928_),
    .ZN(_04154_)
  );
  INV_X1 _38468_ (
    .A(_04154_),
    .ZN(_04155_)
  );
  AND2_X1 _38469_ (
    .A1(_04153_),
    .A2(_04155_),
    .ZN(_04156_)
  );
  INV_X1 _38470_ (
    .A(_04156_),
    .ZN(_00207_)
  );
  AND2_X1 _38471_ (
    .A1(reg_next_pc[24]),
    .A2(_02928_),
    .ZN(_04157_)
  );
  INV_X1 _38472_ (
    .A(_04157_),
    .ZN(_04158_)
  );
  AND2_X1 _38473_ (
    .A1(_04105_),
    .A2(_04131_),
    .ZN(_04159_)
  );
  INV_X1 _38474_ (
    .A(_04159_),
    .ZN(_04160_)
  );
  AND2_X1 _38475_ (
    .A1(_04098_),
    .A2(_04128_),
    .ZN(_04161_)
  );
  AND2_X1 _38476_ (
    .A1(_04160_),
    .A2(_04161_),
    .ZN(_04162_)
  );
  INV_X1 _38477_ (
    .A(_04162_),
    .ZN(_04163_)
  );
  AND2_X1 _38478_ (
    .A1(decoded_imm_j[30]),
    .A2(_03295_),
    .ZN(_04164_)
  );
  INV_X1 _38479_ (
    .A(_04164_),
    .ZN(_04165_)
  );
  AND2_X1 _38480_ (
    .A1(_22014_),
    .A2(_03296_),
    .ZN(_04166_)
  );
  INV_X1 _38481_ (
    .A(_04166_),
    .ZN(_04167_)
  );
  AND2_X1 _38482_ (
    .A1(_04165_),
    .A2(_04167_),
    .ZN(_04168_)
  );
  INV_X1 _38483_ (
    .A(_04168_),
    .ZN(_04169_)
  );
  AND2_X1 _38484_ (
    .A1(_04162_),
    .A2(_04169_),
    .ZN(_04170_)
  );
  INV_X1 _38485_ (
    .A(_04170_),
    .ZN(_04171_)
  );
  AND2_X1 _38486_ (
    .A1(_04163_),
    .A2(_04168_),
    .ZN(_04172_)
  );
  INV_X1 _38487_ (
    .A(_04172_),
    .ZN(_04173_)
  );
  AND2_X1 _38488_ (
    .A1(instr_jal),
    .A2(_04171_),
    .ZN(_04174_)
  );
  AND2_X1 _38489_ (
    .A1(_04173_),
    .A2(_04174_),
    .ZN(_04175_)
  );
  INV_X1 _38490_ (
    .A(_04175_),
    .ZN(_04176_)
  );
  AND2_X1 _38491_ (
    .A1(_03294_),
    .A2(_04142_),
    .ZN(_04177_)
  );
  INV_X1 _38492_ (
    .A(_04177_),
    .ZN(_04178_)
  );
  AND2_X1 _38493_ (
    .A1(_03296_),
    .A2(_04143_),
    .ZN(_04179_)
  );
  INV_X1 _38494_ (
    .A(_04179_),
    .ZN(_04180_)
  );
  AND2_X1 _38495_ (
    .A1(_04178_),
    .A2(_04180_),
    .ZN(_04181_)
  );
  AND2_X1 _38496_ (
    .A1(_21261_),
    .A2(_04181_),
    .ZN(_04182_)
  );
  INV_X1 _38497_ (
    .A(_04182_),
    .ZN(_04183_)
  );
  AND2_X1 _38498_ (
    .A1(decoder_trigger),
    .A2(_04183_),
    .ZN(_04184_)
  );
  AND2_X1 _38499_ (
    .A1(_04176_),
    .A2(_04184_),
    .ZN(_04185_)
  );
  INV_X1 _38500_ (
    .A(_04185_),
    .ZN(_04186_)
  );
  AND2_X1 _38501_ (
    .A1(_02470_),
    .A2(_03296_),
    .ZN(_04187_)
  );
  INV_X1 _38502_ (
    .A(_04187_),
    .ZN(_04188_)
  );
  AND2_X1 _38503_ (
    .A1(_04186_),
    .A2(_04188_),
    .ZN(_04189_)
  );
  INV_X1 _38504_ (
    .A(_04189_),
    .ZN(_04190_)
  );
  AND2_X1 _38505_ (
    .A1(_04158_),
    .A2(_04190_),
    .ZN(_04191_)
  );
  INV_X1 _38506_ (
    .A(_04191_),
    .ZN(_00208_)
  );
  AND2_X1 _38507_ (
    .A1(_04165_),
    .A2(_04173_),
    .ZN(_04192_)
  );
  INV_X1 _38508_ (
    .A(_04192_),
    .ZN(_04193_)
  );
  AND2_X1 _38509_ (
    .A1(decoded_imm_j[30]),
    .A2(_03311_),
    .ZN(_04194_)
  );
  INV_X1 _38510_ (
    .A(_04194_),
    .ZN(_04195_)
  );
  AND2_X1 _38511_ (
    .A1(_22014_),
    .A2(_03312_),
    .ZN(_04196_)
  );
  INV_X1 _38512_ (
    .A(_04196_),
    .ZN(_04197_)
  );
  AND2_X1 _38513_ (
    .A1(_04195_),
    .A2(_04197_),
    .ZN(_04198_)
  );
  INV_X1 _38514_ (
    .A(_04198_),
    .ZN(_04199_)
  );
  AND2_X1 _38515_ (
    .A1(_04193_),
    .A2(_04198_),
    .ZN(_04200_)
  );
  INV_X1 _38516_ (
    .A(_04200_),
    .ZN(_04201_)
  );
  AND2_X1 _38517_ (
    .A1(_04192_),
    .A2(_04199_),
    .ZN(_04202_)
  );
  INV_X1 _38518_ (
    .A(_04202_),
    .ZN(_04203_)
  );
  AND2_X1 _38519_ (
    .A1(instr_jal),
    .A2(_04203_),
    .ZN(_04204_)
  );
  AND2_X1 _38520_ (
    .A1(_04201_),
    .A2(_04204_),
    .ZN(_04205_)
  );
  INV_X1 _38521_ (
    .A(_04205_),
    .ZN(_04206_)
  );
  AND2_X1 _38522_ (
    .A1(_03312_),
    .A2(_04178_),
    .ZN(_04207_)
  );
  INV_X1 _38523_ (
    .A(_04207_),
    .ZN(_04208_)
  );
  AND2_X1 _38524_ (
    .A1(_03311_),
    .A2(_04177_),
    .ZN(_04209_)
  );
  INV_X1 _38525_ (
    .A(_04209_),
    .ZN(_04210_)
  );
  AND2_X1 _38526_ (
    .A1(_21261_),
    .A2(_04210_),
    .ZN(_04211_)
  );
  AND2_X1 _38527_ (
    .A1(_04208_),
    .A2(_04211_),
    .ZN(_04212_)
  );
  INV_X1 _38528_ (
    .A(_04212_),
    .ZN(_04213_)
  );
  AND2_X1 _38529_ (
    .A1(decoder_trigger),
    .A2(_04213_),
    .ZN(_04214_)
  );
  AND2_X1 _38530_ (
    .A1(_04206_),
    .A2(_04214_),
    .ZN(_04215_)
  );
  INV_X1 _38531_ (
    .A(_04215_),
    .ZN(_04216_)
  );
  AND2_X1 _38532_ (
    .A1(_02470_),
    .A2(_03312_),
    .ZN(_04217_)
  );
  INV_X1 _38533_ (
    .A(_04217_),
    .ZN(_04218_)
  );
  AND2_X1 _38534_ (
    .A1(_04216_),
    .A2(_04218_),
    .ZN(_04219_)
  );
  INV_X1 _38535_ (
    .A(_04219_),
    .ZN(_04220_)
  );
  AND2_X1 _38536_ (
    .A1(reg_next_pc[25]),
    .A2(_02928_),
    .ZN(_04221_)
  );
  INV_X1 _38537_ (
    .A(_04221_),
    .ZN(_04222_)
  );
  AND2_X1 _38538_ (
    .A1(_04220_),
    .A2(_04222_),
    .ZN(_04223_)
  );
  INV_X1 _38539_ (
    .A(_04223_),
    .ZN(_00209_)
  );
  AND2_X1 _38540_ (
    .A1(reg_next_pc[26]),
    .A2(_02928_),
    .ZN(_04224_)
  );
  INV_X1 _38541_ (
    .A(_04224_),
    .ZN(_04225_)
  );
  AND2_X1 _38542_ (
    .A1(_04165_),
    .A2(_04195_),
    .ZN(_04226_)
  );
  INV_X1 _38543_ (
    .A(_04226_),
    .ZN(_04227_)
  );
  AND2_X1 _38544_ (
    .A1(_04172_),
    .A2(_04198_),
    .ZN(_04228_)
  );
  INV_X1 _38545_ (
    .A(_04228_),
    .ZN(_04229_)
  );
  AND2_X1 _38546_ (
    .A1(_04226_),
    .A2(_04229_),
    .ZN(_04230_)
  );
  INV_X1 _38547_ (
    .A(_04230_),
    .ZN(_04231_)
  );
  AND2_X1 _38548_ (
    .A1(decoded_imm_j[30]),
    .A2(_03327_),
    .ZN(_04232_)
  );
  INV_X1 _38549_ (
    .A(_04232_),
    .ZN(_04233_)
  );
  AND2_X1 _38550_ (
    .A1(_22014_),
    .A2(_03328_),
    .ZN(_04234_)
  );
  INV_X1 _38551_ (
    .A(_04234_),
    .ZN(_04235_)
  );
  AND2_X1 _38552_ (
    .A1(_04233_),
    .A2(_04235_),
    .ZN(_04236_)
  );
  INV_X1 _38553_ (
    .A(_04236_),
    .ZN(_04237_)
  );
  AND2_X1 _38554_ (
    .A1(_04230_),
    .A2(_04237_),
    .ZN(_04238_)
  );
  INV_X1 _38555_ (
    .A(_04238_),
    .ZN(_04239_)
  );
  AND2_X1 _38556_ (
    .A1(_04231_),
    .A2(_04236_),
    .ZN(_04240_)
  );
  INV_X1 _38557_ (
    .A(_04240_),
    .ZN(_04241_)
  );
  AND2_X1 _38558_ (
    .A1(instr_jal),
    .A2(_04239_),
    .ZN(_04242_)
  );
  AND2_X1 _38559_ (
    .A1(_04241_),
    .A2(_04242_),
    .ZN(_04243_)
  );
  INV_X1 _38560_ (
    .A(_04243_),
    .ZN(_04244_)
  );
  AND2_X1 _38561_ (
    .A1(_03328_),
    .A2(_04210_),
    .ZN(_04245_)
  );
  INV_X1 _38562_ (
    .A(_04245_),
    .ZN(_04246_)
  );
  AND2_X1 _38563_ (
    .A1(_03326_),
    .A2(_04209_),
    .ZN(_04247_)
  );
  INV_X1 _38564_ (
    .A(_04247_),
    .ZN(_04248_)
  );
  AND2_X1 _38565_ (
    .A1(_21261_),
    .A2(_04248_),
    .ZN(_04249_)
  );
  AND2_X1 _38566_ (
    .A1(_04246_),
    .A2(_04249_),
    .ZN(_04250_)
  );
  INV_X1 _38567_ (
    .A(_04250_),
    .ZN(_04251_)
  );
  AND2_X1 _38568_ (
    .A1(decoder_trigger),
    .A2(_04251_),
    .ZN(_04252_)
  );
  AND2_X1 _38569_ (
    .A1(_04244_),
    .A2(_04252_),
    .ZN(_04253_)
  );
  INV_X1 _38570_ (
    .A(_04253_),
    .ZN(_04254_)
  );
  AND2_X1 _38571_ (
    .A1(_02470_),
    .A2(_03328_),
    .ZN(_04255_)
  );
  INV_X1 _38572_ (
    .A(_04255_),
    .ZN(_04256_)
  );
  AND2_X1 _38573_ (
    .A1(_04254_),
    .A2(_04256_),
    .ZN(_04257_)
  );
  INV_X1 _38574_ (
    .A(_04257_),
    .ZN(_04258_)
  );
  AND2_X1 _38575_ (
    .A1(_04225_),
    .A2(_04258_),
    .ZN(_04259_)
  );
  INV_X1 _38576_ (
    .A(_04259_),
    .ZN(_00210_)
  );
  AND2_X1 _38577_ (
    .A1(reg_next_pc[27]),
    .A2(_02928_),
    .ZN(_04260_)
  );
  INV_X1 _38578_ (
    .A(_04260_),
    .ZN(_04261_)
  );
  AND2_X1 _38579_ (
    .A1(_04233_),
    .A2(_04241_),
    .ZN(_04262_)
  );
  INV_X1 _38580_ (
    .A(_04262_),
    .ZN(_04263_)
  );
  AND2_X1 _38581_ (
    .A1(decoded_imm_j[30]),
    .A2(_03343_),
    .ZN(_04264_)
  );
  INV_X1 _38582_ (
    .A(_04264_),
    .ZN(_04265_)
  );
  AND2_X1 _38583_ (
    .A1(_22014_),
    .A2(_03344_),
    .ZN(_04266_)
  );
  INV_X1 _38584_ (
    .A(_04266_),
    .ZN(_04267_)
  );
  AND2_X1 _38585_ (
    .A1(_04265_),
    .A2(_04267_),
    .ZN(_04268_)
  );
  INV_X1 _38586_ (
    .A(_04268_),
    .ZN(_04269_)
  );
  AND2_X1 _38587_ (
    .A1(_04263_),
    .A2(_04268_),
    .ZN(_04270_)
  );
  INV_X1 _38588_ (
    .A(_04270_),
    .ZN(_04271_)
  );
  AND2_X1 _38589_ (
    .A1(_04262_),
    .A2(_04269_),
    .ZN(_04272_)
  );
  INV_X1 _38590_ (
    .A(_04272_),
    .ZN(_04273_)
  );
  AND2_X1 _38591_ (
    .A1(instr_jal),
    .A2(_04273_),
    .ZN(_04274_)
  );
  AND2_X1 _38592_ (
    .A1(_04271_),
    .A2(_04274_),
    .ZN(_04275_)
  );
  INV_X1 _38593_ (
    .A(_04275_),
    .ZN(_04276_)
  );
  AND2_X1 _38594_ (
    .A1(_03344_),
    .A2(_04248_),
    .ZN(_04277_)
  );
  INV_X1 _38595_ (
    .A(_04277_),
    .ZN(_04278_)
  );
  AND2_X1 _38596_ (
    .A1(_03343_),
    .A2(_04247_),
    .ZN(_04279_)
  );
  INV_X1 _38597_ (
    .A(_04279_),
    .ZN(_04280_)
  );
  AND2_X1 _38598_ (
    .A1(_21261_),
    .A2(_04280_),
    .ZN(_04281_)
  );
  AND2_X1 _38599_ (
    .A1(_04278_),
    .A2(_04281_),
    .ZN(_04282_)
  );
  INV_X1 _38600_ (
    .A(_04282_),
    .ZN(_04283_)
  );
  AND2_X1 _38601_ (
    .A1(decoder_trigger),
    .A2(_04283_),
    .ZN(_04284_)
  );
  AND2_X1 _38602_ (
    .A1(_04276_),
    .A2(_04284_),
    .ZN(_04285_)
  );
  INV_X1 _38603_ (
    .A(_04285_),
    .ZN(_04286_)
  );
  AND2_X1 _38604_ (
    .A1(_02470_),
    .A2(_03344_),
    .ZN(_04287_)
  );
  INV_X1 _38605_ (
    .A(_04287_),
    .ZN(_04288_)
  );
  AND2_X1 _38606_ (
    .A1(_04286_),
    .A2(_04288_),
    .ZN(_04289_)
  );
  INV_X1 _38607_ (
    .A(_04289_),
    .ZN(_04290_)
  );
  AND2_X1 _38608_ (
    .A1(_04261_),
    .A2(_04290_),
    .ZN(_04291_)
  );
  INV_X1 _38609_ (
    .A(_04291_),
    .ZN(_00211_)
  );
  AND2_X1 _38610_ (
    .A1(reg_next_pc[28]),
    .A2(_02928_),
    .ZN(_04292_)
  );
  INV_X1 _38611_ (
    .A(_04292_),
    .ZN(_04293_)
  );
  AND2_X1 _38612_ (
    .A1(_04236_),
    .A2(_04268_),
    .ZN(_04294_)
  );
  AND2_X1 _38613_ (
    .A1(_04228_),
    .A2(_04294_),
    .ZN(_04295_)
  );
  INV_X1 _38614_ (
    .A(_04295_),
    .ZN(_04296_)
  );
  AND2_X1 _38615_ (
    .A1(_04227_),
    .A2(_04294_),
    .ZN(_04297_)
  );
  INV_X1 _38616_ (
    .A(_04297_),
    .ZN(_04298_)
  );
  AND2_X1 _38617_ (
    .A1(_04233_),
    .A2(_04265_),
    .ZN(_04299_)
  );
  AND2_X1 _38618_ (
    .A1(_04298_),
    .A2(_04299_),
    .ZN(_04300_)
  );
  AND2_X1 _38619_ (
    .A1(_04296_),
    .A2(_04300_),
    .ZN(_04301_)
  );
  INV_X1 _38620_ (
    .A(_04301_),
    .ZN(_04302_)
  );
  AND2_X1 _38621_ (
    .A1(decoded_imm_j[30]),
    .A2(_03359_),
    .ZN(_04303_)
  );
  INV_X1 _38622_ (
    .A(_04303_),
    .ZN(_04304_)
  );
  AND2_X1 _38623_ (
    .A1(_22014_),
    .A2(_03360_),
    .ZN(_04305_)
  );
  INV_X1 _38624_ (
    .A(_04305_),
    .ZN(_04306_)
  );
  AND2_X1 _38625_ (
    .A1(_04304_),
    .A2(_04306_),
    .ZN(_04307_)
  );
  INV_X1 _38626_ (
    .A(_04307_),
    .ZN(_04308_)
  );
  AND2_X1 _38627_ (
    .A1(_04301_),
    .A2(_04308_),
    .ZN(_04309_)
  );
  INV_X1 _38628_ (
    .A(_04309_),
    .ZN(_04310_)
  );
  AND2_X1 _38629_ (
    .A1(_04302_),
    .A2(_04307_),
    .ZN(_04311_)
  );
  INV_X1 _38630_ (
    .A(_04311_),
    .ZN(_04312_)
  );
  AND2_X1 _38631_ (
    .A1(_04310_),
    .A2(_04312_),
    .ZN(_04313_)
  );
  AND2_X1 _38632_ (
    .A1(instr_jal),
    .A2(_04313_),
    .ZN(_04314_)
  );
  INV_X1 _38633_ (
    .A(_04314_),
    .ZN(_04315_)
  );
  AND2_X1 _38634_ (
    .A1(_03358_),
    .A2(_04279_),
    .ZN(_04316_)
  );
  INV_X1 _38635_ (
    .A(_04316_),
    .ZN(_04317_)
  );
  AND2_X1 _38636_ (
    .A1(_03360_),
    .A2(_04280_),
    .ZN(_04318_)
  );
  INV_X1 _38637_ (
    .A(_04318_),
    .ZN(_04319_)
  );
  AND2_X1 _38638_ (
    .A1(_04317_),
    .A2(_04319_),
    .ZN(_04320_)
  );
  AND2_X1 _38639_ (
    .A1(_21261_),
    .A2(_04320_),
    .ZN(_04321_)
  );
  INV_X1 _38640_ (
    .A(_04321_),
    .ZN(_04322_)
  );
  AND2_X1 _38641_ (
    .A1(decoder_trigger),
    .A2(_04322_),
    .ZN(_04323_)
  );
  AND2_X1 _38642_ (
    .A1(_04315_),
    .A2(_04323_),
    .ZN(_04324_)
  );
  INV_X1 _38643_ (
    .A(_04324_),
    .ZN(_04325_)
  );
  AND2_X1 _38644_ (
    .A1(_02470_),
    .A2(_03360_),
    .ZN(_04326_)
  );
  INV_X1 _38645_ (
    .A(_04326_),
    .ZN(_04327_)
  );
  AND2_X1 _38646_ (
    .A1(_04325_),
    .A2(_04327_),
    .ZN(_04328_)
  );
  INV_X1 _38647_ (
    .A(_04328_),
    .ZN(_04329_)
  );
  AND2_X1 _38648_ (
    .A1(_04293_),
    .A2(_04329_),
    .ZN(_04330_)
  );
  INV_X1 _38649_ (
    .A(_04330_),
    .ZN(_00212_)
  );
  AND2_X1 _38650_ (
    .A1(_04304_),
    .A2(_04312_),
    .ZN(_04331_)
  );
  INV_X1 _38651_ (
    .A(_04331_),
    .ZN(_04332_)
  );
  AND2_X1 _38652_ (
    .A1(decoded_imm_j[30]),
    .A2(_03375_),
    .ZN(_04333_)
  );
  INV_X1 _38653_ (
    .A(_04333_),
    .ZN(_04334_)
  );
  AND2_X1 _38654_ (
    .A1(_22014_),
    .A2(_03376_),
    .ZN(_04335_)
  );
  INV_X1 _38655_ (
    .A(_04335_),
    .ZN(_04336_)
  );
  AND2_X1 _38656_ (
    .A1(_04334_),
    .A2(_04336_),
    .ZN(_04337_)
  );
  INV_X1 _38657_ (
    .A(_04337_),
    .ZN(_04338_)
  );
  AND2_X1 _38658_ (
    .A1(_04332_),
    .A2(_04337_),
    .ZN(_04339_)
  );
  INV_X1 _38659_ (
    .A(_04339_),
    .ZN(_04340_)
  );
  AND2_X1 _38660_ (
    .A1(_04331_),
    .A2(_04338_),
    .ZN(_04341_)
  );
  INV_X1 _38661_ (
    .A(_04341_),
    .ZN(_04342_)
  );
  AND2_X1 _38662_ (
    .A1(instr_jal),
    .A2(_04342_),
    .ZN(_04343_)
  );
  AND2_X1 _38663_ (
    .A1(_04340_),
    .A2(_04343_),
    .ZN(_04344_)
  );
  INV_X1 _38664_ (
    .A(_04344_),
    .ZN(_04345_)
  );
  AND2_X1 _38665_ (
    .A1(_03375_),
    .A2(_04316_),
    .ZN(_04346_)
  );
  INV_X1 _38666_ (
    .A(_04346_),
    .ZN(_04347_)
  );
  AND2_X1 _38667_ (
    .A1(_03376_),
    .A2(_04317_),
    .ZN(_04348_)
  );
  INV_X1 _38668_ (
    .A(_04348_),
    .ZN(_04349_)
  );
  AND2_X1 _38669_ (
    .A1(_04347_),
    .A2(_04349_),
    .ZN(_04350_)
  );
  AND2_X1 _38670_ (
    .A1(_21261_),
    .A2(_04350_),
    .ZN(_04351_)
  );
  INV_X1 _38671_ (
    .A(_04351_),
    .ZN(_04352_)
  );
  AND2_X1 _38672_ (
    .A1(decoder_trigger),
    .A2(_04352_),
    .ZN(_04353_)
  );
  AND2_X1 _38673_ (
    .A1(_04345_),
    .A2(_04353_),
    .ZN(_04354_)
  );
  INV_X1 _38674_ (
    .A(_04354_),
    .ZN(_04355_)
  );
  AND2_X1 _38675_ (
    .A1(_02470_),
    .A2(_03376_),
    .ZN(_04356_)
  );
  INV_X1 _38676_ (
    .A(_04356_),
    .ZN(_04357_)
  );
  AND2_X1 _38677_ (
    .A1(_04355_),
    .A2(_04357_),
    .ZN(_04358_)
  );
  INV_X1 _38678_ (
    .A(_04358_),
    .ZN(_04359_)
  );
  AND2_X1 _38679_ (
    .A1(reg_next_pc[29]),
    .A2(_02928_),
    .ZN(_04360_)
  );
  INV_X1 _38680_ (
    .A(_04360_),
    .ZN(_04361_)
  );
  AND2_X1 _38681_ (
    .A1(_04359_),
    .A2(_04361_),
    .ZN(_04362_)
  );
  INV_X1 _38682_ (
    .A(_04362_),
    .ZN(_00213_)
  );
  AND2_X1 _38683_ (
    .A1(reg_next_pc[30]),
    .A2(_02928_),
    .ZN(_04363_)
  );
  INV_X1 _38684_ (
    .A(_04363_),
    .ZN(_04364_)
  );
  AND2_X1 _38685_ (
    .A1(_04311_),
    .A2(_04337_),
    .ZN(_04365_)
  );
  INV_X1 _38686_ (
    .A(_04365_),
    .ZN(_04366_)
  );
  AND2_X1 _38687_ (
    .A1(_04304_),
    .A2(_04334_),
    .ZN(_04367_)
  );
  AND2_X1 _38688_ (
    .A1(_04366_),
    .A2(_04367_),
    .ZN(_04368_)
  );
  INV_X1 _38689_ (
    .A(_04368_),
    .ZN(_04369_)
  );
  AND2_X1 _38690_ (
    .A1(decoded_imm_j[30]),
    .A2(_03391_),
    .ZN(_04370_)
  );
  INV_X1 _38691_ (
    .A(_04370_),
    .ZN(_04371_)
  );
  AND2_X1 _38692_ (
    .A1(_22014_),
    .A2(_03392_),
    .ZN(_04372_)
  );
  INV_X1 _38693_ (
    .A(_04372_),
    .ZN(_04373_)
  );
  AND2_X1 _38694_ (
    .A1(_04371_),
    .A2(_04373_),
    .ZN(_04374_)
  );
  INV_X1 _38695_ (
    .A(_04374_),
    .ZN(_04375_)
  );
  AND2_X1 _38696_ (
    .A1(_04368_),
    .A2(_04375_),
    .ZN(_04376_)
  );
  INV_X1 _38697_ (
    .A(_04376_),
    .ZN(_04377_)
  );
  AND2_X1 _38698_ (
    .A1(_04369_),
    .A2(_04374_),
    .ZN(_04378_)
  );
  INV_X1 _38699_ (
    .A(_04378_),
    .ZN(_04379_)
  );
  AND2_X1 _38700_ (
    .A1(instr_jal),
    .A2(_04377_),
    .ZN(_04380_)
  );
  AND2_X1 _38701_ (
    .A1(_04379_),
    .A2(_04380_),
    .ZN(_04381_)
  );
  INV_X1 _38702_ (
    .A(_04381_),
    .ZN(_04382_)
  );
  AND2_X1 _38703_ (
    .A1(_03390_),
    .A2(_04346_),
    .ZN(_04383_)
  );
  INV_X1 _38704_ (
    .A(_04383_),
    .ZN(_04384_)
  );
  AND2_X1 _38705_ (
    .A1(_03392_),
    .A2(_04347_),
    .ZN(_04385_)
  );
  INV_X1 _38706_ (
    .A(_04385_),
    .ZN(_04386_)
  );
  AND2_X1 _38707_ (
    .A1(_04384_),
    .A2(_04386_),
    .ZN(_04387_)
  );
  AND2_X1 _38708_ (
    .A1(_21261_),
    .A2(_04387_),
    .ZN(_04388_)
  );
  INV_X1 _38709_ (
    .A(_04388_),
    .ZN(_04389_)
  );
  AND2_X1 _38710_ (
    .A1(decoder_trigger),
    .A2(_04389_),
    .ZN(_04390_)
  );
  AND2_X1 _38711_ (
    .A1(_04382_),
    .A2(_04390_),
    .ZN(_04391_)
  );
  INV_X1 _38712_ (
    .A(_04391_),
    .ZN(_04392_)
  );
  AND2_X1 _38713_ (
    .A1(_02470_),
    .A2(_03392_),
    .ZN(_04393_)
  );
  INV_X1 _38714_ (
    .A(_04393_),
    .ZN(_04394_)
  );
  AND2_X1 _38715_ (
    .A1(_04392_),
    .A2(_04394_),
    .ZN(_04395_)
  );
  INV_X1 _38716_ (
    .A(_04395_),
    .ZN(_04396_)
  );
  AND2_X1 _38717_ (
    .A1(_04364_),
    .A2(_04396_),
    .ZN(_04397_)
  );
  INV_X1 _38718_ (
    .A(_04397_),
    .ZN(_00214_)
  );
  AND2_X1 _38719_ (
    .A1(_04371_),
    .A2(_04379_),
    .ZN(_04398_)
  );
  INV_X1 _38720_ (
    .A(_04398_),
    .ZN(_04399_)
  );
  AND2_X1 _38721_ (
    .A1(_22014_),
    .A2(_03408_),
    .ZN(_04400_)
  );
  INV_X1 _38722_ (
    .A(_04400_),
    .ZN(_04401_)
  );
  AND2_X1 _38723_ (
    .A1(decoded_imm_j[30]),
    .A2(_03407_),
    .ZN(_04402_)
  );
  INV_X1 _38724_ (
    .A(_04402_),
    .ZN(_04403_)
  );
  AND2_X1 _38725_ (
    .A1(decoded_imm_j[30]),
    .A2(_03408_),
    .ZN(_04404_)
  );
  INV_X1 _38726_ (
    .A(_04404_),
    .ZN(_04405_)
  );
  AND2_X1 _38727_ (
    .A1(_22014_),
    .A2(_03407_),
    .ZN(_04406_)
  );
  INV_X1 _38728_ (
    .A(_04406_),
    .ZN(_04407_)
  );
  AND2_X1 _38729_ (
    .A1(_04401_),
    .A2(_04403_),
    .ZN(_04408_)
  );
  AND2_X1 _38730_ (
    .A1(_04405_),
    .A2(_04407_),
    .ZN(_04409_)
  );
  AND2_X1 _38731_ (
    .A1(_04399_),
    .A2(_04408_),
    .ZN(_04410_)
  );
  INV_X1 _38732_ (
    .A(_04410_),
    .ZN(_04411_)
  );
  AND2_X1 _38733_ (
    .A1(_04398_),
    .A2(_04409_),
    .ZN(_04412_)
  );
  INV_X1 _38734_ (
    .A(_04412_),
    .ZN(_04413_)
  );
  AND2_X1 _38735_ (
    .A1(instr_jal),
    .A2(_04413_),
    .ZN(_04414_)
  );
  AND2_X1 _38736_ (
    .A1(_04411_),
    .A2(_04414_),
    .ZN(_04415_)
  );
  INV_X1 _38737_ (
    .A(_04415_),
    .ZN(_04416_)
  );
  AND2_X1 _38738_ (
    .A1(_03407_),
    .A2(_04383_),
    .ZN(_04417_)
  );
  INV_X1 _38739_ (
    .A(_04417_),
    .ZN(_04418_)
  );
  AND2_X1 _38740_ (
    .A1(_03408_),
    .A2(_04384_),
    .ZN(_04419_)
  );
  INV_X1 _38741_ (
    .A(_04419_),
    .ZN(_04420_)
  );
  AND2_X1 _38742_ (
    .A1(_04418_),
    .A2(_04420_),
    .ZN(_04421_)
  );
  AND2_X1 _38743_ (
    .A1(_21261_),
    .A2(_04421_),
    .ZN(_04422_)
  );
  INV_X1 _38744_ (
    .A(_04422_),
    .ZN(_04423_)
  );
  AND2_X1 _38745_ (
    .A1(decoder_trigger),
    .A2(_04423_),
    .ZN(_04424_)
  );
  AND2_X1 _38746_ (
    .A1(_04416_),
    .A2(_04424_),
    .ZN(_04425_)
  );
  INV_X1 _38747_ (
    .A(_04425_),
    .ZN(_04426_)
  );
  AND2_X1 _38748_ (
    .A1(_02470_),
    .A2(_03408_),
    .ZN(_04427_)
  );
  INV_X1 _38749_ (
    .A(_04427_),
    .ZN(_04428_)
  );
  AND2_X1 _38750_ (
    .A1(_04426_),
    .A2(_04428_),
    .ZN(_04429_)
  );
  INV_X1 _38751_ (
    .A(_04429_),
    .ZN(_04430_)
  );
  AND2_X1 _38752_ (
    .A1(reg_next_pc[31]),
    .A2(_02928_),
    .ZN(_04431_)
  );
  INV_X1 _38753_ (
    .A(_04431_),
    .ZN(_04432_)
  );
  AND2_X1 _38754_ (
    .A1(_04430_),
    .A2(_04432_),
    .ZN(_04433_)
  );
  INV_X1 _38755_ (
    .A(_04433_),
    .ZN(_00215_)
  );
  AND2_X1 _38756_ (
    .A1(resetn),
    .A2(_29147_[0]),
    .ZN(_00216_)
  );
  AND2_X1 _38757_ (
    .A1(count_cycle[0]),
    .A2(count_cycle[1]),
    .ZN(_04434_)
  );
  INV_X1 _38758_ (
    .A(_04434_),
    .ZN(_04435_)
  );
  AND2_X1 _38759_ (
    .A1(_22153_),
    .A2(_22154_),
    .ZN(_04436_)
  );
  INV_X1 _38760_ (
    .A(_04436_),
    .ZN(_04437_)
  );
  AND2_X1 _38761_ (
    .A1(resetn),
    .A2(_04437_),
    .ZN(_04438_)
  );
  AND2_X1 _38762_ (
    .A1(_04435_),
    .A2(_04438_),
    .ZN(_00217_)
  );
  AND2_X1 _38763_ (
    .A1(count_cycle[2]),
    .A2(_04434_),
    .ZN(_04439_)
  );
  INV_X1 _38764_ (
    .A(_04439_),
    .ZN(_04440_)
  );
  AND2_X1 _38765_ (
    .A1(_22155_),
    .A2(_04435_),
    .ZN(_04441_)
  );
  INV_X1 _38766_ (
    .A(_04441_),
    .ZN(_04442_)
  );
  AND2_X1 _38767_ (
    .A1(resetn),
    .A2(_04442_),
    .ZN(_04443_)
  );
  AND2_X1 _38768_ (
    .A1(_04440_),
    .A2(_04443_),
    .ZN(_00218_)
  );
  AND2_X1 _38769_ (
    .A1(count_cycle[3]),
    .A2(_04439_),
    .ZN(_04444_)
  );
  INV_X1 _38770_ (
    .A(_04444_),
    .ZN(_04445_)
  );
  AND2_X1 _38771_ (
    .A1(_22156_),
    .A2(_04440_),
    .ZN(_04446_)
  );
  INV_X1 _38772_ (
    .A(_04446_),
    .ZN(_04447_)
  );
  AND2_X1 _38773_ (
    .A1(resetn),
    .A2(_04447_),
    .ZN(_04448_)
  );
  AND2_X1 _38774_ (
    .A1(_04445_),
    .A2(_04448_),
    .ZN(_00219_)
  );
  AND2_X1 _38775_ (
    .A1(count_cycle[4]),
    .A2(_04444_),
    .ZN(_04449_)
  );
  INV_X1 _38776_ (
    .A(_04449_),
    .ZN(_04450_)
  );
  AND2_X1 _38777_ (
    .A1(_22157_),
    .A2(_04445_),
    .ZN(_04451_)
  );
  INV_X1 _38778_ (
    .A(_04451_),
    .ZN(_04452_)
  );
  AND2_X1 _38779_ (
    .A1(resetn),
    .A2(_04452_),
    .ZN(_04453_)
  );
  AND2_X1 _38780_ (
    .A1(_04450_),
    .A2(_04453_),
    .ZN(_00220_)
  );
  AND2_X1 _38781_ (
    .A1(count_cycle[5]),
    .A2(_04449_),
    .ZN(_04454_)
  );
  INV_X1 _38782_ (
    .A(_04454_),
    .ZN(_04455_)
  );
  AND2_X1 _38783_ (
    .A1(_22158_),
    .A2(_04450_),
    .ZN(_04456_)
  );
  INV_X1 _38784_ (
    .A(_04456_),
    .ZN(_04457_)
  );
  AND2_X1 _38785_ (
    .A1(resetn),
    .A2(_04457_),
    .ZN(_04458_)
  );
  AND2_X1 _38786_ (
    .A1(_04455_),
    .A2(_04458_),
    .ZN(_00221_)
  );
  AND2_X1 _38787_ (
    .A1(count_cycle[6]),
    .A2(_04454_),
    .ZN(_04459_)
  );
  INV_X1 _38788_ (
    .A(_04459_),
    .ZN(_04460_)
  );
  AND2_X1 _38789_ (
    .A1(_22159_),
    .A2(_04455_),
    .ZN(_04461_)
  );
  INV_X1 _38790_ (
    .A(_04461_),
    .ZN(_04462_)
  );
  AND2_X1 _38791_ (
    .A1(resetn),
    .A2(_04462_),
    .ZN(_04463_)
  );
  AND2_X1 _38792_ (
    .A1(_04460_),
    .A2(_04463_),
    .ZN(_00222_)
  );
  AND2_X1 _38793_ (
    .A1(count_cycle[7]),
    .A2(_04459_),
    .ZN(_04464_)
  );
  INV_X1 _38794_ (
    .A(_04464_),
    .ZN(_04465_)
  );
  AND2_X1 _38795_ (
    .A1(_22160_),
    .A2(_04460_),
    .ZN(_04466_)
  );
  INV_X1 _38796_ (
    .A(_04466_),
    .ZN(_04467_)
  );
  AND2_X1 _38797_ (
    .A1(resetn),
    .A2(_04467_),
    .ZN(_04468_)
  );
  AND2_X1 _38798_ (
    .A1(_04465_),
    .A2(_04468_),
    .ZN(_00223_)
  );
  AND2_X1 _38799_ (
    .A1(count_cycle[8]),
    .A2(_04464_),
    .ZN(_04469_)
  );
  INV_X1 _38800_ (
    .A(_04469_),
    .ZN(_04470_)
  );
  AND2_X1 _38801_ (
    .A1(_22161_),
    .A2(_04465_),
    .ZN(_04471_)
  );
  INV_X1 _38802_ (
    .A(_04471_),
    .ZN(_04472_)
  );
  AND2_X1 _38803_ (
    .A1(resetn),
    .A2(_04472_),
    .ZN(_04473_)
  );
  AND2_X1 _38804_ (
    .A1(_04470_),
    .A2(_04473_),
    .ZN(_00224_)
  );
  AND2_X1 _38805_ (
    .A1(count_cycle[9]),
    .A2(_04469_),
    .ZN(_04474_)
  );
  INV_X1 _38806_ (
    .A(_04474_),
    .ZN(_04475_)
  );
  AND2_X1 _38807_ (
    .A1(_22162_),
    .A2(_04470_),
    .ZN(_04476_)
  );
  INV_X1 _38808_ (
    .A(_04476_),
    .ZN(_04477_)
  );
  AND2_X1 _38809_ (
    .A1(resetn),
    .A2(_04477_),
    .ZN(_04478_)
  );
  AND2_X1 _38810_ (
    .A1(_04475_),
    .A2(_04478_),
    .ZN(_00225_)
  );
  AND2_X1 _38811_ (
    .A1(count_cycle[10]),
    .A2(_04474_),
    .ZN(_04479_)
  );
  INV_X1 _38812_ (
    .A(_04479_),
    .ZN(_04480_)
  );
  AND2_X1 _38813_ (
    .A1(_22163_),
    .A2(_04475_),
    .ZN(_04481_)
  );
  INV_X1 _38814_ (
    .A(_04481_),
    .ZN(_04482_)
  );
  AND2_X1 _38815_ (
    .A1(resetn),
    .A2(_04482_),
    .ZN(_04483_)
  );
  AND2_X1 _38816_ (
    .A1(_04480_),
    .A2(_04483_),
    .ZN(_00226_)
  );
  AND2_X1 _38817_ (
    .A1(count_cycle[11]),
    .A2(_04479_),
    .ZN(_04484_)
  );
  INV_X1 _38818_ (
    .A(_04484_),
    .ZN(_04485_)
  );
  AND2_X1 _38819_ (
    .A1(_22164_),
    .A2(_04480_),
    .ZN(_04486_)
  );
  INV_X1 _38820_ (
    .A(_04486_),
    .ZN(_04487_)
  );
  AND2_X1 _38821_ (
    .A1(resetn),
    .A2(_04487_),
    .ZN(_04488_)
  );
  AND2_X1 _38822_ (
    .A1(_04485_),
    .A2(_04488_),
    .ZN(_00227_)
  );
  AND2_X1 _38823_ (
    .A1(count_cycle[12]),
    .A2(_04484_),
    .ZN(_04489_)
  );
  INV_X1 _38824_ (
    .A(_04489_),
    .ZN(_04490_)
  );
  AND2_X1 _38825_ (
    .A1(_22165_),
    .A2(_04485_),
    .ZN(_04491_)
  );
  INV_X1 _38826_ (
    .A(_04491_),
    .ZN(_04492_)
  );
  AND2_X1 _38827_ (
    .A1(resetn),
    .A2(_04492_),
    .ZN(_04493_)
  );
  AND2_X1 _38828_ (
    .A1(_04490_),
    .A2(_04493_),
    .ZN(_00228_)
  );
  AND2_X1 _38829_ (
    .A1(count_cycle[13]),
    .A2(_04489_),
    .ZN(_04494_)
  );
  INV_X1 _38830_ (
    .A(_04494_),
    .ZN(_04495_)
  );
  AND2_X1 _38831_ (
    .A1(_22166_),
    .A2(_04490_),
    .ZN(_04496_)
  );
  INV_X1 _38832_ (
    .A(_04496_),
    .ZN(_04497_)
  );
  AND2_X1 _38833_ (
    .A1(resetn),
    .A2(_04497_),
    .ZN(_04498_)
  );
  AND2_X1 _38834_ (
    .A1(_04495_),
    .A2(_04498_),
    .ZN(_00229_)
  );
  AND2_X1 _38835_ (
    .A1(count_cycle[14]),
    .A2(_04494_),
    .ZN(_04499_)
  );
  INV_X1 _38836_ (
    .A(_04499_),
    .ZN(_04500_)
  );
  AND2_X1 _38837_ (
    .A1(_22167_),
    .A2(_04495_),
    .ZN(_04501_)
  );
  INV_X1 _38838_ (
    .A(_04501_),
    .ZN(_04502_)
  );
  AND2_X1 _38839_ (
    .A1(resetn),
    .A2(_04502_),
    .ZN(_04503_)
  );
  AND2_X1 _38840_ (
    .A1(_04500_),
    .A2(_04503_),
    .ZN(_00230_)
  );
  AND2_X1 _38841_ (
    .A1(count_cycle[15]),
    .A2(_04499_),
    .ZN(_04504_)
  );
  INV_X1 _38842_ (
    .A(_04504_),
    .ZN(_04505_)
  );
  AND2_X1 _38843_ (
    .A1(_22168_),
    .A2(_04500_),
    .ZN(_04506_)
  );
  INV_X1 _38844_ (
    .A(_04506_),
    .ZN(_04507_)
  );
  AND2_X1 _38845_ (
    .A1(resetn),
    .A2(_04507_),
    .ZN(_04508_)
  );
  AND2_X1 _38846_ (
    .A1(_04505_),
    .A2(_04508_),
    .ZN(_00231_)
  );
  AND2_X1 _38847_ (
    .A1(count_cycle[16]),
    .A2(_04504_),
    .ZN(_04509_)
  );
  INV_X1 _38848_ (
    .A(_04509_),
    .ZN(_04510_)
  );
  AND2_X1 _38849_ (
    .A1(_22169_),
    .A2(_04505_),
    .ZN(_04511_)
  );
  INV_X1 _38850_ (
    .A(_04511_),
    .ZN(_04512_)
  );
  AND2_X1 _38851_ (
    .A1(resetn),
    .A2(_04512_),
    .ZN(_04513_)
  );
  AND2_X1 _38852_ (
    .A1(_04510_),
    .A2(_04513_),
    .ZN(_00232_)
  );
  AND2_X1 _38853_ (
    .A1(count_cycle[17]),
    .A2(_04509_),
    .ZN(_04514_)
  );
  INV_X1 _38854_ (
    .A(_04514_),
    .ZN(_04515_)
  );
  AND2_X1 _38855_ (
    .A1(_22170_),
    .A2(_04510_),
    .ZN(_04516_)
  );
  INV_X1 _38856_ (
    .A(_04516_),
    .ZN(_04517_)
  );
  AND2_X1 _38857_ (
    .A1(resetn),
    .A2(_04517_),
    .ZN(_04518_)
  );
  AND2_X1 _38858_ (
    .A1(_04515_),
    .A2(_04518_),
    .ZN(_00233_)
  );
  AND2_X1 _38859_ (
    .A1(count_cycle[18]),
    .A2(_04514_),
    .ZN(_04519_)
  );
  INV_X1 _38860_ (
    .A(_04519_),
    .ZN(_04520_)
  );
  AND2_X1 _38861_ (
    .A1(_22171_),
    .A2(_04515_),
    .ZN(_04521_)
  );
  INV_X1 _38862_ (
    .A(_04521_),
    .ZN(_04522_)
  );
  AND2_X1 _38863_ (
    .A1(resetn),
    .A2(_04522_),
    .ZN(_04523_)
  );
  AND2_X1 _38864_ (
    .A1(_04520_),
    .A2(_04523_),
    .ZN(_00234_)
  );
  AND2_X1 _38865_ (
    .A1(count_cycle[19]),
    .A2(_04519_),
    .ZN(_04524_)
  );
  INV_X1 _38866_ (
    .A(_04524_),
    .ZN(_04525_)
  );
  AND2_X1 _38867_ (
    .A1(_22172_),
    .A2(_04520_),
    .ZN(_04526_)
  );
  INV_X1 _38868_ (
    .A(_04526_),
    .ZN(_04527_)
  );
  AND2_X1 _38869_ (
    .A1(resetn),
    .A2(_04527_),
    .ZN(_04528_)
  );
  AND2_X1 _38870_ (
    .A1(_04525_),
    .A2(_04528_),
    .ZN(_00235_)
  );
  AND2_X1 _38871_ (
    .A1(count_cycle[20]),
    .A2(_04524_),
    .ZN(_04529_)
  );
  INV_X1 _38872_ (
    .A(_04529_),
    .ZN(_04530_)
  );
  AND2_X1 _38873_ (
    .A1(_22173_),
    .A2(_04525_),
    .ZN(_04531_)
  );
  INV_X1 _38874_ (
    .A(_04531_),
    .ZN(_04532_)
  );
  AND2_X1 _38875_ (
    .A1(resetn),
    .A2(_04532_),
    .ZN(_04533_)
  );
  AND2_X1 _38876_ (
    .A1(_04530_),
    .A2(_04533_),
    .ZN(_00236_)
  );
  AND2_X1 _38877_ (
    .A1(count_cycle[21]),
    .A2(_04529_),
    .ZN(_04534_)
  );
  INV_X1 _38878_ (
    .A(_04534_),
    .ZN(_04535_)
  );
  AND2_X1 _38879_ (
    .A1(_22174_),
    .A2(_04530_),
    .ZN(_04536_)
  );
  INV_X1 _38880_ (
    .A(_04536_),
    .ZN(_04537_)
  );
  AND2_X1 _38881_ (
    .A1(resetn),
    .A2(_04537_),
    .ZN(_04538_)
  );
  AND2_X1 _38882_ (
    .A1(_04535_),
    .A2(_04538_),
    .ZN(_00237_)
  );
  AND2_X1 _38883_ (
    .A1(count_cycle[22]),
    .A2(_04534_),
    .ZN(_04539_)
  );
  INV_X1 _38884_ (
    .A(_04539_),
    .ZN(_04540_)
  );
  AND2_X1 _38885_ (
    .A1(_22175_),
    .A2(_04535_),
    .ZN(_04541_)
  );
  INV_X1 _38886_ (
    .A(_04541_),
    .ZN(_04542_)
  );
  AND2_X1 _38887_ (
    .A1(resetn),
    .A2(_04542_),
    .ZN(_04543_)
  );
  AND2_X1 _38888_ (
    .A1(_04540_),
    .A2(_04543_),
    .ZN(_00238_)
  );
  AND2_X1 _38889_ (
    .A1(count_cycle[23]),
    .A2(_04539_),
    .ZN(_04544_)
  );
  INV_X1 _38890_ (
    .A(_04544_),
    .ZN(_04545_)
  );
  AND2_X1 _38891_ (
    .A1(_22176_),
    .A2(_04540_),
    .ZN(_04546_)
  );
  INV_X1 _38892_ (
    .A(_04546_),
    .ZN(_04547_)
  );
  AND2_X1 _38893_ (
    .A1(resetn),
    .A2(_04547_),
    .ZN(_04548_)
  );
  AND2_X1 _38894_ (
    .A1(_04545_),
    .A2(_04548_),
    .ZN(_00239_)
  );
  AND2_X1 _38895_ (
    .A1(count_cycle[24]),
    .A2(_04544_),
    .ZN(_04549_)
  );
  INV_X1 _38896_ (
    .A(_04549_),
    .ZN(_04550_)
  );
  AND2_X1 _38897_ (
    .A1(_22177_),
    .A2(_04545_),
    .ZN(_04551_)
  );
  INV_X1 _38898_ (
    .A(_04551_),
    .ZN(_04552_)
  );
  AND2_X1 _38899_ (
    .A1(resetn),
    .A2(_04552_),
    .ZN(_04553_)
  );
  AND2_X1 _38900_ (
    .A1(_04550_),
    .A2(_04553_),
    .ZN(_00240_)
  );
  AND2_X1 _38901_ (
    .A1(count_cycle[25]),
    .A2(_04549_),
    .ZN(_04554_)
  );
  INV_X1 _38902_ (
    .A(_04554_),
    .ZN(_04555_)
  );
  AND2_X1 _38903_ (
    .A1(_22178_),
    .A2(_04550_),
    .ZN(_04556_)
  );
  INV_X1 _38904_ (
    .A(_04556_),
    .ZN(_04557_)
  );
  AND2_X1 _38905_ (
    .A1(resetn),
    .A2(_04557_),
    .ZN(_04558_)
  );
  AND2_X1 _38906_ (
    .A1(_04555_),
    .A2(_04558_),
    .ZN(_00241_)
  );
  AND2_X1 _38907_ (
    .A1(count_cycle[26]),
    .A2(_04554_),
    .ZN(_04559_)
  );
  INV_X1 _38908_ (
    .A(_04559_),
    .ZN(_04560_)
  );
  AND2_X1 _38909_ (
    .A1(_22179_),
    .A2(_04555_),
    .ZN(_04561_)
  );
  INV_X1 _38910_ (
    .A(_04561_),
    .ZN(_04562_)
  );
  AND2_X1 _38911_ (
    .A1(resetn),
    .A2(_04562_),
    .ZN(_04563_)
  );
  AND2_X1 _38912_ (
    .A1(_04560_),
    .A2(_04563_),
    .ZN(_00242_)
  );
  AND2_X1 _38913_ (
    .A1(count_cycle[27]),
    .A2(_04559_),
    .ZN(_04564_)
  );
  INV_X1 _38914_ (
    .A(_04564_),
    .ZN(_04565_)
  );
  AND2_X1 _38915_ (
    .A1(_22180_),
    .A2(_04560_),
    .ZN(_04566_)
  );
  INV_X1 _38916_ (
    .A(_04566_),
    .ZN(_04567_)
  );
  AND2_X1 _38917_ (
    .A1(resetn),
    .A2(_04567_),
    .ZN(_04568_)
  );
  AND2_X1 _38918_ (
    .A1(_04565_),
    .A2(_04568_),
    .ZN(_00243_)
  );
  AND2_X1 _38919_ (
    .A1(count_cycle[28]),
    .A2(_04564_),
    .ZN(_04569_)
  );
  INV_X1 _38920_ (
    .A(_04569_),
    .ZN(_04570_)
  );
  AND2_X1 _38921_ (
    .A1(_22181_),
    .A2(_04565_),
    .ZN(_04571_)
  );
  INV_X1 _38922_ (
    .A(_04571_),
    .ZN(_04572_)
  );
  AND2_X1 _38923_ (
    .A1(resetn),
    .A2(_04572_),
    .ZN(_04573_)
  );
  AND2_X1 _38924_ (
    .A1(_04570_),
    .A2(_04573_),
    .ZN(_00244_)
  );
  AND2_X1 _38925_ (
    .A1(count_cycle[29]),
    .A2(_04569_),
    .ZN(_04574_)
  );
  INV_X1 _38926_ (
    .A(_04574_),
    .ZN(_04575_)
  );
  AND2_X1 _38927_ (
    .A1(_22182_),
    .A2(_04570_),
    .ZN(_04576_)
  );
  INV_X1 _38928_ (
    .A(_04576_),
    .ZN(_04577_)
  );
  AND2_X1 _38929_ (
    .A1(resetn),
    .A2(_04577_),
    .ZN(_04578_)
  );
  AND2_X1 _38930_ (
    .A1(_04575_),
    .A2(_04578_),
    .ZN(_00245_)
  );
  AND2_X1 _38931_ (
    .A1(count_cycle[30]),
    .A2(_04574_),
    .ZN(_04579_)
  );
  INV_X1 _38932_ (
    .A(_04579_),
    .ZN(_04580_)
  );
  AND2_X1 _38933_ (
    .A1(_22183_),
    .A2(_04575_),
    .ZN(_04581_)
  );
  INV_X1 _38934_ (
    .A(_04581_),
    .ZN(_04582_)
  );
  AND2_X1 _38935_ (
    .A1(resetn),
    .A2(_04582_),
    .ZN(_04583_)
  );
  AND2_X1 _38936_ (
    .A1(_04580_),
    .A2(_04583_),
    .ZN(_00246_)
  );
  AND2_X1 _38937_ (
    .A1(count_cycle[31]),
    .A2(_04579_),
    .ZN(_04584_)
  );
  INV_X1 _38938_ (
    .A(_04584_),
    .ZN(_04585_)
  );
  AND2_X1 _38939_ (
    .A1(_22184_),
    .A2(_04580_),
    .ZN(_04586_)
  );
  INV_X1 _38940_ (
    .A(_04586_),
    .ZN(_04587_)
  );
  AND2_X1 _38941_ (
    .A1(resetn),
    .A2(_04587_),
    .ZN(_04588_)
  );
  AND2_X1 _38942_ (
    .A1(_04585_),
    .A2(_04588_),
    .ZN(_00247_)
  );
  AND2_X1 _38943_ (
    .A1(count_cycle[32]),
    .A2(_04584_),
    .ZN(_04589_)
  );
  INV_X1 _38944_ (
    .A(_04589_),
    .ZN(_04590_)
  );
  AND2_X1 _38945_ (
    .A1(_22185_),
    .A2(_04585_),
    .ZN(_04591_)
  );
  INV_X1 _38946_ (
    .A(_04591_),
    .ZN(_04592_)
  );
  AND2_X1 _38947_ (
    .A1(resetn),
    .A2(_04592_),
    .ZN(_04593_)
  );
  AND2_X1 _38948_ (
    .A1(_04590_),
    .A2(_04593_),
    .ZN(_00248_)
  );
  AND2_X1 _38949_ (
    .A1(count_cycle[33]),
    .A2(_04589_),
    .ZN(_04594_)
  );
  INV_X1 _38950_ (
    .A(_04594_),
    .ZN(_04595_)
  );
  AND2_X1 _38951_ (
    .A1(_22186_),
    .A2(_04590_),
    .ZN(_04596_)
  );
  INV_X1 _38952_ (
    .A(_04596_),
    .ZN(_04597_)
  );
  AND2_X1 _38953_ (
    .A1(resetn),
    .A2(_04597_),
    .ZN(_04598_)
  );
  AND2_X1 _38954_ (
    .A1(_04595_),
    .A2(_04598_),
    .ZN(_00249_)
  );
  AND2_X1 _38955_ (
    .A1(count_cycle[34]),
    .A2(_04594_),
    .ZN(_04599_)
  );
  INV_X1 _38956_ (
    .A(_04599_),
    .ZN(_04600_)
  );
  AND2_X1 _38957_ (
    .A1(_22187_),
    .A2(_04595_),
    .ZN(_04601_)
  );
  INV_X1 _38958_ (
    .A(_04601_),
    .ZN(_04602_)
  );
  AND2_X1 _38959_ (
    .A1(resetn),
    .A2(_04602_),
    .ZN(_04603_)
  );
  AND2_X1 _38960_ (
    .A1(_04600_),
    .A2(_04603_),
    .ZN(_00250_)
  );
  AND2_X1 _38961_ (
    .A1(count_cycle[35]),
    .A2(_04599_),
    .ZN(_04604_)
  );
  INV_X1 _38962_ (
    .A(_04604_),
    .ZN(_04605_)
  );
  AND2_X1 _38963_ (
    .A1(_22188_),
    .A2(_04600_),
    .ZN(_04606_)
  );
  INV_X1 _38964_ (
    .A(_04606_),
    .ZN(_04607_)
  );
  AND2_X1 _38965_ (
    .A1(resetn),
    .A2(_04607_),
    .ZN(_04608_)
  );
  AND2_X1 _38966_ (
    .A1(_04605_),
    .A2(_04608_),
    .ZN(_00251_)
  );
  AND2_X1 _38967_ (
    .A1(count_cycle[36]),
    .A2(_04604_),
    .ZN(_04609_)
  );
  INV_X1 _38968_ (
    .A(_04609_),
    .ZN(_04610_)
  );
  AND2_X1 _38969_ (
    .A1(_22189_),
    .A2(_04605_),
    .ZN(_04611_)
  );
  INV_X1 _38970_ (
    .A(_04611_),
    .ZN(_04612_)
  );
  AND2_X1 _38971_ (
    .A1(resetn),
    .A2(_04612_),
    .ZN(_04613_)
  );
  AND2_X1 _38972_ (
    .A1(_04610_),
    .A2(_04613_),
    .ZN(_00252_)
  );
  AND2_X1 _38973_ (
    .A1(count_cycle[37]),
    .A2(_04609_),
    .ZN(_04614_)
  );
  INV_X1 _38974_ (
    .A(_04614_),
    .ZN(_04615_)
  );
  AND2_X1 _38975_ (
    .A1(_22190_),
    .A2(_04610_),
    .ZN(_04616_)
  );
  INV_X1 _38976_ (
    .A(_04616_),
    .ZN(_04617_)
  );
  AND2_X1 _38977_ (
    .A1(resetn),
    .A2(_04617_),
    .ZN(_04618_)
  );
  AND2_X1 _38978_ (
    .A1(_04615_),
    .A2(_04618_),
    .ZN(_00253_)
  );
  AND2_X1 _38979_ (
    .A1(count_cycle[38]),
    .A2(_04614_),
    .ZN(_04619_)
  );
  INV_X1 _38980_ (
    .A(_04619_),
    .ZN(_04620_)
  );
  AND2_X1 _38981_ (
    .A1(_22191_),
    .A2(_04615_),
    .ZN(_04621_)
  );
  INV_X1 _38982_ (
    .A(_04621_),
    .ZN(_04622_)
  );
  AND2_X1 _38983_ (
    .A1(resetn),
    .A2(_04622_),
    .ZN(_04623_)
  );
  AND2_X1 _38984_ (
    .A1(_04620_),
    .A2(_04623_),
    .ZN(_00254_)
  );
  AND2_X1 _38985_ (
    .A1(count_cycle[39]),
    .A2(_04619_),
    .ZN(_04624_)
  );
  INV_X1 _38986_ (
    .A(_04624_),
    .ZN(_04625_)
  );
  AND2_X1 _38987_ (
    .A1(_22192_),
    .A2(_04620_),
    .ZN(_04626_)
  );
  INV_X1 _38988_ (
    .A(_04626_),
    .ZN(_04627_)
  );
  AND2_X1 _38989_ (
    .A1(resetn),
    .A2(_04627_),
    .ZN(_04628_)
  );
  AND2_X1 _38990_ (
    .A1(_04625_),
    .A2(_04628_),
    .ZN(_00255_)
  );
  AND2_X1 _38991_ (
    .A1(count_cycle[40]),
    .A2(_04624_),
    .ZN(_04629_)
  );
  INV_X1 _38992_ (
    .A(_04629_),
    .ZN(_04630_)
  );
  AND2_X1 _38993_ (
    .A1(_22193_),
    .A2(_04625_),
    .ZN(_04631_)
  );
  INV_X1 _38994_ (
    .A(_04631_),
    .ZN(_04632_)
  );
  AND2_X1 _38995_ (
    .A1(resetn),
    .A2(_04632_),
    .ZN(_04633_)
  );
  AND2_X1 _38996_ (
    .A1(_04630_),
    .A2(_04633_),
    .ZN(_00256_)
  );
  AND2_X1 _38997_ (
    .A1(count_cycle[41]),
    .A2(_04629_),
    .ZN(_04634_)
  );
  INV_X1 _38998_ (
    .A(_04634_),
    .ZN(_04635_)
  );
  AND2_X1 _38999_ (
    .A1(_22194_),
    .A2(_04630_),
    .ZN(_04636_)
  );
  INV_X1 _39000_ (
    .A(_04636_),
    .ZN(_04637_)
  );
  AND2_X1 _39001_ (
    .A1(resetn),
    .A2(_04637_),
    .ZN(_04638_)
  );
  AND2_X1 _39002_ (
    .A1(_04635_),
    .A2(_04638_),
    .ZN(_00257_)
  );
  AND2_X1 _39003_ (
    .A1(count_cycle[42]),
    .A2(_04634_),
    .ZN(_04639_)
  );
  INV_X1 _39004_ (
    .A(_04639_),
    .ZN(_04640_)
  );
  AND2_X1 _39005_ (
    .A1(_22195_),
    .A2(_04635_),
    .ZN(_04641_)
  );
  INV_X1 _39006_ (
    .A(_04641_),
    .ZN(_04642_)
  );
  AND2_X1 _39007_ (
    .A1(resetn),
    .A2(_04642_),
    .ZN(_04643_)
  );
  AND2_X1 _39008_ (
    .A1(_04640_),
    .A2(_04643_),
    .ZN(_00258_)
  );
  AND2_X1 _39009_ (
    .A1(count_cycle[43]),
    .A2(_04639_),
    .ZN(_04644_)
  );
  INV_X1 _39010_ (
    .A(_04644_),
    .ZN(_04645_)
  );
  AND2_X1 _39011_ (
    .A1(_22196_),
    .A2(_04640_),
    .ZN(_04646_)
  );
  INV_X1 _39012_ (
    .A(_04646_),
    .ZN(_04647_)
  );
  AND2_X1 _39013_ (
    .A1(resetn),
    .A2(_04647_),
    .ZN(_04648_)
  );
  AND2_X1 _39014_ (
    .A1(_04645_),
    .A2(_04648_),
    .ZN(_00259_)
  );
  AND2_X1 _39015_ (
    .A1(count_cycle[44]),
    .A2(_04644_),
    .ZN(_04649_)
  );
  INV_X1 _39016_ (
    .A(_04649_),
    .ZN(_04650_)
  );
  AND2_X1 _39017_ (
    .A1(_22197_),
    .A2(_04645_),
    .ZN(_04651_)
  );
  INV_X1 _39018_ (
    .A(_04651_),
    .ZN(_04652_)
  );
  AND2_X1 _39019_ (
    .A1(resetn),
    .A2(_04652_),
    .ZN(_04653_)
  );
  AND2_X1 _39020_ (
    .A1(_04650_),
    .A2(_04653_),
    .ZN(_00260_)
  );
  AND2_X1 _39021_ (
    .A1(count_cycle[45]),
    .A2(_04649_),
    .ZN(_04654_)
  );
  INV_X1 _39022_ (
    .A(_04654_),
    .ZN(_04655_)
  );
  AND2_X1 _39023_ (
    .A1(_22198_),
    .A2(_04650_),
    .ZN(_04656_)
  );
  INV_X1 _39024_ (
    .A(_04656_),
    .ZN(_04657_)
  );
  AND2_X1 _39025_ (
    .A1(resetn),
    .A2(_04657_),
    .ZN(_04658_)
  );
  AND2_X1 _39026_ (
    .A1(_04655_),
    .A2(_04658_),
    .ZN(_00261_)
  );
  AND2_X1 _39027_ (
    .A1(count_cycle[46]),
    .A2(_04654_),
    .ZN(_04659_)
  );
  INV_X1 _39028_ (
    .A(_04659_),
    .ZN(_04660_)
  );
  AND2_X1 _39029_ (
    .A1(_22199_),
    .A2(_04655_),
    .ZN(_04661_)
  );
  INV_X1 _39030_ (
    .A(_04661_),
    .ZN(_04662_)
  );
  AND2_X1 _39031_ (
    .A1(resetn),
    .A2(_04662_),
    .ZN(_04663_)
  );
  AND2_X1 _39032_ (
    .A1(_04660_),
    .A2(_04663_),
    .ZN(_00262_)
  );
  AND2_X1 _39033_ (
    .A1(count_cycle[47]),
    .A2(_04659_),
    .ZN(_04664_)
  );
  INV_X1 _39034_ (
    .A(_04664_),
    .ZN(_04665_)
  );
  AND2_X1 _39035_ (
    .A1(_22200_),
    .A2(_04660_),
    .ZN(_04666_)
  );
  INV_X1 _39036_ (
    .A(_04666_),
    .ZN(_04667_)
  );
  AND2_X1 _39037_ (
    .A1(resetn),
    .A2(_04667_),
    .ZN(_04668_)
  );
  AND2_X1 _39038_ (
    .A1(_04665_),
    .A2(_04668_),
    .ZN(_00263_)
  );
  AND2_X1 _39039_ (
    .A1(count_cycle[48]),
    .A2(_04664_),
    .ZN(_04669_)
  );
  INV_X1 _39040_ (
    .A(_04669_),
    .ZN(_04670_)
  );
  AND2_X1 _39041_ (
    .A1(_22201_),
    .A2(_04665_),
    .ZN(_04671_)
  );
  INV_X1 _39042_ (
    .A(_04671_),
    .ZN(_04672_)
  );
  AND2_X1 _39043_ (
    .A1(resetn),
    .A2(_04672_),
    .ZN(_04673_)
  );
  AND2_X1 _39044_ (
    .A1(_04670_),
    .A2(_04673_),
    .ZN(_00264_)
  );
  AND2_X1 _39045_ (
    .A1(count_cycle[49]),
    .A2(_04669_),
    .ZN(_04674_)
  );
  INV_X1 _39046_ (
    .A(_04674_),
    .ZN(_04675_)
  );
  AND2_X1 _39047_ (
    .A1(_22202_),
    .A2(_04670_),
    .ZN(_04676_)
  );
  INV_X1 _39048_ (
    .A(_04676_),
    .ZN(_04677_)
  );
  AND2_X1 _39049_ (
    .A1(resetn),
    .A2(_04677_),
    .ZN(_04678_)
  );
  AND2_X1 _39050_ (
    .A1(_04675_),
    .A2(_04678_),
    .ZN(_00265_)
  );
  AND2_X1 _39051_ (
    .A1(count_cycle[50]),
    .A2(_04674_),
    .ZN(_04679_)
  );
  INV_X1 _39052_ (
    .A(_04679_),
    .ZN(_04680_)
  );
  AND2_X1 _39053_ (
    .A1(_22203_),
    .A2(_04675_),
    .ZN(_04681_)
  );
  INV_X1 _39054_ (
    .A(_04681_),
    .ZN(_04682_)
  );
  AND2_X1 _39055_ (
    .A1(resetn),
    .A2(_04682_),
    .ZN(_04683_)
  );
  AND2_X1 _39056_ (
    .A1(_04680_),
    .A2(_04683_),
    .ZN(_00266_)
  );
  AND2_X1 _39057_ (
    .A1(count_cycle[51]),
    .A2(_04679_),
    .ZN(_04684_)
  );
  INV_X1 _39058_ (
    .A(_04684_),
    .ZN(_04685_)
  );
  AND2_X1 _39059_ (
    .A1(_22204_),
    .A2(_04680_),
    .ZN(_04686_)
  );
  INV_X1 _39060_ (
    .A(_04686_),
    .ZN(_04687_)
  );
  AND2_X1 _39061_ (
    .A1(resetn),
    .A2(_04687_),
    .ZN(_04688_)
  );
  AND2_X1 _39062_ (
    .A1(_04685_),
    .A2(_04688_),
    .ZN(_00267_)
  );
  AND2_X1 _39063_ (
    .A1(count_cycle[52]),
    .A2(_04684_),
    .ZN(_04689_)
  );
  INV_X1 _39064_ (
    .A(_04689_),
    .ZN(_04690_)
  );
  AND2_X1 _39065_ (
    .A1(_22205_),
    .A2(_04685_),
    .ZN(_04691_)
  );
  INV_X1 _39066_ (
    .A(_04691_),
    .ZN(_04692_)
  );
  AND2_X1 _39067_ (
    .A1(resetn),
    .A2(_04692_),
    .ZN(_04693_)
  );
  AND2_X1 _39068_ (
    .A1(_04690_),
    .A2(_04693_),
    .ZN(_00268_)
  );
  AND2_X1 _39069_ (
    .A1(count_cycle[53]),
    .A2(_04689_),
    .ZN(_04694_)
  );
  INV_X1 _39070_ (
    .A(_04694_),
    .ZN(_04695_)
  );
  AND2_X1 _39071_ (
    .A1(_22206_),
    .A2(_04690_),
    .ZN(_04696_)
  );
  INV_X1 _39072_ (
    .A(_04696_),
    .ZN(_04697_)
  );
  AND2_X1 _39073_ (
    .A1(resetn),
    .A2(_04697_),
    .ZN(_04698_)
  );
  AND2_X1 _39074_ (
    .A1(_04695_),
    .A2(_04698_),
    .ZN(_00269_)
  );
  AND2_X1 _39075_ (
    .A1(count_cycle[54]),
    .A2(_04694_),
    .ZN(_04699_)
  );
  INV_X1 _39076_ (
    .A(_04699_),
    .ZN(_04700_)
  );
  AND2_X1 _39077_ (
    .A1(_22207_),
    .A2(_04695_),
    .ZN(_04701_)
  );
  INV_X1 _39078_ (
    .A(_04701_),
    .ZN(_04702_)
  );
  AND2_X1 _39079_ (
    .A1(resetn),
    .A2(_04702_),
    .ZN(_04703_)
  );
  AND2_X1 _39080_ (
    .A1(_04700_),
    .A2(_04703_),
    .ZN(_00270_)
  );
  AND2_X1 _39081_ (
    .A1(count_cycle[55]),
    .A2(_04699_),
    .ZN(_04704_)
  );
  INV_X1 _39082_ (
    .A(_04704_),
    .ZN(_04705_)
  );
  AND2_X1 _39083_ (
    .A1(_22208_),
    .A2(_04700_),
    .ZN(_04706_)
  );
  INV_X1 _39084_ (
    .A(_04706_),
    .ZN(_04707_)
  );
  AND2_X1 _39085_ (
    .A1(resetn),
    .A2(_04707_),
    .ZN(_04708_)
  );
  AND2_X1 _39086_ (
    .A1(_04705_),
    .A2(_04708_),
    .ZN(_00271_)
  );
  AND2_X1 _39087_ (
    .A1(count_cycle[56]),
    .A2(_04704_),
    .ZN(_04709_)
  );
  INV_X1 _39088_ (
    .A(_04709_),
    .ZN(_04710_)
  );
  AND2_X1 _39089_ (
    .A1(_22209_),
    .A2(_04705_),
    .ZN(_04711_)
  );
  INV_X1 _39090_ (
    .A(_04711_),
    .ZN(_04712_)
  );
  AND2_X1 _39091_ (
    .A1(resetn),
    .A2(_04712_),
    .ZN(_04713_)
  );
  AND2_X1 _39092_ (
    .A1(_04710_),
    .A2(_04713_),
    .ZN(_00272_)
  );
  AND2_X1 _39093_ (
    .A1(count_cycle[57]),
    .A2(_04709_),
    .ZN(_04714_)
  );
  INV_X1 _39094_ (
    .A(_04714_),
    .ZN(_04715_)
  );
  AND2_X1 _39095_ (
    .A1(_22210_),
    .A2(_04710_),
    .ZN(_04716_)
  );
  INV_X1 _39096_ (
    .A(_04716_),
    .ZN(_04717_)
  );
  AND2_X1 _39097_ (
    .A1(resetn),
    .A2(_04717_),
    .ZN(_04718_)
  );
  AND2_X1 _39098_ (
    .A1(_04715_),
    .A2(_04718_),
    .ZN(_00273_)
  );
  AND2_X1 _39099_ (
    .A1(count_cycle[58]),
    .A2(_04714_),
    .ZN(_04719_)
  );
  INV_X1 _39100_ (
    .A(_04719_),
    .ZN(_04720_)
  );
  AND2_X1 _39101_ (
    .A1(_22211_),
    .A2(_04715_),
    .ZN(_04721_)
  );
  INV_X1 _39102_ (
    .A(_04721_),
    .ZN(_04722_)
  );
  AND2_X1 _39103_ (
    .A1(resetn),
    .A2(_04722_),
    .ZN(_04723_)
  );
  AND2_X1 _39104_ (
    .A1(_04720_),
    .A2(_04723_),
    .ZN(_00274_)
  );
  AND2_X1 _39105_ (
    .A1(count_cycle[59]),
    .A2(_04719_),
    .ZN(_04724_)
  );
  INV_X1 _39106_ (
    .A(_04724_),
    .ZN(_04725_)
  );
  AND2_X1 _39107_ (
    .A1(_22212_),
    .A2(_04720_),
    .ZN(_04726_)
  );
  INV_X1 _39108_ (
    .A(_04726_),
    .ZN(_04727_)
  );
  AND2_X1 _39109_ (
    .A1(resetn),
    .A2(_04727_),
    .ZN(_04728_)
  );
  AND2_X1 _39110_ (
    .A1(_04725_),
    .A2(_04728_),
    .ZN(_00275_)
  );
  AND2_X1 _39111_ (
    .A1(count_cycle[60]),
    .A2(_04724_),
    .ZN(_04729_)
  );
  INV_X1 _39112_ (
    .A(_04729_),
    .ZN(_04730_)
  );
  AND2_X1 _39113_ (
    .A1(_22213_),
    .A2(_04725_),
    .ZN(_04731_)
  );
  INV_X1 _39114_ (
    .A(_04731_),
    .ZN(_04732_)
  );
  AND2_X1 _39115_ (
    .A1(resetn),
    .A2(_04732_),
    .ZN(_04733_)
  );
  AND2_X1 _39116_ (
    .A1(_04730_),
    .A2(_04733_),
    .ZN(_00276_)
  );
  AND2_X1 _39117_ (
    .A1(count_cycle[61]),
    .A2(_04729_),
    .ZN(_04734_)
  );
  INV_X1 _39118_ (
    .A(_04734_),
    .ZN(_04735_)
  );
  AND2_X1 _39119_ (
    .A1(_22214_),
    .A2(_04730_),
    .ZN(_04736_)
  );
  INV_X1 _39120_ (
    .A(_04736_),
    .ZN(_04737_)
  );
  AND2_X1 _39121_ (
    .A1(resetn),
    .A2(_04737_),
    .ZN(_04738_)
  );
  AND2_X1 _39122_ (
    .A1(_04735_),
    .A2(_04738_),
    .ZN(_00277_)
  );
  AND2_X1 _39123_ (
    .A1(count_cycle[62]),
    .A2(_04734_),
    .ZN(_04739_)
  );
  INV_X1 _39124_ (
    .A(_04739_),
    .ZN(_04740_)
  );
  AND2_X1 _39125_ (
    .A1(_22215_),
    .A2(_04735_),
    .ZN(_04741_)
  );
  INV_X1 _39126_ (
    .A(_04741_),
    .ZN(_04742_)
  );
  AND2_X1 _39127_ (
    .A1(resetn),
    .A2(_04742_),
    .ZN(_04743_)
  );
  AND2_X1 _39128_ (
    .A1(_04740_),
    .A2(_04743_),
    .ZN(_00278_)
  );
  AND2_X1 _39129_ (
    .A1(count_cycle[63]),
    .A2(_04739_),
    .ZN(_04744_)
  );
  INV_X1 _39130_ (
    .A(_04744_),
    .ZN(_04745_)
  );
  AND2_X1 _39131_ (
    .A1(_22216_),
    .A2(_04740_),
    .ZN(_04746_)
  );
  INV_X1 _39132_ (
    .A(_04746_),
    .ZN(_04747_)
  );
  AND2_X1 _39133_ (
    .A1(resetn),
    .A2(_04747_),
    .ZN(_04748_)
  );
  AND2_X1 _39134_ (
    .A1(_04745_),
    .A2(_04748_),
    .ZN(_00279_)
  );
  AND2_X1 _39135_ (
    .A1(_22288_),
    .A2(_22295_),
    .ZN(_04749_)
  );
  INV_X1 _39136_ (
    .A(_04749_),
    .ZN(_04750_)
  );
  AND2_X1 _39137_ (
    .A1(_22333_),
    .A2(_04750_),
    .ZN(_04751_)
  );
  INV_X1 _39138_ (
    .A(_04751_),
    .ZN(_04752_)
  );
  AND2_X1 _39139_ (
    .A1(_21199_),
    .A2(_04752_),
    .ZN(_04753_)
  );
  INV_X1 _39140_ (
    .A(_04753_),
    .ZN(_04754_)
  );
  AND2_X1 _39141_ (
    .A1(reg_pc[31]),
    .A2(_22335_),
    .ZN(_04755_)
  );
  INV_X1 _39142_ (
    .A(_04755_),
    .ZN(_04756_)
  );
  AND2_X1 _39143_ (
    .A1(\cpuregs[7] [31]),
    .A2(_00008_[2]),
    .ZN(_04757_)
  );
  INV_X1 _39144_ (
    .A(_04757_),
    .ZN(_04758_)
  );
  AND2_X1 _39145_ (
    .A1(\cpuregs[3] [31]),
    .A2(_22149_),
    .ZN(_04759_)
  );
  INV_X1 _39146_ (
    .A(_04759_),
    .ZN(_04760_)
  );
  AND2_X1 _39147_ (
    .A1(_04758_),
    .A2(_04760_),
    .ZN(_04761_)
  );
  INV_X1 _39148_ (
    .A(_04761_),
    .ZN(_04762_)
  );
  AND2_X1 _39149_ (
    .A1(_00008_[0]),
    .A2(_04762_),
    .ZN(_04763_)
  );
  INV_X1 _39150_ (
    .A(_04763_),
    .ZN(_04764_)
  );
  AND2_X1 _39151_ (
    .A1(_21361_),
    .A2(_22149_),
    .ZN(_04765_)
  );
  INV_X1 _39152_ (
    .A(_04765_),
    .ZN(_04766_)
  );
  AND2_X1 _39153_ (
    .A1(_21360_),
    .A2(_00008_[2]),
    .ZN(_04767_)
  );
  INV_X1 _39154_ (
    .A(_04767_),
    .ZN(_04768_)
  );
  AND2_X1 _39155_ (
    .A1(_04766_),
    .A2(_04768_),
    .ZN(_04769_)
  );
  AND2_X1 _39156_ (
    .A1(_22147_),
    .A2(_04769_),
    .ZN(_04770_)
  );
  INV_X1 _39157_ (
    .A(_04770_),
    .ZN(_04771_)
  );
  AND2_X1 _39158_ (
    .A1(\cpuregs[5] [31]),
    .A2(_00008_[2]),
    .ZN(_04772_)
  );
  INV_X1 _39159_ (
    .A(_04772_),
    .ZN(_04773_)
  );
  AND2_X1 _39160_ (
    .A1(\cpuregs[1] [31]),
    .A2(_22149_),
    .ZN(_04774_)
  );
  INV_X1 _39161_ (
    .A(_04774_),
    .ZN(_04775_)
  );
  AND2_X1 _39162_ (
    .A1(_04773_),
    .A2(_04775_),
    .ZN(_04776_)
  );
  INV_X1 _39163_ (
    .A(_04776_),
    .ZN(_04777_)
  );
  AND2_X1 _39164_ (
    .A1(_00008_[0]),
    .A2(_04777_),
    .ZN(_04778_)
  );
  INV_X1 _39165_ (
    .A(_04778_),
    .ZN(_04779_)
  );
  AND2_X1 _39166_ (
    .A1(\cpuregs[4] [31]),
    .A2(_00008_[2]),
    .ZN(_04780_)
  );
  INV_X1 _39167_ (
    .A(_04780_),
    .ZN(_04781_)
  );
  AND2_X1 _39168_ (
    .A1(\cpuregs[0] [31]),
    .A2(_22149_),
    .ZN(_04782_)
  );
  INV_X1 _39169_ (
    .A(_04782_),
    .ZN(_04783_)
  );
  AND2_X1 _39170_ (
    .A1(_04781_),
    .A2(_04783_),
    .ZN(_04784_)
  );
  INV_X1 _39171_ (
    .A(_04784_),
    .ZN(_04785_)
  );
  AND2_X1 _39172_ (
    .A1(_22147_),
    .A2(_04785_),
    .ZN(_04786_)
  );
  INV_X1 _39173_ (
    .A(_04786_),
    .ZN(_04787_)
  );
  AND2_X1 _39174_ (
    .A1(_04779_),
    .A2(_04787_),
    .ZN(_04788_)
  );
  AND2_X1 _39175_ (
    .A1(_00008_[1]),
    .A2(_04771_),
    .ZN(_04789_)
  );
  AND2_X1 _39176_ (
    .A1(_04764_),
    .A2(_04789_),
    .ZN(_04790_)
  );
  INV_X1 _39177_ (
    .A(_04790_),
    .ZN(_04791_)
  );
  AND2_X1 _39178_ (
    .A1(_22148_),
    .A2(_04788_),
    .ZN(_04792_)
  );
  INV_X1 _39179_ (
    .A(_04792_),
    .ZN(_04793_)
  );
  AND2_X1 _39180_ (
    .A1(_04791_),
    .A2(_04793_),
    .ZN(_04794_)
  );
  AND2_X1 _39181_ (
    .A1(_22150_),
    .A2(_04794_),
    .ZN(_04795_)
  );
  INV_X1 _39182_ (
    .A(_04795_),
    .ZN(_04796_)
  );
  AND2_X1 _39183_ (
    .A1(\cpuregs[13] [31]),
    .A2(_00008_[0]),
    .ZN(_04797_)
  );
  INV_X1 _39184_ (
    .A(_04797_),
    .ZN(_04798_)
  );
  AND2_X1 _39185_ (
    .A1(\cpuregs[12] [31]),
    .A2(_22147_),
    .ZN(_04799_)
  );
  INV_X1 _39186_ (
    .A(_04799_),
    .ZN(_04800_)
  );
  AND2_X1 _39187_ (
    .A1(_00008_[2]),
    .A2(_04800_),
    .ZN(_04801_)
  );
  AND2_X1 _39188_ (
    .A1(_04798_),
    .A2(_04801_),
    .ZN(_04802_)
  );
  INV_X1 _39189_ (
    .A(_04802_),
    .ZN(_04803_)
  );
  AND2_X1 _39190_ (
    .A1(\cpuregs[9] [31]),
    .A2(_00008_[0]),
    .ZN(_04804_)
  );
  INV_X1 _39191_ (
    .A(_04804_),
    .ZN(_04805_)
  );
  AND2_X1 _39192_ (
    .A1(\cpuregs[8] [31]),
    .A2(_22147_),
    .ZN(_04806_)
  );
  INV_X1 _39193_ (
    .A(_04806_),
    .ZN(_04807_)
  );
  AND2_X1 _39194_ (
    .A1(_22149_),
    .A2(_04807_),
    .ZN(_04808_)
  );
  AND2_X1 _39195_ (
    .A1(_04805_),
    .A2(_04808_),
    .ZN(_04809_)
  );
  INV_X1 _39196_ (
    .A(_04809_),
    .ZN(_04810_)
  );
  AND2_X1 _39197_ (
    .A1(_22148_),
    .A2(_04810_),
    .ZN(_04811_)
  );
  AND2_X1 _39198_ (
    .A1(_04803_),
    .A2(_04811_),
    .ZN(_04812_)
  );
  INV_X1 _39199_ (
    .A(_04812_),
    .ZN(_04813_)
  );
  AND2_X1 _39200_ (
    .A1(\cpuregs[15] [31]),
    .A2(_00008_[0]),
    .ZN(_04814_)
  );
  INV_X1 _39201_ (
    .A(_04814_),
    .ZN(_04815_)
  );
  AND2_X1 _39202_ (
    .A1(\cpuregs[14] [31]),
    .A2(_22147_),
    .ZN(_04816_)
  );
  INV_X1 _39203_ (
    .A(_04816_),
    .ZN(_04817_)
  );
  AND2_X1 _39204_ (
    .A1(_00008_[2]),
    .A2(_04817_),
    .ZN(_04818_)
  );
  AND2_X1 _39205_ (
    .A1(_04815_),
    .A2(_04818_),
    .ZN(_04819_)
  );
  INV_X1 _39206_ (
    .A(_04819_),
    .ZN(_04820_)
  );
  AND2_X1 _39207_ (
    .A1(\cpuregs[11] [31]),
    .A2(_00008_[0]),
    .ZN(_04821_)
  );
  INV_X1 _39208_ (
    .A(_04821_),
    .ZN(_04822_)
  );
  AND2_X1 _39209_ (
    .A1(\cpuregs[10] [31]),
    .A2(_22147_),
    .ZN(_04823_)
  );
  INV_X1 _39210_ (
    .A(_04823_),
    .ZN(_04824_)
  );
  AND2_X1 _39211_ (
    .A1(_22149_),
    .A2(_04824_),
    .ZN(_04825_)
  );
  AND2_X1 _39212_ (
    .A1(_04822_),
    .A2(_04825_),
    .ZN(_04826_)
  );
  INV_X1 _39213_ (
    .A(_04826_),
    .ZN(_04827_)
  );
  AND2_X1 _39214_ (
    .A1(_00008_[1]),
    .A2(_04827_),
    .ZN(_04828_)
  );
  AND2_X1 _39215_ (
    .A1(_04820_),
    .A2(_04828_),
    .ZN(_04829_)
  );
  INV_X1 _39216_ (
    .A(_04829_),
    .ZN(_04830_)
  );
  AND2_X1 _39217_ (
    .A1(_04813_),
    .A2(_04830_),
    .ZN(_04831_)
  );
  INV_X1 _39218_ (
    .A(_04831_),
    .ZN(_04832_)
  );
  AND2_X1 _39219_ (
    .A1(_00008_[3]),
    .A2(_04832_),
    .ZN(_04833_)
  );
  INV_X1 _39220_ (
    .A(_04833_),
    .ZN(_04834_)
  );
  AND2_X1 _39221_ (
    .A1(_04796_),
    .A2(_04834_),
    .ZN(_04835_)
  );
  AND2_X1 _39222_ (
    .A1(_22151_),
    .A2(_04835_),
    .ZN(_04836_)
  );
  INV_X1 _39223_ (
    .A(_04836_),
    .ZN(_04837_)
  );
  AND2_X1 _39224_ (
    .A1(\cpuregs[26] [31]),
    .A2(_22149_),
    .ZN(_04838_)
  );
  INV_X1 _39225_ (
    .A(_04838_),
    .ZN(_04839_)
  );
  AND2_X1 _39226_ (
    .A1(\cpuregs[30] [31]),
    .A2(_00008_[2]),
    .ZN(_04840_)
  );
  INV_X1 _39227_ (
    .A(_04840_),
    .ZN(_04841_)
  );
  AND2_X1 _39228_ (
    .A1(_22147_),
    .A2(_04841_),
    .ZN(_04842_)
  );
  AND2_X1 _39229_ (
    .A1(_04839_),
    .A2(_04842_),
    .ZN(_04843_)
  );
  INV_X1 _39230_ (
    .A(_04843_),
    .ZN(_04844_)
  );
  AND2_X1 _39231_ (
    .A1(\cpuregs[31] [31]),
    .A2(_00008_[2]),
    .ZN(_04845_)
  );
  INV_X1 _39232_ (
    .A(_04845_),
    .ZN(_04846_)
  );
  AND2_X1 _39233_ (
    .A1(\cpuregs[27] [31]),
    .A2(_22149_),
    .ZN(_04847_)
  );
  INV_X1 _39234_ (
    .A(_04847_),
    .ZN(_04848_)
  );
  AND2_X1 _39235_ (
    .A1(_00008_[0]),
    .A2(_04848_),
    .ZN(_04849_)
  );
  AND2_X1 _39236_ (
    .A1(_04846_),
    .A2(_04849_),
    .ZN(_04850_)
  );
  INV_X1 _39237_ (
    .A(_04850_),
    .ZN(_04851_)
  );
  AND2_X1 _39238_ (
    .A1(_04844_),
    .A2(_04851_),
    .ZN(_04852_)
  );
  INV_X1 _39239_ (
    .A(_04852_),
    .ZN(_04853_)
  );
  AND2_X1 _39240_ (
    .A1(_00008_[3]),
    .A2(_04853_),
    .ZN(_04854_)
  );
  INV_X1 _39241_ (
    .A(_04854_),
    .ZN(_04855_)
  );
  AND2_X1 _39242_ (
    .A1(\cpuregs[18] [31]),
    .A2(_22149_),
    .ZN(_04856_)
  );
  INV_X1 _39243_ (
    .A(_04856_),
    .ZN(_04857_)
  );
  AND2_X1 _39244_ (
    .A1(\cpuregs[22] [31]),
    .A2(_00008_[2]),
    .ZN(_04858_)
  );
  INV_X1 _39245_ (
    .A(_04858_),
    .ZN(_04859_)
  );
  AND2_X1 _39246_ (
    .A1(_22147_),
    .A2(_04859_),
    .ZN(_04860_)
  );
  AND2_X1 _39247_ (
    .A1(_04857_),
    .A2(_04860_),
    .ZN(_04861_)
  );
  INV_X1 _39248_ (
    .A(_04861_),
    .ZN(_04862_)
  );
  AND2_X1 _39249_ (
    .A1(\cpuregs[19] [31]),
    .A2(_22149_),
    .ZN(_04863_)
  );
  INV_X1 _39250_ (
    .A(_04863_),
    .ZN(_04864_)
  );
  AND2_X1 _39251_ (
    .A1(\cpuregs[23] [31]),
    .A2(_00008_[2]),
    .ZN(_04865_)
  );
  INV_X1 _39252_ (
    .A(_04865_),
    .ZN(_04866_)
  );
  AND2_X1 _39253_ (
    .A1(_00008_[0]),
    .A2(_04866_),
    .ZN(_04867_)
  );
  AND2_X1 _39254_ (
    .A1(_04864_),
    .A2(_04867_),
    .ZN(_04868_)
  );
  INV_X1 _39255_ (
    .A(_04868_),
    .ZN(_04869_)
  );
  AND2_X1 _39256_ (
    .A1(_04862_),
    .A2(_04869_),
    .ZN(_04870_)
  );
  INV_X1 _39257_ (
    .A(_04870_),
    .ZN(_04871_)
  );
  AND2_X1 _39258_ (
    .A1(_22150_),
    .A2(_04871_),
    .ZN(_04872_)
  );
  INV_X1 _39259_ (
    .A(_04872_),
    .ZN(_04873_)
  );
  AND2_X1 _39260_ (
    .A1(\cpuregs[24] [31]),
    .A2(_22149_),
    .ZN(_04874_)
  );
  INV_X1 _39261_ (
    .A(_04874_),
    .ZN(_04875_)
  );
  AND2_X1 _39262_ (
    .A1(\cpuregs[28] [31]),
    .A2(_00008_[2]),
    .ZN(_04876_)
  );
  INV_X1 _39263_ (
    .A(_04876_),
    .ZN(_04877_)
  );
  AND2_X1 _39264_ (
    .A1(_22147_),
    .A2(_04877_),
    .ZN(_04878_)
  );
  AND2_X1 _39265_ (
    .A1(_04875_),
    .A2(_04878_),
    .ZN(_04879_)
  );
  INV_X1 _39266_ (
    .A(_04879_),
    .ZN(_04880_)
  );
  AND2_X1 _39267_ (
    .A1(\cpuregs[29] [31]),
    .A2(_00008_[2]),
    .ZN(_04881_)
  );
  INV_X1 _39268_ (
    .A(_04881_),
    .ZN(_04882_)
  );
  AND2_X1 _39269_ (
    .A1(\cpuregs[25] [31]),
    .A2(_22149_),
    .ZN(_04883_)
  );
  INV_X1 _39270_ (
    .A(_04883_),
    .ZN(_04884_)
  );
  AND2_X1 _39271_ (
    .A1(_00008_[0]),
    .A2(_04884_),
    .ZN(_04885_)
  );
  AND2_X1 _39272_ (
    .A1(_04882_),
    .A2(_04885_),
    .ZN(_04886_)
  );
  INV_X1 _39273_ (
    .A(_04886_),
    .ZN(_04887_)
  );
  AND2_X1 _39274_ (
    .A1(_04880_),
    .A2(_04887_),
    .ZN(_04888_)
  );
  AND2_X1 _39275_ (
    .A1(\cpuregs[16] [31]),
    .A2(_22149_),
    .ZN(_04889_)
  );
  INV_X1 _39276_ (
    .A(_04889_),
    .ZN(_04890_)
  );
  AND2_X1 _39277_ (
    .A1(\cpuregs[20] [31]),
    .A2(_00008_[2]),
    .ZN(_04891_)
  );
  INV_X1 _39278_ (
    .A(_04891_),
    .ZN(_04892_)
  );
  AND2_X1 _39279_ (
    .A1(_22147_),
    .A2(_04892_),
    .ZN(_04893_)
  );
  AND2_X1 _39280_ (
    .A1(_04890_),
    .A2(_04893_),
    .ZN(_04894_)
  );
  INV_X1 _39281_ (
    .A(_04894_),
    .ZN(_04895_)
  );
  AND2_X1 _39282_ (
    .A1(\cpuregs[17] [31]),
    .A2(_22149_),
    .ZN(_04896_)
  );
  INV_X1 _39283_ (
    .A(_04896_),
    .ZN(_04897_)
  );
  AND2_X1 _39284_ (
    .A1(\cpuregs[21] [31]),
    .A2(_00008_[2]),
    .ZN(_04898_)
  );
  INV_X1 _39285_ (
    .A(_04898_),
    .ZN(_04899_)
  );
  AND2_X1 _39286_ (
    .A1(_00008_[0]),
    .A2(_04899_),
    .ZN(_04900_)
  );
  AND2_X1 _39287_ (
    .A1(_04897_),
    .A2(_04900_),
    .ZN(_04901_)
  );
  INV_X1 _39288_ (
    .A(_04901_),
    .ZN(_04902_)
  );
  AND2_X1 _39289_ (
    .A1(_00008_[3]),
    .A2(_04888_),
    .ZN(_04903_)
  );
  INV_X1 _39290_ (
    .A(_04903_),
    .ZN(_04904_)
  );
  AND2_X1 _39291_ (
    .A1(_22150_),
    .A2(_04902_),
    .ZN(_04905_)
  );
  AND2_X1 _39292_ (
    .A1(_04895_),
    .A2(_04905_),
    .ZN(_04906_)
  );
  INV_X1 _39293_ (
    .A(_04906_),
    .ZN(_04907_)
  );
  AND2_X1 _39294_ (
    .A1(_04904_),
    .A2(_04907_),
    .ZN(_04908_)
  );
  INV_X1 _39295_ (
    .A(_04908_),
    .ZN(_04909_)
  );
  AND2_X1 _39296_ (
    .A1(_00008_[1]),
    .A2(_04873_),
    .ZN(_04910_)
  );
  AND2_X1 _39297_ (
    .A1(_04855_),
    .A2(_04910_),
    .ZN(_04911_)
  );
  INV_X1 _39298_ (
    .A(_04911_),
    .ZN(_04912_)
  );
  AND2_X1 _39299_ (
    .A1(_22148_),
    .A2(_04909_),
    .ZN(_04913_)
  );
  INV_X1 _39300_ (
    .A(_04913_),
    .ZN(_04914_)
  );
  AND2_X1 _39301_ (
    .A1(_00008_[4]),
    .A2(_04912_),
    .ZN(_04915_)
  );
  AND2_X1 _39302_ (
    .A1(_04914_),
    .A2(_04915_),
    .ZN(_04916_)
  );
  INV_X1 _39303_ (
    .A(_04916_),
    .ZN(_04917_)
  );
  AND2_X1 _39304_ (
    .A1(_22546_),
    .A2(_04917_),
    .ZN(_04918_)
  );
  AND2_X1 _39305_ (
    .A1(_04837_),
    .A2(_04918_),
    .ZN(_04919_)
  );
  INV_X1 _39306_ (
    .A(_04919_),
    .ZN(_04920_)
  );
  AND2_X1 _39307_ (
    .A1(_04756_),
    .A2(_04920_),
    .ZN(_04921_)
  );
  INV_X1 _39308_ (
    .A(_04921_),
    .ZN(_04922_)
  );
  AND2_X1 _39309_ (
    .A1(_22271_),
    .A2(_04922_),
    .ZN(_04923_)
  );
  INV_X1 _39310_ (
    .A(_04923_),
    .ZN(_04924_)
  );
  AND2_X1 _39311_ (
    .A1(_22573_),
    .A2(_02028_),
    .ZN(_04925_)
  );
  INV_X1 _39312_ (
    .A(_04925_),
    .ZN(_04926_)
  );
  AND2_X1 _39313_ (
    .A1(reg_op1[30]),
    .A2(_22285_),
    .ZN(_04927_)
  );
  AND2_X1 _39314_ (
    .A1(_22572_),
    .A2(_04927_),
    .ZN(_04928_)
  );
  INV_X1 _39315_ (
    .A(_04928_),
    .ZN(_04929_)
  );
  AND2_X1 _39316_ (
    .A1(_04926_),
    .A2(_04929_),
    .ZN(_04930_)
  );
  INV_X1 _39317_ (
    .A(_04930_),
    .ZN(_04931_)
  );
  AND2_X1 _39318_ (
    .A1(_22295_),
    .A2(_04931_),
    .ZN(_04932_)
  );
  INV_X1 _39319_ (
    .A(_04932_),
    .ZN(_04933_)
  );
  AND2_X1 _39320_ (
    .A1(_04751_),
    .A2(_04933_),
    .ZN(_04934_)
  );
  AND2_X1 _39321_ (
    .A1(_04924_),
    .A2(_04934_),
    .ZN(_04935_)
  );
  AND2_X1 _39322_ (
    .A1(_02448_),
    .A2(_02454_),
    .ZN(_04936_)
  );
  INV_X1 _39323_ (
    .A(_04936_),
    .ZN(_04937_)
  );
  AND2_X1 _39324_ (
    .A1(reg_op1[31]),
    .A2(_21978_),
    .ZN(_04938_)
  );
  INV_X1 _39325_ (
    .A(_04938_),
    .ZN(_04939_)
  );
  AND2_X1 _39326_ (
    .A1(_21199_),
    .A2(decoded_imm[31]),
    .ZN(_04940_)
  );
  INV_X1 _39327_ (
    .A(_04940_),
    .ZN(_04941_)
  );
  AND2_X1 _39328_ (
    .A1(_21199_),
    .A2(_21978_),
    .ZN(_04942_)
  );
  INV_X1 _39329_ (
    .A(_04942_),
    .ZN(_04943_)
  );
  AND2_X1 _39330_ (
    .A1(reg_op1[31]),
    .A2(decoded_imm[31]),
    .ZN(_04944_)
  );
  INV_X1 _39331_ (
    .A(_04944_),
    .ZN(_04945_)
  );
  AND2_X1 _39332_ (
    .A1(_04939_),
    .A2(_04941_),
    .ZN(_04946_)
  );
  AND2_X1 _39333_ (
    .A1(_04943_),
    .A2(_04945_),
    .ZN(_04947_)
  );
  AND2_X1 _39334_ (
    .A1(_04937_),
    .A2(_04947_),
    .ZN(_04948_)
  );
  INV_X1 _39335_ (
    .A(_04948_),
    .ZN(_04949_)
  );
  AND2_X1 _39336_ (
    .A1(_04936_),
    .A2(_04946_),
    .ZN(_04950_)
  );
  INV_X1 _39337_ (
    .A(_04950_),
    .ZN(_04951_)
  );
  AND2_X1 _39338_ (
    .A1(_22559_),
    .A2(_04951_),
    .ZN(_04952_)
  );
  AND2_X1 _39339_ (
    .A1(_04949_),
    .A2(_04952_),
    .ZN(_04953_)
  );
  INV_X1 _39340_ (
    .A(_04953_),
    .ZN(_04954_)
  );
  AND2_X1 _39341_ (
    .A1(_04935_),
    .A2(_04954_),
    .ZN(_04955_)
  );
  INV_X1 _39342_ (
    .A(_04955_),
    .ZN(_04956_)
  );
  AND2_X1 _39343_ (
    .A1(_04754_),
    .A2(_04956_),
    .ZN(_00280_)
  );
  AND2_X1 _39344_ (
    .A1(_22026_),
    .A2(_22060_),
    .ZN(_04957_)
  );
  AND2_X1 _39345_ (
    .A1(_22269_),
    .A2(_04957_),
    .ZN(_04958_)
  );
  INV_X1 _39346_ (
    .A(_04958_),
    .ZN(_04959_)
  );
  AND2_X1 _39347_ (
    .A1(_22272_),
    .A2(_04959_),
    .ZN(_04960_)
  );
  INV_X1 _39348_ (
    .A(_04960_),
    .ZN(_04961_)
  );
  AND2_X1 _39349_ (
    .A1(resetn),
    .A2(_04961_),
    .ZN(_04962_)
  );
  INV_X1 _39350_ (
    .A(_04962_),
    .ZN(_04963_)
  );
  AND2_X1 _39351_ (
    .A1(_21293_),
    .A2(_22070_),
    .ZN(_04964_)
  );
  INV_X1 _39352_ (
    .A(_04964_),
    .ZN(_04965_)
  );
  AND2_X1 _39353_ (
    .A1(_22271_),
    .A2(_04965_),
    .ZN(_04966_)
  );
  INV_X1 _39354_ (
    .A(_04966_),
    .ZN(_04967_)
  );
  AND2_X1 _39355_ (
    .A1(decoded_imm[0]),
    .A2(_04966_),
    .ZN(_04968_)
  );
  INV_X1 _39356_ (
    .A(_04968_),
    .ZN(_04969_)
  );
  AND2_X1 _39357_ (
    .A1(_21282_),
    .A2(_21283_),
    .ZN(_04970_)
  );
  AND2_X1 _39358_ (
    .A1(_21284_),
    .A2(_21285_),
    .ZN(_04971_)
  );
  AND2_X1 _39359_ (
    .A1(_22015_),
    .A2(_04971_),
    .ZN(_04972_)
  );
  AND2_X1 _39360_ (
    .A1(_04970_),
    .A2(_04972_),
    .ZN(_04973_)
  );
  INV_X1 _39361_ (
    .A(_04973_),
    .ZN(_04974_)
  );
  AND2_X1 _39362_ (
    .A1(_21889_),
    .A2(_00007_[2]),
    .ZN(_04975_)
  );
  INV_X1 _39363_ (
    .A(_04975_),
    .ZN(_04976_)
  );
  AND2_X1 _39364_ (
    .A1(_21833_),
    .A2(_22077_),
    .ZN(_04977_)
  );
  INV_X1 _39365_ (
    .A(_04977_),
    .ZN(_04978_)
  );
  AND2_X1 _39366_ (
    .A1(_00007_[0]),
    .A2(_04978_),
    .ZN(_04979_)
  );
  AND2_X1 _39367_ (
    .A1(_04976_),
    .A2(_04979_),
    .ZN(_04980_)
  );
  INV_X1 _39368_ (
    .A(_04980_),
    .ZN(_04981_)
  );
  AND2_X1 _39369_ (
    .A1(_21567_),
    .A2(_22077_),
    .ZN(_04982_)
  );
  INV_X1 _39370_ (
    .A(_04982_),
    .ZN(_04983_)
  );
  AND2_X1 _39371_ (
    .A1(_21905_),
    .A2(_00007_[2]),
    .ZN(_04984_)
  );
  INV_X1 _39372_ (
    .A(_04984_),
    .ZN(_04985_)
  );
  AND2_X1 _39373_ (
    .A1(_04983_),
    .A2(_04985_),
    .ZN(_04986_)
  );
  AND2_X1 _39374_ (
    .A1(_22152_),
    .A2(_04986_),
    .ZN(_04987_)
  );
  INV_X1 _39375_ (
    .A(_04987_),
    .ZN(_04988_)
  );
  AND2_X1 _39376_ (
    .A1(_04981_),
    .A2(_04988_),
    .ZN(_04989_)
  );
  AND2_X1 _39377_ (
    .A1(_22078_),
    .A2(_04989_),
    .ZN(_04990_)
  );
  INV_X1 _39378_ (
    .A(_04990_),
    .ZN(_04991_)
  );
  AND2_X1 _39379_ (
    .A1(_21865_),
    .A2(_22077_),
    .ZN(_04992_)
  );
  INV_X1 _39380_ (
    .A(_04992_),
    .ZN(_04993_)
  );
  AND2_X1 _39381_ (
    .A1(_21849_),
    .A2(_00007_[2]),
    .ZN(_04994_)
  );
  INV_X1 _39382_ (
    .A(_04994_),
    .ZN(_04995_)
  );
  AND2_X1 _39383_ (
    .A1(_04993_),
    .A2(_04995_),
    .ZN(_04996_)
  );
  AND2_X1 _39384_ (
    .A1(_22152_),
    .A2(_04996_),
    .ZN(_04997_)
  );
  INV_X1 _39385_ (
    .A(_04997_),
    .ZN(_04998_)
  );
  AND2_X1 _39386_ (
    .A1(_21937_),
    .A2(_00007_[2]),
    .ZN(_04999_)
  );
  INV_X1 _39387_ (
    .A(_04999_),
    .ZN(_05000_)
  );
  AND2_X1 _39388_ (
    .A1(_21921_),
    .A2(_22077_),
    .ZN(_05001_)
  );
  INV_X1 _39389_ (
    .A(_05001_),
    .ZN(_05002_)
  );
  AND2_X1 _39390_ (
    .A1(_00007_[0]),
    .A2(_05002_),
    .ZN(_05003_)
  );
  AND2_X1 _39391_ (
    .A1(_05000_),
    .A2(_05003_),
    .ZN(_05004_)
  );
  INV_X1 _39392_ (
    .A(_05004_),
    .ZN(_05005_)
  );
  AND2_X1 _39393_ (
    .A1(_04998_),
    .A2(_05005_),
    .ZN(_05006_)
  );
  AND2_X1 _39394_ (
    .A1(_00007_[1]),
    .A2(_05006_),
    .ZN(_05007_)
  );
  INV_X1 _39395_ (
    .A(_05007_),
    .ZN(_05008_)
  );
  AND2_X1 _39396_ (
    .A1(_00007_[3]),
    .A2(_04991_),
    .ZN(_05009_)
  );
  AND2_X1 _39397_ (
    .A1(_05008_),
    .A2(_05009_),
    .ZN(_05010_)
  );
  INV_X1 _39398_ (
    .A(_05010_),
    .ZN(_05011_)
  );
  AND2_X1 _39399_ (
    .A1(_21590_),
    .A2(_22077_),
    .ZN(_05012_)
  );
  INV_X1 _39400_ (
    .A(_05012_),
    .ZN(_05013_)
  );
  AND2_X1 _39401_ (
    .A1(_21408_),
    .A2(_00007_[2]),
    .ZN(_05014_)
  );
  INV_X1 _39402_ (
    .A(_05014_),
    .ZN(_05015_)
  );
  AND2_X1 _39403_ (
    .A1(_21436_),
    .A2(_22077_),
    .ZN(_05016_)
  );
  INV_X1 _39404_ (
    .A(_05016_),
    .ZN(_05017_)
  );
  AND2_X1 _39405_ (
    .A1(_21647_),
    .A2(_00007_[2]),
    .ZN(_05018_)
  );
  INV_X1 _39406_ (
    .A(_05018_),
    .ZN(_05019_)
  );
  AND2_X1 _39407_ (
    .A1(_05017_),
    .A2(_05019_),
    .ZN(_05020_)
  );
  AND2_X1 _39408_ (
    .A1(_21370_),
    .A2(_00007_[2]),
    .ZN(_05021_)
  );
  INV_X1 _39409_ (
    .A(_05021_),
    .ZN(_05022_)
  );
  AND2_X1 _39410_ (
    .A1(_21616_),
    .A2(_22077_),
    .ZN(_05023_)
  );
  INV_X1 _39411_ (
    .A(_05023_),
    .ZN(_05024_)
  );
  AND2_X1 _39412_ (
    .A1(_21458_),
    .A2(_22077_),
    .ZN(_05025_)
  );
  INV_X1 _39413_ (
    .A(_05025_),
    .ZN(_05026_)
  );
  AND2_X1 _39414_ (
    .A1(_21757_),
    .A2(_00007_[2]),
    .ZN(_05027_)
  );
  INV_X1 _39415_ (
    .A(_05027_),
    .ZN(_05028_)
  );
  AND2_X1 _39416_ (
    .A1(_00007_[0]),
    .A2(_05024_),
    .ZN(_05029_)
  );
  AND2_X1 _39417_ (
    .A1(_05022_),
    .A2(_05029_),
    .ZN(_05030_)
  );
  INV_X1 _39418_ (
    .A(_05030_),
    .ZN(_05031_)
  );
  AND2_X1 _39419_ (
    .A1(_22152_),
    .A2(_05013_),
    .ZN(_05032_)
  );
  AND2_X1 _39420_ (
    .A1(_05015_),
    .A2(_05032_),
    .ZN(_05033_)
  );
  INV_X1 _39421_ (
    .A(_05033_),
    .ZN(_05034_)
  );
  AND2_X1 _39422_ (
    .A1(_05031_),
    .A2(_05034_),
    .ZN(_05035_)
  );
  AND2_X1 _39423_ (
    .A1(_00007_[1]),
    .A2(_05035_),
    .ZN(_05036_)
  );
  INV_X1 _39424_ (
    .A(_05036_),
    .ZN(_05037_)
  );
  AND2_X1 _39425_ (
    .A1(_00007_[0]),
    .A2(_05026_),
    .ZN(_05038_)
  );
  AND2_X1 _39426_ (
    .A1(_05028_),
    .A2(_05038_),
    .ZN(_05039_)
  );
  INV_X1 _39427_ (
    .A(_05039_),
    .ZN(_05040_)
  );
  AND2_X1 _39428_ (
    .A1(_22152_),
    .A2(_05020_),
    .ZN(_05041_)
  );
  INV_X1 _39429_ (
    .A(_05041_),
    .ZN(_05042_)
  );
  AND2_X1 _39430_ (
    .A1(_05040_),
    .A2(_05042_),
    .ZN(_05043_)
  );
  AND2_X1 _39431_ (
    .A1(_22078_),
    .A2(_05043_),
    .ZN(_05044_)
  );
  INV_X1 _39432_ (
    .A(_05044_),
    .ZN(_05045_)
  );
  AND2_X1 _39433_ (
    .A1(_05037_),
    .A2(_05045_),
    .ZN(_05046_)
  );
  AND2_X1 _39434_ (
    .A1(_22109_),
    .A2(_05046_),
    .ZN(_05047_)
  );
  INV_X1 _39435_ (
    .A(_05047_),
    .ZN(_05048_)
  );
  AND2_X1 _39436_ (
    .A1(_05011_),
    .A2(_05048_),
    .ZN(_05049_)
  );
  AND2_X1 _39437_ (
    .A1(\cpuregs[13] [0]),
    .A2(_22078_),
    .ZN(_05050_)
  );
  INV_X1 _39438_ (
    .A(_05050_),
    .ZN(_05051_)
  );
  AND2_X1 _39439_ (
    .A1(\cpuregs[15] [0]),
    .A2(_00007_[1]),
    .ZN(_05052_)
  );
  INV_X1 _39440_ (
    .A(_05052_),
    .ZN(_05053_)
  );
  AND2_X1 _39441_ (
    .A1(_00007_[2]),
    .A2(_05053_),
    .ZN(_05054_)
  );
  AND2_X1 _39442_ (
    .A1(_05051_),
    .A2(_05054_),
    .ZN(_05055_)
  );
  INV_X1 _39443_ (
    .A(_05055_),
    .ZN(_05056_)
  );
  AND2_X1 _39444_ (
    .A1(\cpuregs[9] [0]),
    .A2(_22078_),
    .ZN(_05057_)
  );
  INV_X1 _39445_ (
    .A(_05057_),
    .ZN(_05058_)
  );
  AND2_X1 _39446_ (
    .A1(\cpuregs[11] [0]),
    .A2(_00007_[1]),
    .ZN(_05059_)
  );
  INV_X1 _39447_ (
    .A(_05059_),
    .ZN(_05060_)
  );
  AND2_X1 _39448_ (
    .A1(_22077_),
    .A2(_05060_),
    .ZN(_05061_)
  );
  AND2_X1 _39449_ (
    .A1(_05058_),
    .A2(_05061_),
    .ZN(_05062_)
  );
  INV_X1 _39450_ (
    .A(_05062_),
    .ZN(_05063_)
  );
  AND2_X1 _39451_ (
    .A1(_00007_[0]),
    .A2(_05063_),
    .ZN(_05064_)
  );
  AND2_X1 _39452_ (
    .A1(_05056_),
    .A2(_05064_),
    .ZN(_05065_)
  );
  INV_X1 _39453_ (
    .A(_05065_),
    .ZN(_05066_)
  );
  AND2_X1 _39454_ (
    .A1(\cpuregs[12] [0]),
    .A2(_22078_),
    .ZN(_05067_)
  );
  INV_X1 _39455_ (
    .A(_05067_),
    .ZN(_05068_)
  );
  AND2_X1 _39456_ (
    .A1(\cpuregs[14] [0]),
    .A2(_00007_[1]),
    .ZN(_05069_)
  );
  INV_X1 _39457_ (
    .A(_05069_),
    .ZN(_05070_)
  );
  AND2_X1 _39458_ (
    .A1(_00007_[2]),
    .A2(_05070_),
    .ZN(_05071_)
  );
  AND2_X1 _39459_ (
    .A1(_05068_),
    .A2(_05071_),
    .ZN(_05072_)
  );
  INV_X1 _39460_ (
    .A(_05072_),
    .ZN(_05073_)
  );
  AND2_X1 _39461_ (
    .A1(\cpuregs[8] [0]),
    .A2(_22078_),
    .ZN(_05074_)
  );
  INV_X1 _39462_ (
    .A(_05074_),
    .ZN(_05075_)
  );
  AND2_X1 _39463_ (
    .A1(\cpuregs[10] [0]),
    .A2(_00007_[1]),
    .ZN(_05076_)
  );
  INV_X1 _39464_ (
    .A(_05076_),
    .ZN(_05077_)
  );
  AND2_X1 _39465_ (
    .A1(_22077_),
    .A2(_05077_),
    .ZN(_05078_)
  );
  AND2_X1 _39466_ (
    .A1(_05075_),
    .A2(_05078_),
    .ZN(_05079_)
  );
  INV_X1 _39467_ (
    .A(_05079_),
    .ZN(_05080_)
  );
  AND2_X1 _39468_ (
    .A1(_22152_),
    .A2(_05080_),
    .ZN(_05081_)
  );
  AND2_X1 _39469_ (
    .A1(_05073_),
    .A2(_05081_),
    .ZN(_05082_)
  );
  INV_X1 _39470_ (
    .A(_05082_),
    .ZN(_05083_)
  );
  AND2_X1 _39471_ (
    .A1(_05066_),
    .A2(_05083_),
    .ZN(_05084_)
  );
  INV_X1 _39472_ (
    .A(_05084_),
    .ZN(_05085_)
  );
  AND2_X1 _39473_ (
    .A1(_00007_[3]),
    .A2(_05085_),
    .ZN(_05086_)
  );
  INV_X1 _39474_ (
    .A(_05086_),
    .ZN(_05087_)
  );
  AND2_X1 _39475_ (
    .A1(_21537_),
    .A2(_22077_),
    .ZN(_05088_)
  );
  INV_X1 _39476_ (
    .A(_05088_),
    .ZN(_05089_)
  );
  AND2_X1 _39477_ (
    .A1(_21804_),
    .A2(_00007_[2]),
    .ZN(_05090_)
  );
  INV_X1 _39478_ (
    .A(_05090_),
    .ZN(_05091_)
  );
  AND2_X1 _39479_ (
    .A1(_22152_),
    .A2(_05091_),
    .ZN(_05092_)
  );
  AND2_X1 _39480_ (
    .A1(_05089_),
    .A2(_05092_),
    .ZN(_05093_)
  );
  INV_X1 _39481_ (
    .A(_05093_),
    .ZN(_05094_)
  );
  AND2_X1 _39482_ (
    .A1(_21779_),
    .A2(_00007_[2]),
    .ZN(_05095_)
  );
  INV_X1 _39483_ (
    .A(_05095_),
    .ZN(_05096_)
  );
  AND2_X1 _39484_ (
    .A1(_21487_),
    .A2(_22077_),
    .ZN(_05097_)
  );
  INV_X1 _39485_ (
    .A(_05097_),
    .ZN(_05098_)
  );
  AND2_X1 _39486_ (
    .A1(_00007_[0]),
    .A2(_05098_),
    .ZN(_05099_)
  );
  AND2_X1 _39487_ (
    .A1(_05096_),
    .A2(_05099_),
    .ZN(_05100_)
  );
  INV_X1 _39488_ (
    .A(_05100_),
    .ZN(_05101_)
  );
  AND2_X1 _39489_ (
    .A1(_05094_),
    .A2(_05101_),
    .ZN(_05102_)
  );
  AND2_X1 _39490_ (
    .A1(_21669_),
    .A2(_00007_[2]),
    .ZN(_05103_)
  );
  INV_X1 _39491_ (
    .A(_05103_),
    .ZN(_05104_)
  );
  AND2_X1 _39492_ (
    .A1(_21953_),
    .A2(_22077_),
    .ZN(_05105_)
  );
  INV_X1 _39493_ (
    .A(_05105_),
    .ZN(_05106_)
  );
  AND2_X1 _39494_ (
    .A1(_05104_),
    .A2(_05106_),
    .ZN(_05107_)
  );
  AND2_X1 _39495_ (
    .A1(_22152_),
    .A2(_05107_),
    .ZN(_05108_)
  );
  INV_X1 _39496_ (
    .A(_05108_),
    .ZN(_05109_)
  );
  AND2_X1 _39497_ (
    .A1(_21732_),
    .A2(_00007_[2]),
    .ZN(_05110_)
  );
  INV_X1 _39498_ (
    .A(_05110_),
    .ZN(_05111_)
  );
  AND2_X1 _39499_ (
    .A1(_21512_),
    .A2(_22077_),
    .ZN(_05112_)
  );
  INV_X1 _39500_ (
    .A(_05112_),
    .ZN(_05113_)
  );
  AND2_X1 _39501_ (
    .A1(_00007_[0]),
    .A2(_05113_),
    .ZN(_05114_)
  );
  AND2_X1 _39502_ (
    .A1(_05111_),
    .A2(_05114_),
    .ZN(_05115_)
  );
  INV_X1 _39503_ (
    .A(_05115_),
    .ZN(_05116_)
  );
  AND2_X1 _39504_ (
    .A1(_05109_),
    .A2(_05116_),
    .ZN(_05117_)
  );
  AND2_X1 _39505_ (
    .A1(_00007_[1]),
    .A2(_05102_),
    .ZN(_05118_)
  );
  INV_X1 _39506_ (
    .A(_05118_),
    .ZN(_05119_)
  );
  AND2_X1 _39507_ (
    .A1(_22078_),
    .A2(_05117_),
    .ZN(_05120_)
  );
  INV_X1 _39508_ (
    .A(_05120_),
    .ZN(_05121_)
  );
  AND2_X1 _39509_ (
    .A1(_05119_),
    .A2(_05121_),
    .ZN(_05122_)
  );
  AND2_X1 _39510_ (
    .A1(_22109_),
    .A2(_05122_),
    .ZN(_05123_)
  );
  INV_X1 _39511_ (
    .A(_05123_),
    .ZN(_05124_)
  );
  AND2_X1 _39512_ (
    .A1(_05087_),
    .A2(_05124_),
    .ZN(_05125_)
  );
  AND2_X1 _39513_ (
    .A1(_00007_[4]),
    .A2(_05049_),
    .ZN(_05126_)
  );
  INV_X1 _39514_ (
    .A(_05126_),
    .ZN(_05127_)
  );
  AND2_X1 _39515_ (
    .A1(_22144_),
    .A2(_05125_),
    .ZN(_05128_)
  );
  INV_X1 _39516_ (
    .A(_05128_),
    .ZN(_05129_)
  );
  AND2_X1 _39517_ (
    .A1(_04974_),
    .A2(_05129_),
    .ZN(_05130_)
  );
  AND2_X1 _39518_ (
    .A1(_05127_),
    .A2(_05130_),
    .ZN(_05131_)
  );
  AND2_X1 _39519_ (
    .A1(_04958_),
    .A2(_05131_),
    .ZN(_05132_)
  );
  INV_X1 _39520_ (
    .A(_05132_),
    .ZN(_05133_)
  );
  AND2_X1 _39521_ (
    .A1(_21288_),
    .A2(_21289_),
    .ZN(_05134_)
  );
  AND2_X1 _39522_ (
    .A1(_21293_),
    .A2(_05134_),
    .ZN(_05135_)
  );
  AND2_X1 _39523_ (
    .A1(_22271_),
    .A2(_05135_),
    .ZN(_05136_)
  );
  AND2_X1 _39524_ (
    .A1(_22540_),
    .A2(_05136_),
    .ZN(_05137_)
  );
  INV_X1 _39525_ (
    .A(_05137_),
    .ZN(_05138_)
  );
  AND2_X1 _39526_ (
    .A1(_05131_),
    .A2(_05137_),
    .ZN(_05139_)
  );
  INV_X1 _39527_ (
    .A(_05139_),
    .ZN(_05140_)
  );
  AND2_X1 _39528_ (
    .A1(_05133_),
    .A2(_05140_),
    .ZN(_05141_)
  );
  AND2_X1 _39529_ (
    .A1(_04969_),
    .A2(_05141_),
    .ZN(_05142_)
  );
  INV_X1 _39530_ (
    .A(_05142_),
    .ZN(_05143_)
  );
  AND2_X1 _39531_ (
    .A1(_04962_),
    .A2(_05143_),
    .ZN(_05144_)
  );
  INV_X1 _39532_ (
    .A(_05144_),
    .ZN(_05145_)
  );
  AND2_X1 _39533_ (
    .A1(reg_op2[0]),
    .A2(_04963_),
    .ZN(_05146_)
  );
  INV_X1 _39534_ (
    .A(_05146_),
    .ZN(_05147_)
  );
  AND2_X1 _39535_ (
    .A1(_05145_),
    .A2(_05147_),
    .ZN(_05148_)
  );
  INV_X1 _39536_ (
    .A(_05148_),
    .ZN(_00281_)
  );
  AND2_X1 _39537_ (
    .A1(decoded_imm[1]),
    .A2(_04966_),
    .ZN(_05149_)
  );
  INV_X1 _39538_ (
    .A(_05149_),
    .ZN(_05150_)
  );
  AND2_X1 _39539_ (
    .A1(_21437_),
    .A2(_22077_),
    .ZN(_05151_)
  );
  INV_X1 _39540_ (
    .A(_05151_),
    .ZN(_05152_)
  );
  AND2_X1 _39541_ (
    .A1(_21648_),
    .A2(_00007_[2]),
    .ZN(_05153_)
  );
  INV_X1 _39542_ (
    .A(_05153_),
    .ZN(_05154_)
  );
  AND2_X1 _39543_ (
    .A1(_05152_),
    .A2(_05154_),
    .ZN(_05155_)
  );
  AND2_X1 _39544_ (
    .A1(_21591_),
    .A2(_22077_),
    .ZN(_05156_)
  );
  INV_X1 _39545_ (
    .A(_05156_),
    .ZN(_05157_)
  );
  AND2_X1 _39546_ (
    .A1(_21409_),
    .A2(_00007_[2]),
    .ZN(_05158_)
  );
  INV_X1 _39547_ (
    .A(_05158_),
    .ZN(_05159_)
  );
  AND2_X1 _39548_ (
    .A1(_21459_),
    .A2(_22077_),
    .ZN(_05160_)
  );
  INV_X1 _39549_ (
    .A(_05160_),
    .ZN(_05161_)
  );
  AND2_X1 _39550_ (
    .A1(_21758_),
    .A2(_00007_[2]),
    .ZN(_05162_)
  );
  INV_X1 _39551_ (
    .A(_05162_),
    .ZN(_05163_)
  );
  AND2_X1 _39552_ (
    .A1(_21371_),
    .A2(_00007_[2]),
    .ZN(_05164_)
  );
  INV_X1 _39553_ (
    .A(_05164_),
    .ZN(_05165_)
  );
  AND2_X1 _39554_ (
    .A1(_21617_),
    .A2(_22077_),
    .ZN(_05166_)
  );
  INV_X1 _39555_ (
    .A(_05166_),
    .ZN(_05167_)
  );
  AND2_X1 _39556_ (
    .A1(_00007_[0]),
    .A2(_05167_),
    .ZN(_05168_)
  );
  AND2_X1 _39557_ (
    .A1(_05165_),
    .A2(_05168_),
    .ZN(_05169_)
  );
  INV_X1 _39558_ (
    .A(_05169_),
    .ZN(_05170_)
  );
  AND2_X1 _39559_ (
    .A1(_22152_),
    .A2(_05157_),
    .ZN(_05171_)
  );
  AND2_X1 _39560_ (
    .A1(_05159_),
    .A2(_05171_),
    .ZN(_05172_)
  );
  INV_X1 _39561_ (
    .A(_05172_),
    .ZN(_05173_)
  );
  AND2_X1 _39562_ (
    .A1(_05170_),
    .A2(_05173_),
    .ZN(_05174_)
  );
  AND2_X1 _39563_ (
    .A1(_00007_[1]),
    .A2(_05174_),
    .ZN(_05175_)
  );
  INV_X1 _39564_ (
    .A(_05175_),
    .ZN(_05176_)
  );
  AND2_X1 _39565_ (
    .A1(_00007_[0]),
    .A2(_05161_),
    .ZN(_05177_)
  );
  AND2_X1 _39566_ (
    .A1(_05163_),
    .A2(_05177_),
    .ZN(_05178_)
  );
  INV_X1 _39567_ (
    .A(_05178_),
    .ZN(_05179_)
  );
  AND2_X1 _39568_ (
    .A1(_22152_),
    .A2(_05155_),
    .ZN(_05180_)
  );
  INV_X1 _39569_ (
    .A(_05180_),
    .ZN(_05181_)
  );
  AND2_X1 _39570_ (
    .A1(_05179_),
    .A2(_05181_),
    .ZN(_05182_)
  );
  AND2_X1 _39571_ (
    .A1(_22078_),
    .A2(_05182_),
    .ZN(_05183_)
  );
  INV_X1 _39572_ (
    .A(_05183_),
    .ZN(_05184_)
  );
  AND2_X1 _39573_ (
    .A1(_05176_),
    .A2(_05184_),
    .ZN(_05185_)
  );
  AND2_X1 _39574_ (
    .A1(_22109_),
    .A2(_05185_),
    .ZN(_05186_)
  );
  INV_X1 _39575_ (
    .A(_05186_),
    .ZN(_05187_)
  );
  AND2_X1 _39576_ (
    .A1(_21890_),
    .A2(_00007_[2]),
    .ZN(_05188_)
  );
  INV_X1 _39577_ (
    .A(_05188_),
    .ZN(_05189_)
  );
  AND2_X1 _39578_ (
    .A1(_21834_),
    .A2(_22077_),
    .ZN(_05190_)
  );
  INV_X1 _39579_ (
    .A(_05190_),
    .ZN(_05191_)
  );
  AND2_X1 _39580_ (
    .A1(_00007_[0]),
    .A2(_05191_),
    .ZN(_05192_)
  );
  AND2_X1 _39581_ (
    .A1(_05189_),
    .A2(_05192_),
    .ZN(_05193_)
  );
  INV_X1 _39582_ (
    .A(_05193_),
    .ZN(_05194_)
  );
  AND2_X1 _39583_ (
    .A1(_21568_),
    .A2(_22077_),
    .ZN(_05195_)
  );
  INV_X1 _39584_ (
    .A(_05195_),
    .ZN(_05196_)
  );
  AND2_X1 _39585_ (
    .A1(_21906_),
    .A2(_00007_[2]),
    .ZN(_05197_)
  );
  INV_X1 _39586_ (
    .A(_05197_),
    .ZN(_05198_)
  );
  AND2_X1 _39587_ (
    .A1(_05196_),
    .A2(_05198_),
    .ZN(_05199_)
  );
  AND2_X1 _39588_ (
    .A1(_22152_),
    .A2(_05199_),
    .ZN(_05200_)
  );
  INV_X1 _39589_ (
    .A(_05200_),
    .ZN(_05201_)
  );
  AND2_X1 _39590_ (
    .A1(_05194_),
    .A2(_05201_),
    .ZN(_05202_)
  );
  AND2_X1 _39591_ (
    .A1(_22078_),
    .A2(_05202_),
    .ZN(_05203_)
  );
  INV_X1 _39592_ (
    .A(_05203_),
    .ZN(_05204_)
  );
  AND2_X1 _39593_ (
    .A1(_21866_),
    .A2(_22077_),
    .ZN(_05205_)
  );
  INV_X1 _39594_ (
    .A(_05205_),
    .ZN(_05206_)
  );
  AND2_X1 _39595_ (
    .A1(_21850_),
    .A2(_00007_[2]),
    .ZN(_05207_)
  );
  INV_X1 _39596_ (
    .A(_05207_),
    .ZN(_05208_)
  );
  AND2_X1 _39597_ (
    .A1(_05206_),
    .A2(_05208_),
    .ZN(_05209_)
  );
  AND2_X1 _39598_ (
    .A1(_22152_),
    .A2(_05209_),
    .ZN(_05210_)
  );
  INV_X1 _39599_ (
    .A(_05210_),
    .ZN(_05211_)
  );
  AND2_X1 _39600_ (
    .A1(_21938_),
    .A2(_00007_[2]),
    .ZN(_05212_)
  );
  INV_X1 _39601_ (
    .A(_05212_),
    .ZN(_05213_)
  );
  AND2_X1 _39602_ (
    .A1(_21922_),
    .A2(_22077_),
    .ZN(_05214_)
  );
  INV_X1 _39603_ (
    .A(_05214_),
    .ZN(_05215_)
  );
  AND2_X1 _39604_ (
    .A1(_00007_[0]),
    .A2(_05215_),
    .ZN(_05216_)
  );
  AND2_X1 _39605_ (
    .A1(_05213_),
    .A2(_05216_),
    .ZN(_05217_)
  );
  INV_X1 _39606_ (
    .A(_05217_),
    .ZN(_05218_)
  );
  AND2_X1 _39607_ (
    .A1(_05211_),
    .A2(_05218_),
    .ZN(_05219_)
  );
  AND2_X1 _39608_ (
    .A1(_00007_[1]),
    .A2(_05219_),
    .ZN(_05220_)
  );
  INV_X1 _39609_ (
    .A(_05220_),
    .ZN(_05221_)
  );
  AND2_X1 _39610_ (
    .A1(_00007_[3]),
    .A2(_05204_),
    .ZN(_05222_)
  );
  AND2_X1 _39611_ (
    .A1(_05221_),
    .A2(_05222_),
    .ZN(_05223_)
  );
  INV_X1 _39612_ (
    .A(_05223_),
    .ZN(_05224_)
  );
  AND2_X1 _39613_ (
    .A1(_05187_),
    .A2(_05224_),
    .ZN(_05225_)
  );
  AND2_X1 _39614_ (
    .A1(\cpuregs[9] [1]),
    .A2(_22077_),
    .ZN(_05226_)
  );
  INV_X1 _39615_ (
    .A(_05226_),
    .ZN(_05227_)
  );
  AND2_X1 _39616_ (
    .A1(\cpuregs[13] [1]),
    .A2(_00007_[2]),
    .ZN(_05228_)
  );
  INV_X1 _39617_ (
    .A(_05228_),
    .ZN(_05229_)
  );
  AND2_X1 _39618_ (
    .A1(_00007_[0]),
    .A2(_05229_),
    .ZN(_05230_)
  );
  AND2_X1 _39619_ (
    .A1(_05227_),
    .A2(_05230_),
    .ZN(_05231_)
  );
  INV_X1 _39620_ (
    .A(_05231_),
    .ZN(_05232_)
  );
  AND2_X1 _39621_ (
    .A1(\cpuregs[8] [1]),
    .A2(_22077_),
    .ZN(_05233_)
  );
  INV_X1 _39622_ (
    .A(_05233_),
    .ZN(_05234_)
  );
  AND2_X1 _39623_ (
    .A1(\cpuregs[12] [1]),
    .A2(_00007_[2]),
    .ZN(_05235_)
  );
  INV_X1 _39624_ (
    .A(_05235_),
    .ZN(_05236_)
  );
  AND2_X1 _39625_ (
    .A1(_22152_),
    .A2(_05236_),
    .ZN(_05237_)
  );
  AND2_X1 _39626_ (
    .A1(_05234_),
    .A2(_05237_),
    .ZN(_05238_)
  );
  INV_X1 _39627_ (
    .A(_05238_),
    .ZN(_05239_)
  );
  AND2_X1 _39628_ (
    .A1(_22078_),
    .A2(_05239_),
    .ZN(_05240_)
  );
  AND2_X1 _39629_ (
    .A1(_05232_),
    .A2(_05240_),
    .ZN(_05241_)
  );
  INV_X1 _39630_ (
    .A(_05241_),
    .ZN(_05242_)
  );
  AND2_X1 _39631_ (
    .A1(\cpuregs[15] [1]),
    .A2(_00007_[2]),
    .ZN(_05243_)
  );
  INV_X1 _39632_ (
    .A(_05243_),
    .ZN(_05244_)
  );
  AND2_X1 _39633_ (
    .A1(\cpuregs[11] [1]),
    .A2(_22077_),
    .ZN(_05245_)
  );
  INV_X1 _39634_ (
    .A(_05245_),
    .ZN(_05246_)
  );
  AND2_X1 _39635_ (
    .A1(_00007_[0]),
    .A2(_05246_),
    .ZN(_05247_)
  );
  AND2_X1 _39636_ (
    .A1(_05244_),
    .A2(_05247_),
    .ZN(_05248_)
  );
  INV_X1 _39637_ (
    .A(_05248_),
    .ZN(_05249_)
  );
  AND2_X1 _39638_ (
    .A1(\cpuregs[14] [1]),
    .A2(_00007_[2]),
    .ZN(_05250_)
  );
  INV_X1 _39639_ (
    .A(_05250_),
    .ZN(_05251_)
  );
  AND2_X1 _39640_ (
    .A1(\cpuregs[10] [1]),
    .A2(_22077_),
    .ZN(_05252_)
  );
  INV_X1 _39641_ (
    .A(_05252_),
    .ZN(_05253_)
  );
  AND2_X1 _39642_ (
    .A1(_22152_),
    .A2(_05253_),
    .ZN(_05254_)
  );
  AND2_X1 _39643_ (
    .A1(_05251_),
    .A2(_05254_),
    .ZN(_05255_)
  );
  INV_X1 _39644_ (
    .A(_05255_),
    .ZN(_05256_)
  );
  AND2_X1 _39645_ (
    .A1(_00007_[1]),
    .A2(_05256_),
    .ZN(_05257_)
  );
  AND2_X1 _39646_ (
    .A1(_05249_),
    .A2(_05257_),
    .ZN(_05258_)
  );
  INV_X1 _39647_ (
    .A(_05258_),
    .ZN(_05259_)
  );
  AND2_X1 _39648_ (
    .A1(_05242_),
    .A2(_05259_),
    .ZN(_05260_)
  );
  INV_X1 _39649_ (
    .A(_05260_),
    .ZN(_05261_)
  );
  AND2_X1 _39650_ (
    .A1(_00007_[3]),
    .A2(_05261_),
    .ZN(_05262_)
  );
  INV_X1 _39651_ (
    .A(_05262_),
    .ZN(_05263_)
  );
  AND2_X1 _39652_ (
    .A1(_21780_),
    .A2(_00007_[2]),
    .ZN(_05264_)
  );
  INV_X1 _39653_ (
    .A(_05264_),
    .ZN(_05265_)
  );
  AND2_X1 _39654_ (
    .A1(_21488_),
    .A2(_22077_),
    .ZN(_05266_)
  );
  INV_X1 _39655_ (
    .A(_05266_),
    .ZN(_05267_)
  );
  AND2_X1 _39656_ (
    .A1(_00007_[0]),
    .A2(_05267_),
    .ZN(_05268_)
  );
  AND2_X1 _39657_ (
    .A1(_05265_),
    .A2(_05268_),
    .ZN(_05269_)
  );
  INV_X1 _39658_ (
    .A(_05269_),
    .ZN(_05270_)
  );
  AND2_X1 _39659_ (
    .A1(_21805_),
    .A2(_00007_[2]),
    .ZN(_05271_)
  );
  INV_X1 _39660_ (
    .A(_05271_),
    .ZN(_05272_)
  );
  AND2_X1 _39661_ (
    .A1(_21538_),
    .A2(_22077_),
    .ZN(_05273_)
  );
  INV_X1 _39662_ (
    .A(_05273_),
    .ZN(_05274_)
  );
  AND2_X1 _39663_ (
    .A1(_22152_),
    .A2(_05274_),
    .ZN(_05275_)
  );
  AND2_X1 _39664_ (
    .A1(_05272_),
    .A2(_05275_),
    .ZN(_05276_)
  );
  INV_X1 _39665_ (
    .A(_05276_),
    .ZN(_05277_)
  );
  AND2_X1 _39666_ (
    .A1(_05270_),
    .A2(_05277_),
    .ZN(_05278_)
  );
  AND2_X1 _39667_ (
    .A1(_00007_[1]),
    .A2(_05278_),
    .ZN(_05279_)
  );
  INV_X1 _39668_ (
    .A(_05279_),
    .ZN(_05280_)
  );
  AND2_X1 _39669_ (
    .A1(_21733_),
    .A2(_00007_[2]),
    .ZN(_05281_)
  );
  INV_X1 _39670_ (
    .A(_05281_),
    .ZN(_05282_)
  );
  AND2_X1 _39671_ (
    .A1(_21513_),
    .A2(_22077_),
    .ZN(_05283_)
  );
  INV_X1 _39672_ (
    .A(_05283_),
    .ZN(_05284_)
  );
  AND2_X1 _39673_ (
    .A1(_00007_[0]),
    .A2(_05284_),
    .ZN(_05285_)
  );
  AND2_X1 _39674_ (
    .A1(_05282_),
    .A2(_05285_),
    .ZN(_05286_)
  );
  INV_X1 _39675_ (
    .A(_05286_),
    .ZN(_05287_)
  );
  AND2_X1 _39676_ (
    .A1(_21954_),
    .A2(_22077_),
    .ZN(_05288_)
  );
  INV_X1 _39677_ (
    .A(_05288_),
    .ZN(_05289_)
  );
  AND2_X1 _39678_ (
    .A1(_21670_),
    .A2(_00007_[2]),
    .ZN(_05290_)
  );
  INV_X1 _39679_ (
    .A(_05290_),
    .ZN(_05291_)
  );
  AND2_X1 _39680_ (
    .A1(_05289_),
    .A2(_05291_),
    .ZN(_05292_)
  );
  AND2_X1 _39681_ (
    .A1(_22152_),
    .A2(_05292_),
    .ZN(_05293_)
  );
  INV_X1 _39682_ (
    .A(_05293_),
    .ZN(_05294_)
  );
  AND2_X1 _39683_ (
    .A1(_05287_),
    .A2(_05294_),
    .ZN(_05295_)
  );
  AND2_X1 _39684_ (
    .A1(_22078_),
    .A2(_05295_),
    .ZN(_05296_)
  );
  INV_X1 _39685_ (
    .A(_05296_),
    .ZN(_05297_)
  );
  AND2_X1 _39686_ (
    .A1(_05280_),
    .A2(_05297_),
    .ZN(_05298_)
  );
  AND2_X1 _39687_ (
    .A1(_22109_),
    .A2(_05298_),
    .ZN(_05299_)
  );
  INV_X1 _39688_ (
    .A(_05299_),
    .ZN(_05300_)
  );
  AND2_X1 _39689_ (
    .A1(_00007_[4]),
    .A2(_05225_),
    .ZN(_05301_)
  );
  INV_X1 _39690_ (
    .A(_05301_),
    .ZN(_05302_)
  );
  AND2_X1 _39691_ (
    .A1(_22144_),
    .A2(_05300_),
    .ZN(_05303_)
  );
  AND2_X1 _39692_ (
    .A1(_05263_),
    .A2(_05303_),
    .ZN(_05304_)
  );
  INV_X1 _39693_ (
    .A(_05304_),
    .ZN(_05305_)
  );
  AND2_X1 _39694_ (
    .A1(_04974_),
    .A2(_05305_),
    .ZN(_05306_)
  );
  AND2_X1 _39695_ (
    .A1(_05302_),
    .A2(_05306_),
    .ZN(_05307_)
  );
  AND2_X1 _39696_ (
    .A1(_04958_),
    .A2(_05307_),
    .ZN(_05308_)
  );
  INV_X1 _39697_ (
    .A(_05308_),
    .ZN(_05309_)
  );
  AND2_X1 _39698_ (
    .A1(_05137_),
    .A2(_05307_),
    .ZN(_05310_)
  );
  INV_X1 _39699_ (
    .A(_05310_),
    .ZN(_05311_)
  );
  AND2_X1 _39700_ (
    .A1(_05309_),
    .A2(_05311_),
    .ZN(_05312_)
  );
  AND2_X1 _39701_ (
    .A1(_05150_),
    .A2(_05312_),
    .ZN(_05313_)
  );
  INV_X1 _39702_ (
    .A(_05313_),
    .ZN(_05314_)
  );
  AND2_X1 _39703_ (
    .A1(_04962_),
    .A2(_05314_),
    .ZN(_05315_)
  );
  INV_X1 _39704_ (
    .A(_05315_),
    .ZN(_05316_)
  );
  AND2_X1 _39705_ (
    .A1(reg_op2[1]),
    .A2(_04963_),
    .ZN(_05317_)
  );
  INV_X1 _39706_ (
    .A(_05317_),
    .ZN(_05318_)
  );
  AND2_X1 _39707_ (
    .A1(_05316_),
    .A2(_05318_),
    .ZN(_05319_)
  );
  INV_X1 _39708_ (
    .A(_05319_),
    .ZN(_00282_)
  );
  AND2_X1 _39709_ (
    .A1(decoded_imm[2]),
    .A2(_04966_),
    .ZN(_05320_)
  );
  INV_X1 _39710_ (
    .A(_05320_),
    .ZN(_05321_)
  );
  AND2_X1 _39711_ (
    .A1(_21438_),
    .A2(_22077_),
    .ZN(_05322_)
  );
  INV_X1 _39712_ (
    .A(_05322_),
    .ZN(_05323_)
  );
  AND2_X1 _39713_ (
    .A1(_21649_),
    .A2(_00007_[2]),
    .ZN(_05324_)
  );
  INV_X1 _39714_ (
    .A(_05324_),
    .ZN(_05325_)
  );
  AND2_X1 _39715_ (
    .A1(_05323_),
    .A2(_05325_),
    .ZN(_05326_)
  );
  AND2_X1 _39716_ (
    .A1(_21592_),
    .A2(_22077_),
    .ZN(_05327_)
  );
  INV_X1 _39717_ (
    .A(_05327_),
    .ZN(_05328_)
  );
  AND2_X1 _39718_ (
    .A1(_21410_),
    .A2(_00007_[2]),
    .ZN(_05329_)
  );
  INV_X1 _39719_ (
    .A(_05329_),
    .ZN(_05330_)
  );
  AND2_X1 _39720_ (
    .A1(_21460_),
    .A2(_22077_),
    .ZN(_05331_)
  );
  INV_X1 _39721_ (
    .A(_05331_),
    .ZN(_05332_)
  );
  AND2_X1 _39722_ (
    .A1(_21759_),
    .A2(_00007_[2]),
    .ZN(_05333_)
  );
  INV_X1 _39723_ (
    .A(_05333_),
    .ZN(_05334_)
  );
  AND2_X1 _39724_ (
    .A1(_21372_),
    .A2(_00007_[2]),
    .ZN(_05335_)
  );
  INV_X1 _39725_ (
    .A(_05335_),
    .ZN(_05336_)
  );
  AND2_X1 _39726_ (
    .A1(_21618_),
    .A2(_22077_),
    .ZN(_05337_)
  );
  INV_X1 _39727_ (
    .A(_05337_),
    .ZN(_05338_)
  );
  AND2_X1 _39728_ (
    .A1(_00007_[0]),
    .A2(_05338_),
    .ZN(_05339_)
  );
  AND2_X1 _39729_ (
    .A1(_05336_),
    .A2(_05339_),
    .ZN(_05340_)
  );
  INV_X1 _39730_ (
    .A(_05340_),
    .ZN(_05341_)
  );
  AND2_X1 _39731_ (
    .A1(_22152_),
    .A2(_05328_),
    .ZN(_05342_)
  );
  AND2_X1 _39732_ (
    .A1(_05330_),
    .A2(_05342_),
    .ZN(_05343_)
  );
  INV_X1 _39733_ (
    .A(_05343_),
    .ZN(_05344_)
  );
  AND2_X1 _39734_ (
    .A1(_05341_),
    .A2(_05344_),
    .ZN(_05345_)
  );
  AND2_X1 _39735_ (
    .A1(_00007_[1]),
    .A2(_05345_),
    .ZN(_05346_)
  );
  INV_X1 _39736_ (
    .A(_05346_),
    .ZN(_05347_)
  );
  AND2_X1 _39737_ (
    .A1(_00007_[0]),
    .A2(_05332_),
    .ZN(_05348_)
  );
  AND2_X1 _39738_ (
    .A1(_05334_),
    .A2(_05348_),
    .ZN(_05349_)
  );
  INV_X1 _39739_ (
    .A(_05349_),
    .ZN(_05350_)
  );
  AND2_X1 _39740_ (
    .A1(_22152_),
    .A2(_05326_),
    .ZN(_05351_)
  );
  INV_X1 _39741_ (
    .A(_05351_),
    .ZN(_05352_)
  );
  AND2_X1 _39742_ (
    .A1(_05350_),
    .A2(_05352_),
    .ZN(_05353_)
  );
  AND2_X1 _39743_ (
    .A1(_22078_),
    .A2(_05353_),
    .ZN(_05354_)
  );
  INV_X1 _39744_ (
    .A(_05354_),
    .ZN(_05355_)
  );
  AND2_X1 _39745_ (
    .A1(_05347_),
    .A2(_05355_),
    .ZN(_05356_)
  );
  AND2_X1 _39746_ (
    .A1(_22109_),
    .A2(_05356_),
    .ZN(_05357_)
  );
  INV_X1 _39747_ (
    .A(_05357_),
    .ZN(_05358_)
  );
  AND2_X1 _39748_ (
    .A1(_21891_),
    .A2(_00007_[2]),
    .ZN(_05359_)
  );
  INV_X1 _39749_ (
    .A(_05359_),
    .ZN(_05360_)
  );
  AND2_X1 _39750_ (
    .A1(_21835_),
    .A2(_22077_),
    .ZN(_05361_)
  );
  INV_X1 _39751_ (
    .A(_05361_),
    .ZN(_05362_)
  );
  AND2_X1 _39752_ (
    .A1(_00007_[0]),
    .A2(_05362_),
    .ZN(_05363_)
  );
  AND2_X1 _39753_ (
    .A1(_05360_),
    .A2(_05363_),
    .ZN(_05364_)
  );
  INV_X1 _39754_ (
    .A(_05364_),
    .ZN(_05365_)
  );
  AND2_X1 _39755_ (
    .A1(_21569_),
    .A2(_22077_),
    .ZN(_05366_)
  );
  INV_X1 _39756_ (
    .A(_05366_),
    .ZN(_05367_)
  );
  AND2_X1 _39757_ (
    .A1(_21907_),
    .A2(_00007_[2]),
    .ZN(_05368_)
  );
  INV_X1 _39758_ (
    .A(_05368_),
    .ZN(_05369_)
  );
  AND2_X1 _39759_ (
    .A1(_05367_),
    .A2(_05369_),
    .ZN(_05370_)
  );
  AND2_X1 _39760_ (
    .A1(_22152_),
    .A2(_05370_),
    .ZN(_05371_)
  );
  INV_X1 _39761_ (
    .A(_05371_),
    .ZN(_05372_)
  );
  AND2_X1 _39762_ (
    .A1(_05365_),
    .A2(_05372_),
    .ZN(_05373_)
  );
  AND2_X1 _39763_ (
    .A1(_22078_),
    .A2(_05373_),
    .ZN(_05374_)
  );
  INV_X1 _39764_ (
    .A(_05374_),
    .ZN(_05375_)
  );
  AND2_X1 _39765_ (
    .A1(_21867_),
    .A2(_22077_),
    .ZN(_05376_)
  );
  INV_X1 _39766_ (
    .A(_05376_),
    .ZN(_05377_)
  );
  AND2_X1 _39767_ (
    .A1(_21851_),
    .A2(_00007_[2]),
    .ZN(_05378_)
  );
  INV_X1 _39768_ (
    .A(_05378_),
    .ZN(_05379_)
  );
  AND2_X1 _39769_ (
    .A1(_05377_),
    .A2(_05379_),
    .ZN(_05380_)
  );
  AND2_X1 _39770_ (
    .A1(_22152_),
    .A2(_05380_),
    .ZN(_05381_)
  );
  INV_X1 _39771_ (
    .A(_05381_),
    .ZN(_05382_)
  );
  AND2_X1 _39772_ (
    .A1(_21939_),
    .A2(_00007_[2]),
    .ZN(_05383_)
  );
  INV_X1 _39773_ (
    .A(_05383_),
    .ZN(_05384_)
  );
  AND2_X1 _39774_ (
    .A1(_21923_),
    .A2(_22077_),
    .ZN(_05385_)
  );
  INV_X1 _39775_ (
    .A(_05385_),
    .ZN(_05386_)
  );
  AND2_X1 _39776_ (
    .A1(_00007_[0]),
    .A2(_05386_),
    .ZN(_05387_)
  );
  AND2_X1 _39777_ (
    .A1(_05384_),
    .A2(_05387_),
    .ZN(_05388_)
  );
  INV_X1 _39778_ (
    .A(_05388_),
    .ZN(_05389_)
  );
  AND2_X1 _39779_ (
    .A1(_05382_),
    .A2(_05389_),
    .ZN(_05390_)
  );
  AND2_X1 _39780_ (
    .A1(_00007_[1]),
    .A2(_05390_),
    .ZN(_05391_)
  );
  INV_X1 _39781_ (
    .A(_05391_),
    .ZN(_05392_)
  );
  AND2_X1 _39782_ (
    .A1(_00007_[3]),
    .A2(_05375_),
    .ZN(_05393_)
  );
  AND2_X1 _39783_ (
    .A1(_05392_),
    .A2(_05393_),
    .ZN(_05394_)
  );
  INV_X1 _39784_ (
    .A(_05394_),
    .ZN(_05395_)
  );
  AND2_X1 _39785_ (
    .A1(_05358_),
    .A2(_05395_),
    .ZN(_05396_)
  );
  AND2_X1 _39786_ (
    .A1(\cpuregs[9] [2]),
    .A2(_22077_),
    .ZN(_05397_)
  );
  INV_X1 _39787_ (
    .A(_05397_),
    .ZN(_05398_)
  );
  AND2_X1 _39788_ (
    .A1(\cpuregs[13] [2]),
    .A2(_00007_[2]),
    .ZN(_05399_)
  );
  INV_X1 _39789_ (
    .A(_05399_),
    .ZN(_05400_)
  );
  AND2_X1 _39790_ (
    .A1(_00007_[0]),
    .A2(_05400_),
    .ZN(_05401_)
  );
  AND2_X1 _39791_ (
    .A1(_05398_),
    .A2(_05401_),
    .ZN(_05402_)
  );
  INV_X1 _39792_ (
    .A(_05402_),
    .ZN(_05403_)
  );
  AND2_X1 _39793_ (
    .A1(\cpuregs[8] [2]),
    .A2(_22077_),
    .ZN(_05404_)
  );
  INV_X1 _39794_ (
    .A(_05404_),
    .ZN(_05405_)
  );
  AND2_X1 _39795_ (
    .A1(\cpuregs[12] [2]),
    .A2(_00007_[2]),
    .ZN(_05406_)
  );
  INV_X1 _39796_ (
    .A(_05406_),
    .ZN(_05407_)
  );
  AND2_X1 _39797_ (
    .A1(_22152_),
    .A2(_05407_),
    .ZN(_05408_)
  );
  AND2_X1 _39798_ (
    .A1(_05405_),
    .A2(_05408_),
    .ZN(_05409_)
  );
  INV_X1 _39799_ (
    .A(_05409_),
    .ZN(_05410_)
  );
  AND2_X1 _39800_ (
    .A1(_22078_),
    .A2(_05410_),
    .ZN(_05411_)
  );
  AND2_X1 _39801_ (
    .A1(_05403_),
    .A2(_05411_),
    .ZN(_05412_)
  );
  INV_X1 _39802_ (
    .A(_05412_),
    .ZN(_05413_)
  );
  AND2_X1 _39803_ (
    .A1(\cpuregs[15] [2]),
    .A2(_00007_[2]),
    .ZN(_05414_)
  );
  INV_X1 _39804_ (
    .A(_05414_),
    .ZN(_05415_)
  );
  AND2_X1 _39805_ (
    .A1(\cpuregs[11] [2]),
    .A2(_22077_),
    .ZN(_05416_)
  );
  INV_X1 _39806_ (
    .A(_05416_),
    .ZN(_05417_)
  );
  AND2_X1 _39807_ (
    .A1(_00007_[0]),
    .A2(_05417_),
    .ZN(_05418_)
  );
  AND2_X1 _39808_ (
    .A1(_05415_),
    .A2(_05418_),
    .ZN(_05419_)
  );
  INV_X1 _39809_ (
    .A(_05419_),
    .ZN(_05420_)
  );
  AND2_X1 _39810_ (
    .A1(\cpuregs[14] [2]),
    .A2(_00007_[2]),
    .ZN(_05421_)
  );
  INV_X1 _39811_ (
    .A(_05421_),
    .ZN(_05422_)
  );
  AND2_X1 _39812_ (
    .A1(\cpuregs[10] [2]),
    .A2(_22077_),
    .ZN(_05423_)
  );
  INV_X1 _39813_ (
    .A(_05423_),
    .ZN(_05424_)
  );
  AND2_X1 _39814_ (
    .A1(_22152_),
    .A2(_05424_),
    .ZN(_05425_)
  );
  AND2_X1 _39815_ (
    .A1(_05422_),
    .A2(_05425_),
    .ZN(_05426_)
  );
  INV_X1 _39816_ (
    .A(_05426_),
    .ZN(_05427_)
  );
  AND2_X1 _39817_ (
    .A1(_00007_[1]),
    .A2(_05427_),
    .ZN(_05428_)
  );
  AND2_X1 _39818_ (
    .A1(_05420_),
    .A2(_05428_),
    .ZN(_05429_)
  );
  INV_X1 _39819_ (
    .A(_05429_),
    .ZN(_05430_)
  );
  AND2_X1 _39820_ (
    .A1(_05413_),
    .A2(_05430_),
    .ZN(_05431_)
  );
  INV_X1 _39821_ (
    .A(_05431_),
    .ZN(_05432_)
  );
  AND2_X1 _39822_ (
    .A1(_00007_[3]),
    .A2(_05432_),
    .ZN(_05433_)
  );
  INV_X1 _39823_ (
    .A(_05433_),
    .ZN(_05434_)
  );
  AND2_X1 _39824_ (
    .A1(_21781_),
    .A2(_00007_[2]),
    .ZN(_05435_)
  );
  INV_X1 _39825_ (
    .A(_05435_),
    .ZN(_05436_)
  );
  AND2_X1 _39826_ (
    .A1(_21489_),
    .A2(_22077_),
    .ZN(_05437_)
  );
  INV_X1 _39827_ (
    .A(_05437_),
    .ZN(_05438_)
  );
  AND2_X1 _39828_ (
    .A1(_00007_[0]),
    .A2(_05438_),
    .ZN(_05439_)
  );
  AND2_X1 _39829_ (
    .A1(_05436_),
    .A2(_05439_),
    .ZN(_05440_)
  );
  INV_X1 _39830_ (
    .A(_05440_),
    .ZN(_05441_)
  );
  AND2_X1 _39831_ (
    .A1(_21806_),
    .A2(_00007_[2]),
    .ZN(_05442_)
  );
  INV_X1 _39832_ (
    .A(_05442_),
    .ZN(_05443_)
  );
  AND2_X1 _39833_ (
    .A1(_21539_),
    .A2(_22077_),
    .ZN(_05444_)
  );
  INV_X1 _39834_ (
    .A(_05444_),
    .ZN(_05445_)
  );
  AND2_X1 _39835_ (
    .A1(_22152_),
    .A2(_05445_),
    .ZN(_05446_)
  );
  AND2_X1 _39836_ (
    .A1(_05443_),
    .A2(_05446_),
    .ZN(_05447_)
  );
  INV_X1 _39837_ (
    .A(_05447_),
    .ZN(_05448_)
  );
  AND2_X1 _39838_ (
    .A1(_05441_),
    .A2(_05448_),
    .ZN(_05449_)
  );
  AND2_X1 _39839_ (
    .A1(_00007_[1]),
    .A2(_05449_),
    .ZN(_05450_)
  );
  INV_X1 _39840_ (
    .A(_05450_),
    .ZN(_05451_)
  );
  AND2_X1 _39841_ (
    .A1(_21734_),
    .A2(_00007_[2]),
    .ZN(_05452_)
  );
  INV_X1 _39842_ (
    .A(_05452_),
    .ZN(_05453_)
  );
  AND2_X1 _39843_ (
    .A1(_21514_),
    .A2(_22077_),
    .ZN(_05454_)
  );
  INV_X1 _39844_ (
    .A(_05454_),
    .ZN(_05455_)
  );
  AND2_X1 _39845_ (
    .A1(_00007_[0]),
    .A2(_05455_),
    .ZN(_05456_)
  );
  AND2_X1 _39846_ (
    .A1(_05453_),
    .A2(_05456_),
    .ZN(_05457_)
  );
  INV_X1 _39847_ (
    .A(_05457_),
    .ZN(_05458_)
  );
  AND2_X1 _39848_ (
    .A1(_21955_),
    .A2(_22077_),
    .ZN(_05459_)
  );
  INV_X1 _39849_ (
    .A(_05459_),
    .ZN(_05460_)
  );
  AND2_X1 _39850_ (
    .A1(_21671_),
    .A2(_00007_[2]),
    .ZN(_05461_)
  );
  INV_X1 _39851_ (
    .A(_05461_),
    .ZN(_05462_)
  );
  AND2_X1 _39852_ (
    .A1(_05460_),
    .A2(_05462_),
    .ZN(_05463_)
  );
  AND2_X1 _39853_ (
    .A1(_22152_),
    .A2(_05463_),
    .ZN(_05464_)
  );
  INV_X1 _39854_ (
    .A(_05464_),
    .ZN(_05465_)
  );
  AND2_X1 _39855_ (
    .A1(_05458_),
    .A2(_05465_),
    .ZN(_05466_)
  );
  AND2_X1 _39856_ (
    .A1(_22078_),
    .A2(_05466_),
    .ZN(_05467_)
  );
  INV_X1 _39857_ (
    .A(_05467_),
    .ZN(_05468_)
  );
  AND2_X1 _39858_ (
    .A1(_05451_),
    .A2(_05468_),
    .ZN(_05469_)
  );
  AND2_X1 _39859_ (
    .A1(_22109_),
    .A2(_05469_),
    .ZN(_05470_)
  );
  INV_X1 _39860_ (
    .A(_05470_),
    .ZN(_05471_)
  );
  AND2_X1 _39861_ (
    .A1(_00007_[4]),
    .A2(_05396_),
    .ZN(_05472_)
  );
  INV_X1 _39862_ (
    .A(_05472_),
    .ZN(_05473_)
  );
  AND2_X1 _39863_ (
    .A1(_22144_),
    .A2(_05471_),
    .ZN(_05474_)
  );
  AND2_X1 _39864_ (
    .A1(_05434_),
    .A2(_05474_),
    .ZN(_05475_)
  );
  INV_X1 _39865_ (
    .A(_05475_),
    .ZN(_05476_)
  );
  AND2_X1 _39866_ (
    .A1(_04974_),
    .A2(_05476_),
    .ZN(_05477_)
  );
  AND2_X1 _39867_ (
    .A1(_05473_),
    .A2(_05477_),
    .ZN(_05478_)
  );
  AND2_X1 _39868_ (
    .A1(_04958_),
    .A2(_05478_),
    .ZN(_05479_)
  );
  INV_X1 _39869_ (
    .A(_05479_),
    .ZN(_05480_)
  );
  AND2_X1 _39870_ (
    .A1(_05137_),
    .A2(_05478_),
    .ZN(_05481_)
  );
  INV_X1 _39871_ (
    .A(_05481_),
    .ZN(_05482_)
  );
  AND2_X1 _39872_ (
    .A1(_05480_),
    .A2(_05482_),
    .ZN(_05483_)
  );
  AND2_X1 _39873_ (
    .A1(_05321_),
    .A2(_05483_),
    .ZN(_05484_)
  );
  AND2_X1 _39874_ (
    .A1(_21202_),
    .A2(_04963_),
    .ZN(_05485_)
  );
  INV_X1 _39875_ (
    .A(_05485_),
    .ZN(_05486_)
  );
  AND2_X1 _39876_ (
    .A1(_04962_),
    .A2(_05484_),
    .ZN(_05487_)
  );
  INV_X1 _39877_ (
    .A(_05487_),
    .ZN(_05488_)
  );
  AND2_X1 _39878_ (
    .A1(_05486_),
    .A2(_05488_),
    .ZN(_00283_)
  );
  AND2_X1 _39879_ (
    .A1(decoded_imm[3]),
    .A2(_04966_),
    .ZN(_05489_)
  );
  INV_X1 _39880_ (
    .A(_05489_),
    .ZN(_05490_)
  );
  AND2_X1 _39881_ (
    .A1(\cpuregs[31] [3]),
    .A2(_00007_[1]),
    .ZN(_05491_)
  );
  INV_X1 _39882_ (
    .A(_05491_),
    .ZN(_05492_)
  );
  AND2_X1 _39883_ (
    .A1(\cpuregs[29] [3]),
    .A2(_22078_),
    .ZN(_05493_)
  );
  INV_X1 _39884_ (
    .A(_05493_),
    .ZN(_05494_)
  );
  AND2_X1 _39885_ (
    .A1(_05492_),
    .A2(_05494_),
    .ZN(_05495_)
  );
  INV_X1 _39886_ (
    .A(_05495_),
    .ZN(_05496_)
  );
  AND2_X1 _39887_ (
    .A1(_00007_[2]),
    .A2(_05496_),
    .ZN(_05497_)
  );
  INV_X1 _39888_ (
    .A(_05497_),
    .ZN(_05498_)
  );
  AND2_X1 _39889_ (
    .A1(\cpuregs[27] [3]),
    .A2(_00007_[1]),
    .ZN(_05499_)
  );
  INV_X1 _39890_ (
    .A(_05499_),
    .ZN(_05500_)
  );
  AND2_X1 _39891_ (
    .A1(\cpuregs[25] [3]),
    .A2(_22078_),
    .ZN(_05501_)
  );
  INV_X1 _39892_ (
    .A(_05501_),
    .ZN(_05502_)
  );
  AND2_X1 _39893_ (
    .A1(_05500_),
    .A2(_05502_),
    .ZN(_05503_)
  );
  INV_X1 _39894_ (
    .A(_05503_),
    .ZN(_05504_)
  );
  AND2_X1 _39895_ (
    .A1(_22077_),
    .A2(_05504_),
    .ZN(_05505_)
  );
  INV_X1 _39896_ (
    .A(_05505_),
    .ZN(_05506_)
  );
  AND2_X1 _39897_ (
    .A1(_05498_),
    .A2(_05506_),
    .ZN(_05507_)
  );
  INV_X1 _39898_ (
    .A(_05507_),
    .ZN(_05508_)
  );
  AND2_X1 _39899_ (
    .A1(_00007_[0]),
    .A2(_05508_),
    .ZN(_05509_)
  );
  INV_X1 _39900_ (
    .A(_05509_),
    .ZN(_05510_)
  );
  AND2_X1 _39901_ (
    .A1(\cpuregs[30] [3]),
    .A2(_00007_[1]),
    .ZN(_05511_)
  );
  INV_X1 _39902_ (
    .A(_05511_),
    .ZN(_05512_)
  );
  AND2_X1 _39903_ (
    .A1(\cpuregs[28] [3]),
    .A2(_22078_),
    .ZN(_05513_)
  );
  INV_X1 _39904_ (
    .A(_05513_),
    .ZN(_05514_)
  );
  AND2_X1 _39905_ (
    .A1(_05512_),
    .A2(_05514_),
    .ZN(_05515_)
  );
  INV_X1 _39906_ (
    .A(_05515_),
    .ZN(_05516_)
  );
  AND2_X1 _39907_ (
    .A1(_00007_[2]),
    .A2(_05516_),
    .ZN(_05517_)
  );
  INV_X1 _39908_ (
    .A(_05517_),
    .ZN(_05518_)
  );
  AND2_X1 _39909_ (
    .A1(\cpuregs[26] [3]),
    .A2(_00007_[1]),
    .ZN(_05519_)
  );
  INV_X1 _39910_ (
    .A(_05519_),
    .ZN(_05520_)
  );
  AND2_X1 _39911_ (
    .A1(\cpuregs[24] [3]),
    .A2(_22078_),
    .ZN(_05521_)
  );
  INV_X1 _39912_ (
    .A(_05521_),
    .ZN(_05522_)
  );
  AND2_X1 _39913_ (
    .A1(_05520_),
    .A2(_05522_),
    .ZN(_05523_)
  );
  INV_X1 _39914_ (
    .A(_05523_),
    .ZN(_05524_)
  );
  AND2_X1 _39915_ (
    .A1(_22077_),
    .A2(_05524_),
    .ZN(_05525_)
  );
  INV_X1 _39916_ (
    .A(_05525_),
    .ZN(_05526_)
  );
  AND2_X1 _39917_ (
    .A1(_05518_),
    .A2(_05526_),
    .ZN(_05527_)
  );
  INV_X1 _39918_ (
    .A(_05527_),
    .ZN(_05528_)
  );
  AND2_X1 _39919_ (
    .A1(_22152_),
    .A2(_05528_),
    .ZN(_05529_)
  );
  INV_X1 _39920_ (
    .A(_05529_),
    .ZN(_05530_)
  );
  AND2_X1 _39921_ (
    .A1(_05510_),
    .A2(_05530_),
    .ZN(_05531_)
  );
  INV_X1 _39922_ (
    .A(_05531_),
    .ZN(_05532_)
  );
  AND2_X1 _39923_ (
    .A1(_00007_[3]),
    .A2(_05532_),
    .ZN(_05533_)
  );
  INV_X1 _39924_ (
    .A(_05533_),
    .ZN(_05534_)
  );
  AND2_X1 _39925_ (
    .A1(_21593_),
    .A2(_22077_),
    .ZN(_05535_)
  );
  INV_X1 _39926_ (
    .A(_05535_),
    .ZN(_05536_)
  );
  AND2_X1 _39927_ (
    .A1(_21411_),
    .A2(_00007_[2]),
    .ZN(_05537_)
  );
  INV_X1 _39928_ (
    .A(_05537_),
    .ZN(_05538_)
  );
  AND2_X1 _39929_ (
    .A1(_21439_),
    .A2(_22077_),
    .ZN(_05539_)
  );
  INV_X1 _39930_ (
    .A(_05539_),
    .ZN(_05540_)
  );
  AND2_X1 _39931_ (
    .A1(_21650_),
    .A2(_00007_[2]),
    .ZN(_05541_)
  );
  INV_X1 _39932_ (
    .A(_05541_),
    .ZN(_05542_)
  );
  AND2_X1 _39933_ (
    .A1(_05540_),
    .A2(_05542_),
    .ZN(_05543_)
  );
  AND2_X1 _39934_ (
    .A1(_21373_),
    .A2(_00007_[2]),
    .ZN(_05544_)
  );
  INV_X1 _39935_ (
    .A(_05544_),
    .ZN(_05545_)
  );
  AND2_X1 _39936_ (
    .A1(_21619_),
    .A2(_22077_),
    .ZN(_05546_)
  );
  INV_X1 _39937_ (
    .A(_05546_),
    .ZN(_05547_)
  );
  AND2_X1 _39938_ (
    .A1(_21461_),
    .A2(_22077_),
    .ZN(_05548_)
  );
  INV_X1 _39939_ (
    .A(_05548_),
    .ZN(_05549_)
  );
  AND2_X1 _39940_ (
    .A1(_21760_),
    .A2(_00007_[2]),
    .ZN(_05550_)
  );
  INV_X1 _39941_ (
    .A(_05550_),
    .ZN(_05551_)
  );
  AND2_X1 _39942_ (
    .A1(_00007_[0]),
    .A2(_05547_),
    .ZN(_05552_)
  );
  AND2_X1 _39943_ (
    .A1(_05545_),
    .A2(_05552_),
    .ZN(_05553_)
  );
  INV_X1 _39944_ (
    .A(_05553_),
    .ZN(_05554_)
  );
  AND2_X1 _39945_ (
    .A1(_22152_),
    .A2(_05536_),
    .ZN(_05555_)
  );
  AND2_X1 _39946_ (
    .A1(_05538_),
    .A2(_05555_),
    .ZN(_05556_)
  );
  INV_X1 _39947_ (
    .A(_05556_),
    .ZN(_05557_)
  );
  AND2_X1 _39948_ (
    .A1(_05554_),
    .A2(_05557_),
    .ZN(_05558_)
  );
  AND2_X1 _39949_ (
    .A1(_00007_[1]),
    .A2(_05558_),
    .ZN(_05559_)
  );
  INV_X1 _39950_ (
    .A(_05559_),
    .ZN(_05560_)
  );
  AND2_X1 _39951_ (
    .A1(_00007_[0]),
    .A2(_05549_),
    .ZN(_05561_)
  );
  AND2_X1 _39952_ (
    .A1(_05551_),
    .A2(_05561_),
    .ZN(_05562_)
  );
  INV_X1 _39953_ (
    .A(_05562_),
    .ZN(_05563_)
  );
  AND2_X1 _39954_ (
    .A1(_22152_),
    .A2(_05543_),
    .ZN(_05564_)
  );
  INV_X1 _39955_ (
    .A(_05564_),
    .ZN(_05565_)
  );
  AND2_X1 _39956_ (
    .A1(_05563_),
    .A2(_05565_),
    .ZN(_05566_)
  );
  AND2_X1 _39957_ (
    .A1(_22078_),
    .A2(_05566_),
    .ZN(_05567_)
  );
  INV_X1 _39958_ (
    .A(_05567_),
    .ZN(_05568_)
  );
  AND2_X1 _39959_ (
    .A1(_05560_),
    .A2(_05568_),
    .ZN(_05569_)
  );
  AND2_X1 _39960_ (
    .A1(_22109_),
    .A2(_05569_),
    .ZN(_05570_)
  );
  INV_X1 _39961_ (
    .A(_05570_),
    .ZN(_05571_)
  );
  AND2_X1 _39962_ (
    .A1(_05534_),
    .A2(_05571_),
    .ZN(_05572_)
  );
  AND2_X1 _39963_ (
    .A1(\cpuregs[13] [3]),
    .A2(_22078_),
    .ZN(_05573_)
  );
  INV_X1 _39964_ (
    .A(_05573_),
    .ZN(_05574_)
  );
  AND2_X1 _39965_ (
    .A1(\cpuregs[15] [3]),
    .A2(_00007_[1]),
    .ZN(_05575_)
  );
  INV_X1 _39966_ (
    .A(_05575_),
    .ZN(_05576_)
  );
  AND2_X1 _39967_ (
    .A1(_00007_[2]),
    .A2(_05576_),
    .ZN(_05577_)
  );
  AND2_X1 _39968_ (
    .A1(_05574_),
    .A2(_05577_),
    .ZN(_05578_)
  );
  INV_X1 _39969_ (
    .A(_05578_),
    .ZN(_05579_)
  );
  AND2_X1 _39970_ (
    .A1(\cpuregs[9] [3]),
    .A2(_22078_),
    .ZN(_05580_)
  );
  INV_X1 _39971_ (
    .A(_05580_),
    .ZN(_05581_)
  );
  AND2_X1 _39972_ (
    .A1(\cpuregs[11] [3]),
    .A2(_00007_[1]),
    .ZN(_05582_)
  );
  INV_X1 _39973_ (
    .A(_05582_),
    .ZN(_05583_)
  );
  AND2_X1 _39974_ (
    .A1(_22077_),
    .A2(_05583_),
    .ZN(_05584_)
  );
  AND2_X1 _39975_ (
    .A1(_05581_),
    .A2(_05584_),
    .ZN(_05585_)
  );
  INV_X1 _39976_ (
    .A(_05585_),
    .ZN(_05586_)
  );
  AND2_X1 _39977_ (
    .A1(_00007_[0]),
    .A2(_05586_),
    .ZN(_05587_)
  );
  AND2_X1 _39978_ (
    .A1(_05579_),
    .A2(_05587_),
    .ZN(_05588_)
  );
  INV_X1 _39979_ (
    .A(_05588_),
    .ZN(_05589_)
  );
  AND2_X1 _39980_ (
    .A1(\cpuregs[12] [3]),
    .A2(_22078_),
    .ZN(_05590_)
  );
  INV_X1 _39981_ (
    .A(_05590_),
    .ZN(_05591_)
  );
  AND2_X1 _39982_ (
    .A1(\cpuregs[14] [3]),
    .A2(_00007_[1]),
    .ZN(_05592_)
  );
  INV_X1 _39983_ (
    .A(_05592_),
    .ZN(_05593_)
  );
  AND2_X1 _39984_ (
    .A1(_00007_[2]),
    .A2(_05593_),
    .ZN(_05594_)
  );
  AND2_X1 _39985_ (
    .A1(_05591_),
    .A2(_05594_),
    .ZN(_05595_)
  );
  INV_X1 _39986_ (
    .A(_05595_),
    .ZN(_05596_)
  );
  AND2_X1 _39987_ (
    .A1(\cpuregs[8] [3]),
    .A2(_22078_),
    .ZN(_05597_)
  );
  INV_X1 _39988_ (
    .A(_05597_),
    .ZN(_05598_)
  );
  AND2_X1 _39989_ (
    .A1(\cpuregs[10] [3]),
    .A2(_00007_[1]),
    .ZN(_05599_)
  );
  INV_X1 _39990_ (
    .A(_05599_),
    .ZN(_05600_)
  );
  AND2_X1 _39991_ (
    .A1(_22077_),
    .A2(_05600_),
    .ZN(_05601_)
  );
  AND2_X1 _39992_ (
    .A1(_05598_),
    .A2(_05601_),
    .ZN(_05602_)
  );
  INV_X1 _39993_ (
    .A(_05602_),
    .ZN(_05603_)
  );
  AND2_X1 _39994_ (
    .A1(_22152_),
    .A2(_05603_),
    .ZN(_05604_)
  );
  AND2_X1 _39995_ (
    .A1(_05596_),
    .A2(_05604_),
    .ZN(_05605_)
  );
  INV_X1 _39996_ (
    .A(_05605_),
    .ZN(_05606_)
  );
  AND2_X1 _39997_ (
    .A1(_05589_),
    .A2(_05606_),
    .ZN(_05607_)
  );
  INV_X1 _39998_ (
    .A(_05607_),
    .ZN(_05608_)
  );
  AND2_X1 _39999_ (
    .A1(_00007_[3]),
    .A2(_05608_),
    .ZN(_05609_)
  );
  INV_X1 _40000_ (
    .A(_05609_),
    .ZN(_05610_)
  );
  AND2_X1 _40001_ (
    .A1(_21540_),
    .A2(_22077_),
    .ZN(_05611_)
  );
  INV_X1 _40002_ (
    .A(_05611_),
    .ZN(_05612_)
  );
  AND2_X1 _40003_ (
    .A1(_21807_),
    .A2(_00007_[2]),
    .ZN(_05613_)
  );
  INV_X1 _40004_ (
    .A(_05613_),
    .ZN(_05614_)
  );
  AND2_X1 _40005_ (
    .A1(_22152_),
    .A2(_05614_),
    .ZN(_05615_)
  );
  AND2_X1 _40006_ (
    .A1(_05612_),
    .A2(_05615_),
    .ZN(_05616_)
  );
  INV_X1 _40007_ (
    .A(_05616_),
    .ZN(_05617_)
  );
  AND2_X1 _40008_ (
    .A1(_21782_),
    .A2(_00007_[2]),
    .ZN(_05618_)
  );
  INV_X1 _40009_ (
    .A(_05618_),
    .ZN(_05619_)
  );
  AND2_X1 _40010_ (
    .A1(_21490_),
    .A2(_22077_),
    .ZN(_05620_)
  );
  INV_X1 _40011_ (
    .A(_05620_),
    .ZN(_05621_)
  );
  AND2_X1 _40012_ (
    .A1(_00007_[0]),
    .A2(_05621_),
    .ZN(_05622_)
  );
  AND2_X1 _40013_ (
    .A1(_05619_),
    .A2(_05622_),
    .ZN(_05623_)
  );
  INV_X1 _40014_ (
    .A(_05623_),
    .ZN(_05624_)
  );
  AND2_X1 _40015_ (
    .A1(_05617_),
    .A2(_05624_),
    .ZN(_05625_)
  );
  AND2_X1 _40016_ (
    .A1(_21672_),
    .A2(_00007_[2]),
    .ZN(_05626_)
  );
  INV_X1 _40017_ (
    .A(_05626_),
    .ZN(_05627_)
  );
  AND2_X1 _40018_ (
    .A1(_21956_),
    .A2(_22077_),
    .ZN(_05628_)
  );
  INV_X1 _40019_ (
    .A(_05628_),
    .ZN(_05629_)
  );
  AND2_X1 _40020_ (
    .A1(_05627_),
    .A2(_05629_),
    .ZN(_05630_)
  );
  AND2_X1 _40021_ (
    .A1(_22152_),
    .A2(_05630_),
    .ZN(_05631_)
  );
  INV_X1 _40022_ (
    .A(_05631_),
    .ZN(_05632_)
  );
  AND2_X1 _40023_ (
    .A1(_21735_),
    .A2(_00007_[2]),
    .ZN(_05633_)
  );
  INV_X1 _40024_ (
    .A(_05633_),
    .ZN(_05634_)
  );
  AND2_X1 _40025_ (
    .A1(_21515_),
    .A2(_22077_),
    .ZN(_05635_)
  );
  INV_X1 _40026_ (
    .A(_05635_),
    .ZN(_05636_)
  );
  AND2_X1 _40027_ (
    .A1(_00007_[0]),
    .A2(_05636_),
    .ZN(_05637_)
  );
  AND2_X1 _40028_ (
    .A1(_05634_),
    .A2(_05637_),
    .ZN(_05638_)
  );
  INV_X1 _40029_ (
    .A(_05638_),
    .ZN(_05639_)
  );
  AND2_X1 _40030_ (
    .A1(_05632_),
    .A2(_05639_),
    .ZN(_05640_)
  );
  AND2_X1 _40031_ (
    .A1(_00007_[1]),
    .A2(_05625_),
    .ZN(_05641_)
  );
  INV_X1 _40032_ (
    .A(_05641_),
    .ZN(_05642_)
  );
  AND2_X1 _40033_ (
    .A1(_22078_),
    .A2(_05640_),
    .ZN(_05643_)
  );
  INV_X1 _40034_ (
    .A(_05643_),
    .ZN(_05644_)
  );
  AND2_X1 _40035_ (
    .A1(_05642_),
    .A2(_05644_),
    .ZN(_05645_)
  );
  AND2_X1 _40036_ (
    .A1(_22109_),
    .A2(_05645_),
    .ZN(_05646_)
  );
  INV_X1 _40037_ (
    .A(_05646_),
    .ZN(_05647_)
  );
  AND2_X1 _40038_ (
    .A1(_05610_),
    .A2(_05647_),
    .ZN(_05648_)
  );
  AND2_X1 _40039_ (
    .A1(_00007_[4]),
    .A2(_05572_),
    .ZN(_05649_)
  );
  INV_X1 _40040_ (
    .A(_05649_),
    .ZN(_05650_)
  );
  AND2_X1 _40041_ (
    .A1(_22144_),
    .A2(_05648_),
    .ZN(_05651_)
  );
  INV_X1 _40042_ (
    .A(_05651_),
    .ZN(_05652_)
  );
  AND2_X1 _40043_ (
    .A1(_04974_),
    .A2(_05652_),
    .ZN(_05653_)
  );
  AND2_X1 _40044_ (
    .A1(_05650_),
    .A2(_05653_),
    .ZN(_05654_)
  );
  AND2_X1 _40045_ (
    .A1(_04958_),
    .A2(_05654_),
    .ZN(_05655_)
  );
  INV_X1 _40046_ (
    .A(_05655_),
    .ZN(_05656_)
  );
  AND2_X1 _40047_ (
    .A1(_05137_),
    .A2(_05654_),
    .ZN(_05657_)
  );
  INV_X1 _40048_ (
    .A(_05657_),
    .ZN(_05658_)
  );
  AND2_X1 _40049_ (
    .A1(_05656_),
    .A2(_05658_),
    .ZN(_05659_)
  );
  AND2_X1 _40050_ (
    .A1(_05490_),
    .A2(_05659_),
    .ZN(_05660_)
  );
  AND2_X1 _40051_ (
    .A1(_21203_),
    .A2(_04963_),
    .ZN(_05661_)
  );
  INV_X1 _40052_ (
    .A(_05661_),
    .ZN(_05662_)
  );
  AND2_X1 _40053_ (
    .A1(_04962_),
    .A2(_05660_),
    .ZN(_05663_)
  );
  INV_X1 _40054_ (
    .A(_05663_),
    .ZN(_05664_)
  );
  AND2_X1 _40055_ (
    .A1(_05662_),
    .A2(_05664_),
    .ZN(_00284_)
  );
  AND2_X1 _40056_ (
    .A1(decoded_imm[4]),
    .A2(_04966_),
    .ZN(_05665_)
  );
  INV_X1 _40057_ (
    .A(_05665_),
    .ZN(_05666_)
  );
  AND2_X1 _40058_ (
    .A1(_21440_),
    .A2(_22077_),
    .ZN(_05667_)
  );
  INV_X1 _40059_ (
    .A(_05667_),
    .ZN(_05668_)
  );
  AND2_X1 _40060_ (
    .A1(_21651_),
    .A2(_00007_[2]),
    .ZN(_05669_)
  );
  INV_X1 _40061_ (
    .A(_05669_),
    .ZN(_05670_)
  );
  AND2_X1 _40062_ (
    .A1(_05668_),
    .A2(_05670_),
    .ZN(_05671_)
  );
  AND2_X1 _40063_ (
    .A1(_21594_),
    .A2(_22077_),
    .ZN(_05672_)
  );
  INV_X1 _40064_ (
    .A(_05672_),
    .ZN(_05673_)
  );
  AND2_X1 _40065_ (
    .A1(_21412_),
    .A2(_00007_[2]),
    .ZN(_05674_)
  );
  INV_X1 _40066_ (
    .A(_05674_),
    .ZN(_05675_)
  );
  AND2_X1 _40067_ (
    .A1(_21462_),
    .A2(_22077_),
    .ZN(_05676_)
  );
  INV_X1 _40068_ (
    .A(_05676_),
    .ZN(_05677_)
  );
  AND2_X1 _40069_ (
    .A1(_21761_),
    .A2(_00007_[2]),
    .ZN(_05678_)
  );
  INV_X1 _40070_ (
    .A(_05678_),
    .ZN(_05679_)
  );
  AND2_X1 _40071_ (
    .A1(_21374_),
    .A2(_00007_[2]),
    .ZN(_05680_)
  );
  INV_X1 _40072_ (
    .A(_05680_),
    .ZN(_05681_)
  );
  AND2_X1 _40073_ (
    .A1(_21620_),
    .A2(_22077_),
    .ZN(_05682_)
  );
  INV_X1 _40074_ (
    .A(_05682_),
    .ZN(_05683_)
  );
  AND2_X1 _40075_ (
    .A1(_00007_[0]),
    .A2(_05683_),
    .ZN(_05684_)
  );
  AND2_X1 _40076_ (
    .A1(_05681_),
    .A2(_05684_),
    .ZN(_05685_)
  );
  INV_X1 _40077_ (
    .A(_05685_),
    .ZN(_05686_)
  );
  AND2_X1 _40078_ (
    .A1(_22152_),
    .A2(_05673_),
    .ZN(_05687_)
  );
  AND2_X1 _40079_ (
    .A1(_05675_),
    .A2(_05687_),
    .ZN(_05688_)
  );
  INV_X1 _40080_ (
    .A(_05688_),
    .ZN(_05689_)
  );
  AND2_X1 _40081_ (
    .A1(_05686_),
    .A2(_05689_),
    .ZN(_05690_)
  );
  AND2_X1 _40082_ (
    .A1(_00007_[1]),
    .A2(_05690_),
    .ZN(_05691_)
  );
  INV_X1 _40083_ (
    .A(_05691_),
    .ZN(_05692_)
  );
  AND2_X1 _40084_ (
    .A1(_00007_[0]),
    .A2(_05677_),
    .ZN(_05693_)
  );
  AND2_X1 _40085_ (
    .A1(_05679_),
    .A2(_05693_),
    .ZN(_05694_)
  );
  INV_X1 _40086_ (
    .A(_05694_),
    .ZN(_05695_)
  );
  AND2_X1 _40087_ (
    .A1(_22152_),
    .A2(_05671_),
    .ZN(_05696_)
  );
  INV_X1 _40088_ (
    .A(_05696_),
    .ZN(_05697_)
  );
  AND2_X1 _40089_ (
    .A1(_05695_),
    .A2(_05697_),
    .ZN(_05698_)
  );
  AND2_X1 _40090_ (
    .A1(_22078_),
    .A2(_05698_),
    .ZN(_05699_)
  );
  INV_X1 _40091_ (
    .A(_05699_),
    .ZN(_05700_)
  );
  AND2_X1 _40092_ (
    .A1(_22109_),
    .A2(_05700_),
    .ZN(_05701_)
  );
  AND2_X1 _40093_ (
    .A1(_05692_),
    .A2(_05701_),
    .ZN(_05702_)
  );
  INV_X1 _40094_ (
    .A(_05702_),
    .ZN(_05703_)
  );
  AND2_X1 _40095_ (
    .A1(\cpuregs[27] [4]),
    .A2(_00007_[1]),
    .ZN(_05704_)
  );
  INV_X1 _40096_ (
    .A(_05704_),
    .ZN(_05705_)
  );
  AND2_X1 _40097_ (
    .A1(\cpuregs[25] [4]),
    .A2(_22078_),
    .ZN(_05706_)
  );
  INV_X1 _40098_ (
    .A(_05706_),
    .ZN(_05707_)
  );
  AND2_X1 _40099_ (
    .A1(_05705_),
    .A2(_05707_),
    .ZN(_05708_)
  );
  INV_X1 _40100_ (
    .A(_05708_),
    .ZN(_05709_)
  );
  AND2_X1 _40101_ (
    .A1(_22077_),
    .A2(_05709_),
    .ZN(_05710_)
  );
  INV_X1 _40102_ (
    .A(_05710_),
    .ZN(_05711_)
  );
  AND2_X1 _40103_ (
    .A1(\cpuregs[31] [4]),
    .A2(_00007_[1]),
    .ZN(_05712_)
  );
  INV_X1 _40104_ (
    .A(_05712_),
    .ZN(_05713_)
  );
  AND2_X1 _40105_ (
    .A1(\cpuregs[29] [4]),
    .A2(_22078_),
    .ZN(_05714_)
  );
  INV_X1 _40106_ (
    .A(_05714_),
    .ZN(_05715_)
  );
  AND2_X1 _40107_ (
    .A1(_05713_),
    .A2(_05715_),
    .ZN(_05716_)
  );
  INV_X1 _40108_ (
    .A(_05716_),
    .ZN(_05717_)
  );
  AND2_X1 _40109_ (
    .A1(_00007_[2]),
    .A2(_05717_),
    .ZN(_05718_)
  );
  INV_X1 _40110_ (
    .A(_05718_),
    .ZN(_05719_)
  );
  AND2_X1 _40111_ (
    .A1(_00007_[0]),
    .A2(_05719_),
    .ZN(_05720_)
  );
  AND2_X1 _40112_ (
    .A1(_05711_),
    .A2(_05720_),
    .ZN(_05721_)
  );
  INV_X1 _40113_ (
    .A(_05721_),
    .ZN(_05722_)
  );
  AND2_X1 _40114_ (
    .A1(\cpuregs[26] [4]),
    .A2(_00007_[1]),
    .ZN(_05723_)
  );
  INV_X1 _40115_ (
    .A(_05723_),
    .ZN(_05724_)
  );
  AND2_X1 _40116_ (
    .A1(\cpuregs[24] [4]),
    .A2(_22078_),
    .ZN(_05725_)
  );
  INV_X1 _40117_ (
    .A(_05725_),
    .ZN(_05726_)
  );
  AND2_X1 _40118_ (
    .A1(_05724_),
    .A2(_05726_),
    .ZN(_05727_)
  );
  INV_X1 _40119_ (
    .A(_05727_),
    .ZN(_05728_)
  );
  AND2_X1 _40120_ (
    .A1(_22077_),
    .A2(_05728_),
    .ZN(_05729_)
  );
  INV_X1 _40121_ (
    .A(_05729_),
    .ZN(_05730_)
  );
  AND2_X1 _40122_ (
    .A1(\cpuregs[30] [4]),
    .A2(_00007_[1]),
    .ZN(_05731_)
  );
  INV_X1 _40123_ (
    .A(_05731_),
    .ZN(_05732_)
  );
  AND2_X1 _40124_ (
    .A1(\cpuregs[28] [4]),
    .A2(_22078_),
    .ZN(_05733_)
  );
  INV_X1 _40125_ (
    .A(_05733_),
    .ZN(_05734_)
  );
  AND2_X1 _40126_ (
    .A1(_05732_),
    .A2(_05734_),
    .ZN(_05735_)
  );
  INV_X1 _40127_ (
    .A(_05735_),
    .ZN(_05736_)
  );
  AND2_X1 _40128_ (
    .A1(_00007_[2]),
    .A2(_05736_),
    .ZN(_05737_)
  );
  INV_X1 _40129_ (
    .A(_05737_),
    .ZN(_05738_)
  );
  AND2_X1 _40130_ (
    .A1(_22152_),
    .A2(_05738_),
    .ZN(_05739_)
  );
  AND2_X1 _40131_ (
    .A1(_05730_),
    .A2(_05739_),
    .ZN(_05740_)
  );
  INV_X1 _40132_ (
    .A(_05740_),
    .ZN(_05741_)
  );
  AND2_X1 _40133_ (
    .A1(_00007_[3]),
    .A2(_05741_),
    .ZN(_05742_)
  );
  AND2_X1 _40134_ (
    .A1(_05722_),
    .A2(_05742_),
    .ZN(_05743_)
  );
  INV_X1 _40135_ (
    .A(_05743_),
    .ZN(_05744_)
  );
  AND2_X1 _40136_ (
    .A1(_05703_),
    .A2(_05744_),
    .ZN(_05745_)
  );
  AND2_X1 _40137_ (
    .A1(\cpuregs[9] [4]),
    .A2(_22077_),
    .ZN(_05746_)
  );
  INV_X1 _40138_ (
    .A(_05746_),
    .ZN(_05747_)
  );
  AND2_X1 _40139_ (
    .A1(\cpuregs[13] [4]),
    .A2(_00007_[2]),
    .ZN(_05748_)
  );
  INV_X1 _40140_ (
    .A(_05748_),
    .ZN(_05749_)
  );
  AND2_X1 _40141_ (
    .A1(_00007_[0]),
    .A2(_05749_),
    .ZN(_05750_)
  );
  AND2_X1 _40142_ (
    .A1(_05747_),
    .A2(_05750_),
    .ZN(_05751_)
  );
  INV_X1 _40143_ (
    .A(_05751_),
    .ZN(_05752_)
  );
  AND2_X1 _40144_ (
    .A1(\cpuregs[8] [4]),
    .A2(_22077_),
    .ZN(_05753_)
  );
  INV_X1 _40145_ (
    .A(_05753_),
    .ZN(_05754_)
  );
  AND2_X1 _40146_ (
    .A1(\cpuregs[12] [4]),
    .A2(_00007_[2]),
    .ZN(_05755_)
  );
  INV_X1 _40147_ (
    .A(_05755_),
    .ZN(_05756_)
  );
  AND2_X1 _40148_ (
    .A1(_22152_),
    .A2(_05756_),
    .ZN(_05757_)
  );
  AND2_X1 _40149_ (
    .A1(_05754_),
    .A2(_05757_),
    .ZN(_05758_)
  );
  INV_X1 _40150_ (
    .A(_05758_),
    .ZN(_05759_)
  );
  AND2_X1 _40151_ (
    .A1(_22078_),
    .A2(_05759_),
    .ZN(_05760_)
  );
  AND2_X1 _40152_ (
    .A1(_05752_),
    .A2(_05760_),
    .ZN(_05761_)
  );
  INV_X1 _40153_ (
    .A(_05761_),
    .ZN(_05762_)
  );
  AND2_X1 _40154_ (
    .A1(\cpuregs[15] [4]),
    .A2(_00007_[2]),
    .ZN(_05763_)
  );
  INV_X1 _40155_ (
    .A(_05763_),
    .ZN(_05764_)
  );
  AND2_X1 _40156_ (
    .A1(\cpuregs[11] [4]),
    .A2(_22077_),
    .ZN(_05765_)
  );
  INV_X1 _40157_ (
    .A(_05765_),
    .ZN(_05766_)
  );
  AND2_X1 _40158_ (
    .A1(_00007_[0]),
    .A2(_05766_),
    .ZN(_05767_)
  );
  AND2_X1 _40159_ (
    .A1(_05764_),
    .A2(_05767_),
    .ZN(_05768_)
  );
  INV_X1 _40160_ (
    .A(_05768_),
    .ZN(_05769_)
  );
  AND2_X1 _40161_ (
    .A1(\cpuregs[14] [4]),
    .A2(_00007_[2]),
    .ZN(_05770_)
  );
  INV_X1 _40162_ (
    .A(_05770_),
    .ZN(_05771_)
  );
  AND2_X1 _40163_ (
    .A1(\cpuregs[10] [4]),
    .A2(_22077_),
    .ZN(_05772_)
  );
  INV_X1 _40164_ (
    .A(_05772_),
    .ZN(_05773_)
  );
  AND2_X1 _40165_ (
    .A1(_22152_),
    .A2(_05773_),
    .ZN(_05774_)
  );
  AND2_X1 _40166_ (
    .A1(_05771_),
    .A2(_05774_),
    .ZN(_05775_)
  );
  INV_X1 _40167_ (
    .A(_05775_),
    .ZN(_05776_)
  );
  AND2_X1 _40168_ (
    .A1(_00007_[1]),
    .A2(_05776_),
    .ZN(_05777_)
  );
  AND2_X1 _40169_ (
    .A1(_05769_),
    .A2(_05777_),
    .ZN(_05778_)
  );
  INV_X1 _40170_ (
    .A(_05778_),
    .ZN(_05779_)
  );
  AND2_X1 _40171_ (
    .A1(_05762_),
    .A2(_05779_),
    .ZN(_05780_)
  );
  INV_X1 _40172_ (
    .A(_05780_),
    .ZN(_05781_)
  );
  AND2_X1 _40173_ (
    .A1(_00007_[3]),
    .A2(_05781_),
    .ZN(_05782_)
  );
  INV_X1 _40174_ (
    .A(_05782_),
    .ZN(_05783_)
  );
  AND2_X1 _40175_ (
    .A1(_21783_),
    .A2(_00007_[2]),
    .ZN(_05784_)
  );
  INV_X1 _40176_ (
    .A(_05784_),
    .ZN(_05785_)
  );
  AND2_X1 _40177_ (
    .A1(_21491_),
    .A2(_22077_),
    .ZN(_05786_)
  );
  INV_X1 _40178_ (
    .A(_05786_),
    .ZN(_05787_)
  );
  AND2_X1 _40179_ (
    .A1(_00007_[0]),
    .A2(_05787_),
    .ZN(_05788_)
  );
  AND2_X1 _40180_ (
    .A1(_05785_),
    .A2(_05788_),
    .ZN(_05789_)
  );
  INV_X1 _40181_ (
    .A(_05789_),
    .ZN(_05790_)
  );
  AND2_X1 _40182_ (
    .A1(_21808_),
    .A2(_00007_[2]),
    .ZN(_05791_)
  );
  INV_X1 _40183_ (
    .A(_05791_),
    .ZN(_05792_)
  );
  AND2_X1 _40184_ (
    .A1(_21541_),
    .A2(_22077_),
    .ZN(_05793_)
  );
  INV_X1 _40185_ (
    .A(_05793_),
    .ZN(_05794_)
  );
  AND2_X1 _40186_ (
    .A1(_22152_),
    .A2(_05794_),
    .ZN(_05795_)
  );
  AND2_X1 _40187_ (
    .A1(_05792_),
    .A2(_05795_),
    .ZN(_05796_)
  );
  INV_X1 _40188_ (
    .A(_05796_),
    .ZN(_05797_)
  );
  AND2_X1 _40189_ (
    .A1(_05790_),
    .A2(_05797_),
    .ZN(_05798_)
  );
  AND2_X1 _40190_ (
    .A1(_00007_[1]),
    .A2(_05798_),
    .ZN(_05799_)
  );
  INV_X1 _40191_ (
    .A(_05799_),
    .ZN(_05800_)
  );
  AND2_X1 _40192_ (
    .A1(_21736_),
    .A2(_00007_[2]),
    .ZN(_05801_)
  );
  INV_X1 _40193_ (
    .A(_05801_),
    .ZN(_05802_)
  );
  AND2_X1 _40194_ (
    .A1(_21516_),
    .A2(_22077_),
    .ZN(_05803_)
  );
  INV_X1 _40195_ (
    .A(_05803_),
    .ZN(_05804_)
  );
  AND2_X1 _40196_ (
    .A1(_00007_[0]),
    .A2(_05804_),
    .ZN(_05805_)
  );
  AND2_X1 _40197_ (
    .A1(_05802_),
    .A2(_05805_),
    .ZN(_05806_)
  );
  INV_X1 _40198_ (
    .A(_05806_),
    .ZN(_05807_)
  );
  AND2_X1 _40199_ (
    .A1(_21957_),
    .A2(_22077_),
    .ZN(_05808_)
  );
  INV_X1 _40200_ (
    .A(_05808_),
    .ZN(_05809_)
  );
  AND2_X1 _40201_ (
    .A1(_21673_),
    .A2(_00007_[2]),
    .ZN(_05810_)
  );
  INV_X1 _40202_ (
    .A(_05810_),
    .ZN(_05811_)
  );
  AND2_X1 _40203_ (
    .A1(_05809_),
    .A2(_05811_),
    .ZN(_05812_)
  );
  AND2_X1 _40204_ (
    .A1(_22152_),
    .A2(_05812_),
    .ZN(_05813_)
  );
  INV_X1 _40205_ (
    .A(_05813_),
    .ZN(_05814_)
  );
  AND2_X1 _40206_ (
    .A1(_05807_),
    .A2(_05814_),
    .ZN(_05815_)
  );
  AND2_X1 _40207_ (
    .A1(_22078_),
    .A2(_05815_),
    .ZN(_05816_)
  );
  INV_X1 _40208_ (
    .A(_05816_),
    .ZN(_05817_)
  );
  AND2_X1 _40209_ (
    .A1(_05800_),
    .A2(_05817_),
    .ZN(_05818_)
  );
  AND2_X1 _40210_ (
    .A1(_22109_),
    .A2(_05818_),
    .ZN(_05819_)
  );
  INV_X1 _40211_ (
    .A(_05819_),
    .ZN(_05820_)
  );
  AND2_X1 _40212_ (
    .A1(_00007_[4]),
    .A2(_05745_),
    .ZN(_05821_)
  );
  INV_X1 _40213_ (
    .A(_05821_),
    .ZN(_05822_)
  );
  AND2_X1 _40214_ (
    .A1(_22144_),
    .A2(_05820_),
    .ZN(_05823_)
  );
  AND2_X1 _40215_ (
    .A1(_05783_),
    .A2(_05823_),
    .ZN(_05824_)
  );
  INV_X1 _40216_ (
    .A(_05824_),
    .ZN(_05825_)
  );
  AND2_X1 _40217_ (
    .A1(_04974_),
    .A2(_05825_),
    .ZN(_05826_)
  );
  AND2_X1 _40218_ (
    .A1(_05822_),
    .A2(_05826_),
    .ZN(_05827_)
  );
  AND2_X1 _40219_ (
    .A1(_04958_),
    .A2(_05827_),
    .ZN(_05828_)
  );
  INV_X1 _40220_ (
    .A(_05828_),
    .ZN(_05829_)
  );
  AND2_X1 _40221_ (
    .A1(_05137_),
    .A2(_05827_),
    .ZN(_05830_)
  );
  INV_X1 _40222_ (
    .A(_05830_),
    .ZN(_05831_)
  );
  AND2_X1 _40223_ (
    .A1(_05829_),
    .A2(_05831_),
    .ZN(_05832_)
  );
  AND2_X1 _40224_ (
    .A1(_05666_),
    .A2(_05832_),
    .ZN(_05833_)
  );
  AND2_X1 _40225_ (
    .A1(_21204_),
    .A2(_04963_),
    .ZN(_05834_)
  );
  INV_X1 _40226_ (
    .A(_05834_),
    .ZN(_05835_)
  );
  AND2_X1 _40227_ (
    .A1(_04962_),
    .A2(_05833_),
    .ZN(_05836_)
  );
  INV_X1 _40228_ (
    .A(_05836_),
    .ZN(_05837_)
  );
  AND2_X1 _40229_ (
    .A1(_05835_),
    .A2(_05837_),
    .ZN(_00285_)
  );
  AND2_X1 _40230_ (
    .A1(decoded_imm[5]),
    .A2(_04966_),
    .ZN(_05838_)
  );
  INV_X1 _40231_ (
    .A(_05838_),
    .ZN(_05839_)
  );
  AND2_X1 _40232_ (
    .A1(_04959_),
    .A2(_05138_),
    .ZN(_05840_)
  );
  INV_X1 _40233_ (
    .A(_05840_),
    .ZN(_05841_)
  );
  AND2_X1 _40234_ (
    .A1(_04974_),
    .A2(_05841_),
    .ZN(_05842_)
  );
  AND2_X1 _40235_ (
    .A1(_21621_),
    .A2(_22077_),
    .ZN(_05843_)
  );
  INV_X1 _40236_ (
    .A(_05843_),
    .ZN(_05844_)
  );
  AND2_X1 _40237_ (
    .A1(_21375_),
    .A2(_00007_[2]),
    .ZN(_05845_)
  );
  INV_X1 _40238_ (
    .A(_05845_),
    .ZN(_05846_)
  );
  AND2_X1 _40239_ (
    .A1(_00007_[0]),
    .A2(_05844_),
    .ZN(_05847_)
  );
  AND2_X1 _40240_ (
    .A1(_05846_),
    .A2(_05847_),
    .ZN(_05848_)
  );
  INV_X1 _40241_ (
    .A(_05848_),
    .ZN(_05849_)
  );
  AND2_X1 _40242_ (
    .A1(_21595_),
    .A2(_22077_),
    .ZN(_05850_)
  );
  INV_X1 _40243_ (
    .A(_05850_),
    .ZN(_05851_)
  );
  AND2_X1 _40244_ (
    .A1(_21413_),
    .A2(_00007_[2]),
    .ZN(_05852_)
  );
  INV_X1 _40245_ (
    .A(_05852_),
    .ZN(_05853_)
  );
  AND2_X1 _40246_ (
    .A1(_22152_),
    .A2(_05853_),
    .ZN(_05854_)
  );
  AND2_X1 _40247_ (
    .A1(_05851_),
    .A2(_05854_),
    .ZN(_05855_)
  );
  INV_X1 _40248_ (
    .A(_05855_),
    .ZN(_05856_)
  );
  AND2_X1 _40249_ (
    .A1(_21762_),
    .A2(_00007_[2]),
    .ZN(_05857_)
  );
  INV_X1 _40250_ (
    .A(_05857_),
    .ZN(_05858_)
  );
  AND2_X1 _40251_ (
    .A1(_21463_),
    .A2(_22077_),
    .ZN(_05859_)
  );
  INV_X1 _40252_ (
    .A(_05859_),
    .ZN(_05860_)
  );
  AND2_X1 _40253_ (
    .A1(_00007_[0]),
    .A2(_05858_),
    .ZN(_05861_)
  );
  AND2_X1 _40254_ (
    .A1(_05860_),
    .A2(_05861_),
    .ZN(_05862_)
  );
  INV_X1 _40255_ (
    .A(_05862_),
    .ZN(_05863_)
  );
  AND2_X1 _40256_ (
    .A1(_21441_),
    .A2(_22077_),
    .ZN(_05864_)
  );
  INV_X1 _40257_ (
    .A(_05864_),
    .ZN(_05865_)
  );
  AND2_X1 _40258_ (
    .A1(_21652_),
    .A2(_00007_[2]),
    .ZN(_05866_)
  );
  INV_X1 _40259_ (
    .A(_05866_),
    .ZN(_05867_)
  );
  AND2_X1 _40260_ (
    .A1(_05865_),
    .A2(_05867_),
    .ZN(_05868_)
  );
  AND2_X1 _40261_ (
    .A1(_22152_),
    .A2(_05868_),
    .ZN(_05869_)
  );
  INV_X1 _40262_ (
    .A(_05869_),
    .ZN(_05870_)
  );
  AND2_X1 _40263_ (
    .A1(_21480_),
    .A2(_00007_[2]),
    .ZN(_05871_)
  );
  INV_X1 _40264_ (
    .A(_05871_),
    .ZN(_05872_)
  );
  AND2_X1 _40265_ (
    .A1(_21725_),
    .A2(_22077_),
    .ZN(_05873_)
  );
  INV_X1 _40266_ (
    .A(_05873_),
    .ZN(_05874_)
  );
  AND2_X1 _40267_ (
    .A1(_05872_),
    .A2(_05874_),
    .ZN(_05875_)
  );
  AND2_X1 _40268_ (
    .A1(_21717_),
    .A2(_22077_),
    .ZN(_05876_)
  );
  INV_X1 _40269_ (
    .A(_05876_),
    .ZN(_05877_)
  );
  AND2_X1 _40270_ (
    .A1(_21639_),
    .A2(_00007_[2]),
    .ZN(_05878_)
  );
  INV_X1 _40271_ (
    .A(_05878_),
    .ZN(_05879_)
  );
  AND2_X1 _40272_ (
    .A1(_21698_),
    .A2(_22077_),
    .ZN(_05880_)
  );
  INV_X1 _40273_ (
    .A(_05880_),
    .ZN(_05881_)
  );
  AND2_X1 _40274_ (
    .A1(_21393_),
    .A2(_00007_[2]),
    .ZN(_05882_)
  );
  INV_X1 _40275_ (
    .A(_05882_),
    .ZN(_05883_)
  );
  AND2_X1 _40276_ (
    .A1(_05881_),
    .A2(_05883_),
    .ZN(_05884_)
  );
  AND2_X1 _40277_ (
    .A1(_21583_),
    .A2(_22077_),
    .ZN(_05885_)
  );
  INV_X1 _40278_ (
    .A(_05885_),
    .ZN(_05886_)
  );
  AND2_X1 _40279_ (
    .A1(_21401_),
    .A2(_00007_[2]),
    .ZN(_05887_)
  );
  INV_X1 _40280_ (
    .A(_05887_),
    .ZN(_05888_)
  );
  AND2_X1 _40281_ (
    .A1(_00007_[0]),
    .A2(_05877_),
    .ZN(_05889_)
  );
  AND2_X1 _40282_ (
    .A1(_05879_),
    .A2(_05889_),
    .ZN(_05890_)
  );
  INV_X1 _40283_ (
    .A(_05890_),
    .ZN(_05891_)
  );
  AND2_X1 _40284_ (
    .A1(_22152_),
    .A2(_05875_),
    .ZN(_05892_)
  );
  INV_X1 _40285_ (
    .A(_05892_),
    .ZN(_05893_)
  );
  AND2_X1 _40286_ (
    .A1(_05891_),
    .A2(_05893_),
    .ZN(_05894_)
  );
  AND2_X1 _40287_ (
    .A1(_22078_),
    .A2(_05894_),
    .ZN(_05895_)
  );
  INV_X1 _40288_ (
    .A(_05895_),
    .ZN(_05896_)
  );
  AND2_X1 _40289_ (
    .A1(_22152_),
    .A2(_05884_),
    .ZN(_05897_)
  );
  INV_X1 _40290_ (
    .A(_05897_),
    .ZN(_05898_)
  );
  AND2_X1 _40291_ (
    .A1(_00007_[0]),
    .A2(_05888_),
    .ZN(_05899_)
  );
  AND2_X1 _40292_ (
    .A1(_05886_),
    .A2(_05899_),
    .ZN(_05900_)
  );
  INV_X1 _40293_ (
    .A(_05900_),
    .ZN(_05901_)
  );
  AND2_X1 _40294_ (
    .A1(_00007_[1]),
    .A2(_05901_),
    .ZN(_05902_)
  );
  AND2_X1 _40295_ (
    .A1(_05898_),
    .A2(_05902_),
    .ZN(_05903_)
  );
  INV_X1 _40296_ (
    .A(_05903_),
    .ZN(_05904_)
  );
  AND2_X1 _40297_ (
    .A1(_05896_),
    .A2(_05904_),
    .ZN(_05905_)
  );
  AND2_X1 _40298_ (
    .A1(_21492_),
    .A2(_22077_),
    .ZN(_05906_)
  );
  INV_X1 _40299_ (
    .A(_05906_),
    .ZN(_05907_)
  );
  AND2_X1 _40300_ (
    .A1(_21784_),
    .A2(_00007_[2]),
    .ZN(_05908_)
  );
  INV_X1 _40301_ (
    .A(_05908_),
    .ZN(_05909_)
  );
  AND2_X1 _40302_ (
    .A1(_00007_[0]),
    .A2(_05907_),
    .ZN(_05910_)
  );
  AND2_X1 _40303_ (
    .A1(_05909_),
    .A2(_05910_),
    .ZN(_05911_)
  );
  INV_X1 _40304_ (
    .A(_05911_),
    .ZN(_05912_)
  );
  AND2_X1 _40305_ (
    .A1(_21542_),
    .A2(_22077_),
    .ZN(_05913_)
  );
  INV_X1 _40306_ (
    .A(_05913_),
    .ZN(_05914_)
  );
  AND2_X1 _40307_ (
    .A1(_21809_),
    .A2(_00007_[2]),
    .ZN(_05915_)
  );
  INV_X1 _40308_ (
    .A(_05915_),
    .ZN(_05916_)
  );
  AND2_X1 _40309_ (
    .A1(_22152_),
    .A2(_05916_),
    .ZN(_05917_)
  );
  AND2_X1 _40310_ (
    .A1(_05914_),
    .A2(_05917_),
    .ZN(_05918_)
  );
  INV_X1 _40311_ (
    .A(_05918_),
    .ZN(_05919_)
  );
  AND2_X1 _40312_ (
    .A1(_21737_),
    .A2(_00007_[2]),
    .ZN(_05920_)
  );
  INV_X1 _40313_ (
    .A(_05920_),
    .ZN(_05921_)
  );
  AND2_X1 _40314_ (
    .A1(_21517_),
    .A2(_22077_),
    .ZN(_05922_)
  );
  INV_X1 _40315_ (
    .A(_05922_),
    .ZN(_05923_)
  );
  AND2_X1 _40316_ (
    .A1(_00007_[0]),
    .A2(_05921_),
    .ZN(_05924_)
  );
  AND2_X1 _40317_ (
    .A1(_05923_),
    .A2(_05924_),
    .ZN(_05925_)
  );
  INV_X1 _40318_ (
    .A(_05925_),
    .ZN(_05926_)
  );
  AND2_X1 _40319_ (
    .A1(_21958_),
    .A2(_22077_),
    .ZN(_05927_)
  );
  INV_X1 _40320_ (
    .A(_05927_),
    .ZN(_05928_)
  );
  AND2_X1 _40321_ (
    .A1(_21674_),
    .A2(_00007_[2]),
    .ZN(_05929_)
  );
  INV_X1 _40322_ (
    .A(_05929_),
    .ZN(_05930_)
  );
  AND2_X1 _40323_ (
    .A1(_05928_),
    .A2(_05930_),
    .ZN(_05931_)
  );
  AND2_X1 _40324_ (
    .A1(_22152_),
    .A2(_05931_),
    .ZN(_05932_)
  );
  INV_X1 _40325_ (
    .A(_05932_),
    .ZN(_05933_)
  );
  AND2_X1 _40326_ (
    .A1(_05926_),
    .A2(_05933_),
    .ZN(_05934_)
  );
  AND2_X1 _40327_ (
    .A1(_22078_),
    .A2(_05934_),
    .ZN(_05935_)
  );
  INV_X1 _40328_ (
    .A(_05935_),
    .ZN(_05936_)
  );
  AND2_X1 _40329_ (
    .A1(_00007_[1]),
    .A2(_05919_),
    .ZN(_05937_)
  );
  AND2_X1 _40330_ (
    .A1(_05912_),
    .A2(_05937_),
    .ZN(_05938_)
  );
  INV_X1 _40331_ (
    .A(_05938_),
    .ZN(_05939_)
  );
  AND2_X1 _40332_ (
    .A1(_05936_),
    .A2(_05939_),
    .ZN(_05940_)
  );
  AND2_X1 _40333_ (
    .A1(_22144_),
    .A2(_05905_),
    .ZN(_05941_)
  );
  INV_X1 _40334_ (
    .A(_05941_),
    .ZN(_05942_)
  );
  AND2_X1 _40335_ (
    .A1(_21924_),
    .A2(_22077_),
    .ZN(_05943_)
  );
  INV_X1 _40336_ (
    .A(_05943_),
    .ZN(_05944_)
  );
  AND2_X1 _40337_ (
    .A1(_21940_),
    .A2(_00007_[2]),
    .ZN(_05945_)
  );
  INV_X1 _40338_ (
    .A(_05945_),
    .ZN(_05946_)
  );
  AND2_X1 _40339_ (
    .A1(_00007_[0]),
    .A2(_05946_),
    .ZN(_05947_)
  );
  AND2_X1 _40340_ (
    .A1(_05944_),
    .A2(_05947_),
    .ZN(_05948_)
  );
  INV_X1 _40341_ (
    .A(_05948_),
    .ZN(_05949_)
  );
  AND2_X1 _40342_ (
    .A1(_21852_),
    .A2(_00007_[2]),
    .ZN(_05950_)
  );
  INV_X1 _40343_ (
    .A(_05950_),
    .ZN(_05951_)
  );
  AND2_X1 _40344_ (
    .A1(_21868_),
    .A2(_22077_),
    .ZN(_05952_)
  );
  INV_X1 _40345_ (
    .A(_05952_),
    .ZN(_05953_)
  );
  AND2_X1 _40346_ (
    .A1(_05951_),
    .A2(_05953_),
    .ZN(_05954_)
  );
  AND2_X1 _40347_ (
    .A1(_22152_),
    .A2(_05954_),
    .ZN(_05955_)
  );
  INV_X1 _40348_ (
    .A(_05955_),
    .ZN(_05956_)
  );
  AND2_X1 _40349_ (
    .A1(_00007_[1]),
    .A2(_05949_),
    .ZN(_05957_)
  );
  AND2_X1 _40350_ (
    .A1(_05956_),
    .A2(_05957_),
    .ZN(_05958_)
  );
  INV_X1 _40351_ (
    .A(_05958_),
    .ZN(_05959_)
  );
  AND2_X1 _40352_ (
    .A1(_21892_),
    .A2(_00007_[2]),
    .ZN(_05960_)
  );
  INV_X1 _40353_ (
    .A(_05960_),
    .ZN(_05961_)
  );
  AND2_X1 _40354_ (
    .A1(_21836_),
    .A2(_22077_),
    .ZN(_05962_)
  );
  INV_X1 _40355_ (
    .A(_05962_),
    .ZN(_05963_)
  );
  AND2_X1 _40356_ (
    .A1(_00007_[0]),
    .A2(_05963_),
    .ZN(_05964_)
  );
  AND2_X1 _40357_ (
    .A1(_05961_),
    .A2(_05964_),
    .ZN(_05965_)
  );
  INV_X1 _40358_ (
    .A(_05965_),
    .ZN(_05966_)
  );
  AND2_X1 _40359_ (
    .A1(_21570_),
    .A2(_22077_),
    .ZN(_05967_)
  );
  INV_X1 _40360_ (
    .A(_05967_),
    .ZN(_05968_)
  );
  AND2_X1 _40361_ (
    .A1(_21908_),
    .A2(_00007_[2]),
    .ZN(_05969_)
  );
  INV_X1 _40362_ (
    .A(_05969_),
    .ZN(_05970_)
  );
  AND2_X1 _40363_ (
    .A1(_05968_),
    .A2(_05970_),
    .ZN(_05971_)
  );
  AND2_X1 _40364_ (
    .A1(_22152_),
    .A2(_05971_),
    .ZN(_05972_)
  );
  INV_X1 _40365_ (
    .A(_05972_),
    .ZN(_05973_)
  );
  AND2_X1 _40366_ (
    .A1(_22078_),
    .A2(_05973_),
    .ZN(_05974_)
  );
  AND2_X1 _40367_ (
    .A1(_05966_),
    .A2(_05974_),
    .ZN(_05975_)
  );
  INV_X1 _40368_ (
    .A(_05975_),
    .ZN(_05976_)
  );
  AND2_X1 _40369_ (
    .A1(_00007_[4]),
    .A2(_05976_),
    .ZN(_05977_)
  );
  AND2_X1 _40370_ (
    .A1(_05959_),
    .A2(_05977_),
    .ZN(_05978_)
  );
  INV_X1 _40371_ (
    .A(_05978_),
    .ZN(_05979_)
  );
  AND2_X1 _40372_ (
    .A1(_05942_),
    .A2(_05979_),
    .ZN(_05980_)
  );
  AND2_X1 _40373_ (
    .A1(_00007_[3]),
    .A2(_05980_),
    .ZN(_05981_)
  );
  INV_X1 _40374_ (
    .A(_05981_),
    .ZN(_05982_)
  );
  AND2_X1 _40375_ (
    .A1(_00007_[1]),
    .A2(_05856_),
    .ZN(_05983_)
  );
  AND2_X1 _40376_ (
    .A1(_05849_),
    .A2(_05983_),
    .ZN(_05984_)
  );
  INV_X1 _40377_ (
    .A(_05984_),
    .ZN(_05985_)
  );
  AND2_X1 _40378_ (
    .A1(_22078_),
    .A2(_05870_),
    .ZN(_05986_)
  );
  AND2_X1 _40379_ (
    .A1(_05863_),
    .A2(_05986_),
    .ZN(_05987_)
  );
  INV_X1 _40380_ (
    .A(_05987_),
    .ZN(_05988_)
  );
  AND2_X1 _40381_ (
    .A1(_00007_[4]),
    .A2(_05988_),
    .ZN(_05989_)
  );
  AND2_X1 _40382_ (
    .A1(_05985_),
    .A2(_05989_),
    .ZN(_05990_)
  );
  INV_X1 _40383_ (
    .A(_05990_),
    .ZN(_05991_)
  );
  AND2_X1 _40384_ (
    .A1(_22144_),
    .A2(_05940_),
    .ZN(_05992_)
  );
  INV_X1 _40385_ (
    .A(_05992_),
    .ZN(_05993_)
  );
  AND2_X1 _40386_ (
    .A1(_05991_),
    .A2(_05993_),
    .ZN(_05994_)
  );
  AND2_X1 _40387_ (
    .A1(_22109_),
    .A2(_05994_),
    .ZN(_05995_)
  );
  INV_X1 _40388_ (
    .A(_05995_),
    .ZN(_05996_)
  );
  AND2_X1 _40389_ (
    .A1(_05982_),
    .A2(_05996_),
    .ZN(_05997_)
  );
  AND2_X1 _40390_ (
    .A1(_05842_),
    .A2(_05997_),
    .ZN(_05998_)
  );
  INV_X1 _40391_ (
    .A(_05998_),
    .ZN(_05999_)
  );
  AND2_X1 _40392_ (
    .A1(_21205_),
    .A2(_04963_),
    .ZN(_06000_)
  );
  INV_X1 _40393_ (
    .A(_06000_),
    .ZN(_06001_)
  );
  AND2_X1 _40394_ (
    .A1(_04962_),
    .A2(_05999_),
    .ZN(_06002_)
  );
  AND2_X1 _40395_ (
    .A1(_05839_),
    .A2(_06002_),
    .ZN(_06003_)
  );
  INV_X1 _40396_ (
    .A(_06003_),
    .ZN(_06004_)
  );
  AND2_X1 _40397_ (
    .A1(_06001_),
    .A2(_06004_),
    .ZN(_00286_)
  );
  AND2_X1 _40398_ (
    .A1(decoded_imm[6]),
    .A2(_04966_),
    .ZN(_06005_)
  );
  INV_X1 _40399_ (
    .A(_06005_),
    .ZN(_06006_)
  );
  AND2_X1 _40400_ (
    .A1(_21893_),
    .A2(_00007_[2]),
    .ZN(_06007_)
  );
  INV_X1 _40401_ (
    .A(_06007_),
    .ZN(_06008_)
  );
  AND2_X1 _40402_ (
    .A1(_21837_),
    .A2(_22077_),
    .ZN(_06009_)
  );
  INV_X1 _40403_ (
    .A(_06009_),
    .ZN(_06010_)
  );
  AND2_X1 _40404_ (
    .A1(_00007_[0]),
    .A2(_06010_),
    .ZN(_06011_)
  );
  AND2_X1 _40405_ (
    .A1(_06008_),
    .A2(_06011_),
    .ZN(_06012_)
  );
  INV_X1 _40406_ (
    .A(_06012_),
    .ZN(_06013_)
  );
  AND2_X1 _40407_ (
    .A1(_21571_),
    .A2(_22077_),
    .ZN(_06014_)
  );
  INV_X1 _40408_ (
    .A(_06014_),
    .ZN(_06015_)
  );
  AND2_X1 _40409_ (
    .A1(_21909_),
    .A2(_00007_[2]),
    .ZN(_06016_)
  );
  INV_X1 _40410_ (
    .A(_06016_),
    .ZN(_06017_)
  );
  AND2_X1 _40411_ (
    .A1(_06015_),
    .A2(_06017_),
    .ZN(_06018_)
  );
  AND2_X1 _40412_ (
    .A1(_22152_),
    .A2(_06018_),
    .ZN(_06019_)
  );
  INV_X1 _40413_ (
    .A(_06019_),
    .ZN(_06020_)
  );
  AND2_X1 _40414_ (
    .A1(_06013_),
    .A2(_06020_),
    .ZN(_06021_)
  );
  AND2_X1 _40415_ (
    .A1(_22078_),
    .A2(_06021_),
    .ZN(_06022_)
  );
  INV_X1 _40416_ (
    .A(_06022_),
    .ZN(_06023_)
  );
  AND2_X1 _40417_ (
    .A1(_21869_),
    .A2(_22077_),
    .ZN(_06024_)
  );
  INV_X1 _40418_ (
    .A(_06024_),
    .ZN(_06025_)
  );
  AND2_X1 _40419_ (
    .A1(_21853_),
    .A2(_00007_[2]),
    .ZN(_06026_)
  );
  INV_X1 _40420_ (
    .A(_06026_),
    .ZN(_06027_)
  );
  AND2_X1 _40421_ (
    .A1(_06025_),
    .A2(_06027_),
    .ZN(_06028_)
  );
  AND2_X1 _40422_ (
    .A1(_22152_),
    .A2(_06028_),
    .ZN(_06029_)
  );
  INV_X1 _40423_ (
    .A(_06029_),
    .ZN(_06030_)
  );
  AND2_X1 _40424_ (
    .A1(_21941_),
    .A2(_00007_[2]),
    .ZN(_06031_)
  );
  INV_X1 _40425_ (
    .A(_06031_),
    .ZN(_06032_)
  );
  AND2_X1 _40426_ (
    .A1(_21925_),
    .A2(_22077_),
    .ZN(_06033_)
  );
  INV_X1 _40427_ (
    .A(_06033_),
    .ZN(_06034_)
  );
  AND2_X1 _40428_ (
    .A1(_00007_[0]),
    .A2(_06034_),
    .ZN(_06035_)
  );
  AND2_X1 _40429_ (
    .A1(_06032_),
    .A2(_06035_),
    .ZN(_06036_)
  );
  INV_X1 _40430_ (
    .A(_06036_),
    .ZN(_06037_)
  );
  AND2_X1 _40431_ (
    .A1(_06030_),
    .A2(_06037_),
    .ZN(_06038_)
  );
  AND2_X1 _40432_ (
    .A1(_00007_[1]),
    .A2(_06038_),
    .ZN(_06039_)
  );
  INV_X1 _40433_ (
    .A(_06039_),
    .ZN(_06040_)
  );
  AND2_X1 _40434_ (
    .A1(_00007_[3]),
    .A2(_06023_),
    .ZN(_06041_)
  );
  AND2_X1 _40435_ (
    .A1(_06040_),
    .A2(_06041_),
    .ZN(_06042_)
  );
  INV_X1 _40436_ (
    .A(_06042_),
    .ZN(_06043_)
  );
  AND2_X1 _40437_ (
    .A1(\cpuregs[17] [6]),
    .A2(_22077_),
    .ZN(_06044_)
  );
  INV_X1 _40438_ (
    .A(_06044_),
    .ZN(_06045_)
  );
  AND2_X1 _40439_ (
    .A1(\cpuregs[21] [6]),
    .A2(_00007_[2]),
    .ZN(_06046_)
  );
  INV_X1 _40440_ (
    .A(_06046_),
    .ZN(_06047_)
  );
  AND2_X1 _40441_ (
    .A1(_00007_[0]),
    .A2(_06047_),
    .ZN(_06048_)
  );
  AND2_X1 _40442_ (
    .A1(_06045_),
    .A2(_06048_),
    .ZN(_06049_)
  );
  INV_X1 _40443_ (
    .A(_06049_),
    .ZN(_06050_)
  );
  AND2_X1 _40444_ (
    .A1(\cpuregs[16] [6]),
    .A2(_22077_),
    .ZN(_06051_)
  );
  INV_X1 _40445_ (
    .A(_06051_),
    .ZN(_06052_)
  );
  AND2_X1 _40446_ (
    .A1(\cpuregs[20] [6]),
    .A2(_00007_[2]),
    .ZN(_06053_)
  );
  INV_X1 _40447_ (
    .A(_06053_),
    .ZN(_06054_)
  );
  AND2_X1 _40448_ (
    .A1(_22152_),
    .A2(_06054_),
    .ZN(_06055_)
  );
  AND2_X1 _40449_ (
    .A1(_06052_),
    .A2(_06055_),
    .ZN(_06056_)
  );
  INV_X1 _40450_ (
    .A(_06056_),
    .ZN(_06057_)
  );
  AND2_X1 _40451_ (
    .A1(_22078_),
    .A2(_06057_),
    .ZN(_06058_)
  );
  AND2_X1 _40452_ (
    .A1(_06050_),
    .A2(_06058_),
    .ZN(_06059_)
  );
  INV_X1 _40453_ (
    .A(_06059_),
    .ZN(_06060_)
  );
  AND2_X1 _40454_ (
    .A1(\cpuregs[19] [6]),
    .A2(_22077_),
    .ZN(_06061_)
  );
  INV_X1 _40455_ (
    .A(_06061_),
    .ZN(_06062_)
  );
  AND2_X1 _40456_ (
    .A1(\cpuregs[23] [6]),
    .A2(_00007_[2]),
    .ZN(_06063_)
  );
  INV_X1 _40457_ (
    .A(_06063_),
    .ZN(_06064_)
  );
  AND2_X1 _40458_ (
    .A1(_00007_[0]),
    .A2(_06064_),
    .ZN(_06065_)
  );
  AND2_X1 _40459_ (
    .A1(_06062_),
    .A2(_06065_),
    .ZN(_06066_)
  );
  INV_X1 _40460_ (
    .A(_06066_),
    .ZN(_06067_)
  );
  AND2_X1 _40461_ (
    .A1(\cpuregs[22] [6]),
    .A2(_00007_[2]),
    .ZN(_06068_)
  );
  INV_X1 _40462_ (
    .A(_06068_),
    .ZN(_06069_)
  );
  AND2_X1 _40463_ (
    .A1(\cpuregs[18] [6]),
    .A2(_22077_),
    .ZN(_06070_)
  );
  INV_X1 _40464_ (
    .A(_06070_),
    .ZN(_06071_)
  );
  AND2_X1 _40465_ (
    .A1(_22152_),
    .A2(_06071_),
    .ZN(_06072_)
  );
  AND2_X1 _40466_ (
    .A1(_06069_),
    .A2(_06072_),
    .ZN(_06073_)
  );
  INV_X1 _40467_ (
    .A(_06073_),
    .ZN(_06074_)
  );
  AND2_X1 _40468_ (
    .A1(_00007_[1]),
    .A2(_06074_),
    .ZN(_06075_)
  );
  AND2_X1 _40469_ (
    .A1(_06067_),
    .A2(_06075_),
    .ZN(_06076_)
  );
  INV_X1 _40470_ (
    .A(_06076_),
    .ZN(_06077_)
  );
  AND2_X1 _40471_ (
    .A1(_06060_),
    .A2(_06077_),
    .ZN(_06078_)
  );
  INV_X1 _40472_ (
    .A(_06078_),
    .ZN(_06079_)
  );
  AND2_X1 _40473_ (
    .A1(_22109_),
    .A2(_06079_),
    .ZN(_06080_)
  );
  INV_X1 _40474_ (
    .A(_06080_),
    .ZN(_06081_)
  );
  AND2_X1 _40475_ (
    .A1(_06043_),
    .A2(_06081_),
    .ZN(_06082_)
  );
  AND2_X1 _40476_ (
    .A1(_21640_),
    .A2(_00007_[2]),
    .ZN(_06083_)
  );
  INV_X1 _40477_ (
    .A(_06083_),
    .ZN(_06084_)
  );
  AND2_X1 _40478_ (
    .A1(_21718_),
    .A2(_22077_),
    .ZN(_06085_)
  );
  INV_X1 _40479_ (
    .A(_06085_),
    .ZN(_06086_)
  );
  AND2_X1 _40480_ (
    .A1(_00007_[0]),
    .A2(_06086_),
    .ZN(_06087_)
  );
  AND2_X1 _40481_ (
    .A1(_06084_),
    .A2(_06087_),
    .ZN(_06088_)
  );
  INV_X1 _40482_ (
    .A(_06088_),
    .ZN(_06089_)
  );
  AND2_X1 _40483_ (
    .A1(_21726_),
    .A2(_22077_),
    .ZN(_06090_)
  );
  INV_X1 _40484_ (
    .A(_06090_),
    .ZN(_06091_)
  );
  AND2_X1 _40485_ (
    .A1(_21481_),
    .A2(_00007_[2]),
    .ZN(_06092_)
  );
  INV_X1 _40486_ (
    .A(_06092_),
    .ZN(_06093_)
  );
  AND2_X1 _40487_ (
    .A1(_06091_),
    .A2(_06093_),
    .ZN(_06094_)
  );
  AND2_X1 _40488_ (
    .A1(_22152_),
    .A2(_06094_),
    .ZN(_06095_)
  );
  INV_X1 _40489_ (
    .A(_06095_),
    .ZN(_06096_)
  );
  AND2_X1 _40490_ (
    .A1(_06089_),
    .A2(_06096_),
    .ZN(_06097_)
  );
  AND2_X1 _40491_ (
    .A1(_22078_),
    .A2(_06097_),
    .ZN(_06098_)
  );
  INV_X1 _40492_ (
    .A(_06098_),
    .ZN(_06099_)
  );
  AND2_X1 _40493_ (
    .A1(_21699_),
    .A2(_22077_),
    .ZN(_06100_)
  );
  INV_X1 _40494_ (
    .A(_06100_),
    .ZN(_06101_)
  );
  AND2_X1 _40495_ (
    .A1(_21394_),
    .A2(_00007_[2]),
    .ZN(_06102_)
  );
  INV_X1 _40496_ (
    .A(_06102_),
    .ZN(_06103_)
  );
  AND2_X1 _40497_ (
    .A1(_06101_),
    .A2(_06103_),
    .ZN(_06104_)
  );
  AND2_X1 _40498_ (
    .A1(_22152_),
    .A2(_06104_),
    .ZN(_06105_)
  );
  INV_X1 _40499_ (
    .A(_06105_),
    .ZN(_06106_)
  );
  AND2_X1 _40500_ (
    .A1(_21402_),
    .A2(_00007_[2]),
    .ZN(_06107_)
  );
  INV_X1 _40501_ (
    .A(_06107_),
    .ZN(_06108_)
  );
  AND2_X1 _40502_ (
    .A1(_21584_),
    .A2(_22077_),
    .ZN(_06109_)
  );
  INV_X1 _40503_ (
    .A(_06109_),
    .ZN(_06110_)
  );
  AND2_X1 _40504_ (
    .A1(_00007_[0]),
    .A2(_06110_),
    .ZN(_06111_)
  );
  AND2_X1 _40505_ (
    .A1(_06108_),
    .A2(_06111_),
    .ZN(_06112_)
  );
  INV_X1 _40506_ (
    .A(_06112_),
    .ZN(_06113_)
  );
  AND2_X1 _40507_ (
    .A1(_06106_),
    .A2(_06113_),
    .ZN(_06114_)
  );
  AND2_X1 _40508_ (
    .A1(_00007_[1]),
    .A2(_06114_),
    .ZN(_06115_)
  );
  INV_X1 _40509_ (
    .A(_06115_),
    .ZN(_06116_)
  );
  AND2_X1 _40510_ (
    .A1(_00007_[3]),
    .A2(_06099_),
    .ZN(_06117_)
  );
  AND2_X1 _40511_ (
    .A1(_06116_),
    .A2(_06117_),
    .ZN(_06118_)
  );
  INV_X1 _40512_ (
    .A(_06118_),
    .ZN(_06119_)
  );
  AND2_X1 _40513_ (
    .A1(_21543_),
    .A2(_22077_),
    .ZN(_06120_)
  );
  INV_X1 _40514_ (
    .A(_06120_),
    .ZN(_06121_)
  );
  AND2_X1 _40515_ (
    .A1(_21810_),
    .A2(_00007_[2]),
    .ZN(_06122_)
  );
  INV_X1 _40516_ (
    .A(_06122_),
    .ZN(_06123_)
  );
  AND2_X1 _40517_ (
    .A1(_22152_),
    .A2(_06123_),
    .ZN(_06124_)
  );
  AND2_X1 _40518_ (
    .A1(_06121_),
    .A2(_06124_),
    .ZN(_06125_)
  );
  INV_X1 _40519_ (
    .A(_06125_),
    .ZN(_06126_)
  );
  AND2_X1 _40520_ (
    .A1(_21785_),
    .A2(_00007_[2]),
    .ZN(_06127_)
  );
  INV_X1 _40521_ (
    .A(_06127_),
    .ZN(_06128_)
  );
  AND2_X1 _40522_ (
    .A1(_21493_),
    .A2(_22077_),
    .ZN(_06129_)
  );
  INV_X1 _40523_ (
    .A(_06129_),
    .ZN(_06130_)
  );
  AND2_X1 _40524_ (
    .A1(_00007_[0]),
    .A2(_06130_),
    .ZN(_06131_)
  );
  AND2_X1 _40525_ (
    .A1(_06128_),
    .A2(_06131_),
    .ZN(_06132_)
  );
  INV_X1 _40526_ (
    .A(_06132_),
    .ZN(_06133_)
  );
  AND2_X1 _40527_ (
    .A1(_06126_),
    .A2(_06133_),
    .ZN(_06134_)
  );
  AND2_X1 _40528_ (
    .A1(_21675_),
    .A2(_00007_[2]),
    .ZN(_06135_)
  );
  INV_X1 _40529_ (
    .A(_06135_),
    .ZN(_06136_)
  );
  AND2_X1 _40530_ (
    .A1(_21959_),
    .A2(_22077_),
    .ZN(_06137_)
  );
  INV_X1 _40531_ (
    .A(_06137_),
    .ZN(_06138_)
  );
  AND2_X1 _40532_ (
    .A1(_06136_),
    .A2(_06138_),
    .ZN(_06139_)
  );
  AND2_X1 _40533_ (
    .A1(_22152_),
    .A2(_06139_),
    .ZN(_06140_)
  );
  INV_X1 _40534_ (
    .A(_06140_),
    .ZN(_06141_)
  );
  AND2_X1 _40535_ (
    .A1(_21738_),
    .A2(_00007_[2]),
    .ZN(_06142_)
  );
  INV_X1 _40536_ (
    .A(_06142_),
    .ZN(_06143_)
  );
  AND2_X1 _40537_ (
    .A1(_21518_),
    .A2(_22077_),
    .ZN(_06144_)
  );
  INV_X1 _40538_ (
    .A(_06144_),
    .ZN(_06145_)
  );
  AND2_X1 _40539_ (
    .A1(_00007_[0]),
    .A2(_06145_),
    .ZN(_06146_)
  );
  AND2_X1 _40540_ (
    .A1(_06143_),
    .A2(_06146_),
    .ZN(_06147_)
  );
  INV_X1 _40541_ (
    .A(_06147_),
    .ZN(_06148_)
  );
  AND2_X1 _40542_ (
    .A1(_06141_),
    .A2(_06148_),
    .ZN(_06149_)
  );
  AND2_X1 _40543_ (
    .A1(_00007_[1]),
    .A2(_06134_),
    .ZN(_06150_)
  );
  INV_X1 _40544_ (
    .A(_06150_),
    .ZN(_06151_)
  );
  AND2_X1 _40545_ (
    .A1(_22078_),
    .A2(_06149_),
    .ZN(_06152_)
  );
  INV_X1 _40546_ (
    .A(_06152_),
    .ZN(_06153_)
  );
  AND2_X1 _40547_ (
    .A1(_06151_),
    .A2(_06153_),
    .ZN(_06154_)
  );
  AND2_X1 _40548_ (
    .A1(_22109_),
    .A2(_06154_),
    .ZN(_06155_)
  );
  INV_X1 _40549_ (
    .A(_06155_),
    .ZN(_06156_)
  );
  AND2_X1 _40550_ (
    .A1(_06119_),
    .A2(_06156_),
    .ZN(_06157_)
  );
  AND2_X1 _40551_ (
    .A1(_00007_[4]),
    .A2(_06082_),
    .ZN(_06158_)
  );
  INV_X1 _40552_ (
    .A(_06158_),
    .ZN(_06159_)
  );
  AND2_X1 _40553_ (
    .A1(_22144_),
    .A2(_06157_),
    .ZN(_06160_)
  );
  INV_X1 _40554_ (
    .A(_06160_),
    .ZN(_06161_)
  );
  AND2_X1 _40555_ (
    .A1(_06159_),
    .A2(_06161_),
    .ZN(_06162_)
  );
  AND2_X1 _40556_ (
    .A1(_05842_),
    .A2(_06162_),
    .ZN(_06163_)
  );
  INV_X1 _40557_ (
    .A(_06163_),
    .ZN(_06164_)
  );
  AND2_X1 _40558_ (
    .A1(_06006_),
    .A2(_06164_),
    .ZN(_06165_)
  );
  AND2_X1 _40559_ (
    .A1(_04962_),
    .A2(_06165_),
    .ZN(_06166_)
  );
  INV_X1 _40560_ (
    .A(_06166_),
    .ZN(_06167_)
  );
  AND2_X1 _40561_ (
    .A1(_21206_),
    .A2(_04963_),
    .ZN(_06168_)
  );
  INV_X1 _40562_ (
    .A(_06168_),
    .ZN(_06169_)
  );
  AND2_X1 _40563_ (
    .A1(_06167_),
    .A2(_06169_),
    .ZN(_00287_)
  );
  AND2_X1 _40564_ (
    .A1(_21641_),
    .A2(_00007_[2]),
    .ZN(_06170_)
  );
  INV_X1 _40565_ (
    .A(_06170_),
    .ZN(_06171_)
  );
  AND2_X1 _40566_ (
    .A1(_21719_),
    .A2(_22077_),
    .ZN(_06172_)
  );
  INV_X1 _40567_ (
    .A(_06172_),
    .ZN(_06173_)
  );
  AND2_X1 _40568_ (
    .A1(_00007_[0]),
    .A2(_06173_),
    .ZN(_06174_)
  );
  AND2_X1 _40569_ (
    .A1(_06171_),
    .A2(_06174_),
    .ZN(_06175_)
  );
  INV_X1 _40570_ (
    .A(_06175_),
    .ZN(_06176_)
  );
  AND2_X1 _40571_ (
    .A1(_21727_),
    .A2(_22077_),
    .ZN(_06177_)
  );
  INV_X1 _40572_ (
    .A(_06177_),
    .ZN(_06178_)
  );
  AND2_X1 _40573_ (
    .A1(_21482_),
    .A2(_00007_[2]),
    .ZN(_06179_)
  );
  INV_X1 _40574_ (
    .A(_06179_),
    .ZN(_06180_)
  );
  AND2_X1 _40575_ (
    .A1(_06178_),
    .A2(_06180_),
    .ZN(_06181_)
  );
  AND2_X1 _40576_ (
    .A1(_22152_),
    .A2(_06181_),
    .ZN(_06182_)
  );
  INV_X1 _40577_ (
    .A(_06182_),
    .ZN(_06183_)
  );
  AND2_X1 _40578_ (
    .A1(_06176_),
    .A2(_06183_),
    .ZN(_06184_)
  );
  AND2_X1 _40579_ (
    .A1(_22078_),
    .A2(_06184_),
    .ZN(_06185_)
  );
  INV_X1 _40580_ (
    .A(_06185_),
    .ZN(_06186_)
  );
  AND2_X1 _40581_ (
    .A1(_21700_),
    .A2(_22077_),
    .ZN(_06187_)
  );
  INV_X1 _40582_ (
    .A(_06187_),
    .ZN(_06188_)
  );
  AND2_X1 _40583_ (
    .A1(_21395_),
    .A2(_00007_[2]),
    .ZN(_06189_)
  );
  INV_X1 _40584_ (
    .A(_06189_),
    .ZN(_06190_)
  );
  AND2_X1 _40585_ (
    .A1(_06188_),
    .A2(_06190_),
    .ZN(_06191_)
  );
  AND2_X1 _40586_ (
    .A1(_22152_),
    .A2(_06191_),
    .ZN(_06192_)
  );
  INV_X1 _40587_ (
    .A(_06192_),
    .ZN(_06193_)
  );
  AND2_X1 _40588_ (
    .A1(_21403_),
    .A2(_00007_[2]),
    .ZN(_06194_)
  );
  INV_X1 _40589_ (
    .A(_06194_),
    .ZN(_06195_)
  );
  AND2_X1 _40590_ (
    .A1(_21585_),
    .A2(_22077_),
    .ZN(_06196_)
  );
  INV_X1 _40591_ (
    .A(_06196_),
    .ZN(_06197_)
  );
  AND2_X1 _40592_ (
    .A1(_00007_[0]),
    .A2(_06197_),
    .ZN(_06198_)
  );
  AND2_X1 _40593_ (
    .A1(_06195_),
    .A2(_06198_),
    .ZN(_06199_)
  );
  INV_X1 _40594_ (
    .A(_06199_),
    .ZN(_06200_)
  );
  AND2_X1 _40595_ (
    .A1(_06193_),
    .A2(_06200_),
    .ZN(_06201_)
  );
  AND2_X1 _40596_ (
    .A1(_00007_[1]),
    .A2(_06201_),
    .ZN(_06202_)
  );
  INV_X1 _40597_ (
    .A(_06202_),
    .ZN(_06203_)
  );
  AND2_X1 _40598_ (
    .A1(_00007_[3]),
    .A2(_06186_),
    .ZN(_06204_)
  );
  AND2_X1 _40599_ (
    .A1(_06203_),
    .A2(_06204_),
    .ZN(_06205_)
  );
  INV_X1 _40600_ (
    .A(_06205_),
    .ZN(_06206_)
  );
  AND2_X1 _40601_ (
    .A1(_21786_),
    .A2(_00007_[2]),
    .ZN(_06207_)
  );
  INV_X1 _40602_ (
    .A(_06207_),
    .ZN(_06208_)
  );
  AND2_X1 _40603_ (
    .A1(_21494_),
    .A2(_22077_),
    .ZN(_06209_)
  );
  INV_X1 _40604_ (
    .A(_06209_),
    .ZN(_06210_)
  );
  AND2_X1 _40605_ (
    .A1(_00007_[0]),
    .A2(_06210_),
    .ZN(_06211_)
  );
  AND2_X1 _40606_ (
    .A1(_06208_),
    .A2(_06211_),
    .ZN(_06212_)
  );
  INV_X1 _40607_ (
    .A(_06212_),
    .ZN(_06213_)
  );
  AND2_X1 _40608_ (
    .A1(_21811_),
    .A2(_00007_[2]),
    .ZN(_06214_)
  );
  INV_X1 _40609_ (
    .A(_06214_),
    .ZN(_06215_)
  );
  AND2_X1 _40610_ (
    .A1(_21544_),
    .A2(_22077_),
    .ZN(_06216_)
  );
  INV_X1 _40611_ (
    .A(_06216_),
    .ZN(_06217_)
  );
  AND2_X1 _40612_ (
    .A1(_22152_),
    .A2(_06217_),
    .ZN(_06218_)
  );
  AND2_X1 _40613_ (
    .A1(_06215_),
    .A2(_06218_),
    .ZN(_06219_)
  );
  INV_X1 _40614_ (
    .A(_06219_),
    .ZN(_06220_)
  );
  AND2_X1 _40615_ (
    .A1(_06213_),
    .A2(_06220_),
    .ZN(_06221_)
  );
  AND2_X1 _40616_ (
    .A1(_00007_[1]),
    .A2(_06221_),
    .ZN(_06222_)
  );
  INV_X1 _40617_ (
    .A(_06222_),
    .ZN(_06223_)
  );
  AND2_X1 _40618_ (
    .A1(_21739_),
    .A2(_00007_[2]),
    .ZN(_06224_)
  );
  INV_X1 _40619_ (
    .A(_06224_),
    .ZN(_06225_)
  );
  AND2_X1 _40620_ (
    .A1(_21519_),
    .A2(_22077_),
    .ZN(_06226_)
  );
  INV_X1 _40621_ (
    .A(_06226_),
    .ZN(_06227_)
  );
  AND2_X1 _40622_ (
    .A1(_00007_[0]),
    .A2(_06227_),
    .ZN(_06228_)
  );
  AND2_X1 _40623_ (
    .A1(_06225_),
    .A2(_06228_),
    .ZN(_06229_)
  );
  INV_X1 _40624_ (
    .A(_06229_),
    .ZN(_06230_)
  );
  AND2_X1 _40625_ (
    .A1(_21960_),
    .A2(_22077_),
    .ZN(_06231_)
  );
  INV_X1 _40626_ (
    .A(_06231_),
    .ZN(_06232_)
  );
  AND2_X1 _40627_ (
    .A1(_21676_),
    .A2(_00007_[2]),
    .ZN(_06233_)
  );
  INV_X1 _40628_ (
    .A(_06233_),
    .ZN(_06234_)
  );
  AND2_X1 _40629_ (
    .A1(_06232_),
    .A2(_06234_),
    .ZN(_06235_)
  );
  AND2_X1 _40630_ (
    .A1(_22152_),
    .A2(_06235_),
    .ZN(_06236_)
  );
  INV_X1 _40631_ (
    .A(_06236_),
    .ZN(_06237_)
  );
  AND2_X1 _40632_ (
    .A1(_06230_),
    .A2(_06237_),
    .ZN(_06238_)
  );
  AND2_X1 _40633_ (
    .A1(_22078_),
    .A2(_06238_),
    .ZN(_06239_)
  );
  INV_X1 _40634_ (
    .A(_06239_),
    .ZN(_06240_)
  );
  AND2_X1 _40635_ (
    .A1(_06223_),
    .A2(_06240_),
    .ZN(_06241_)
  );
  AND2_X1 _40636_ (
    .A1(_22109_),
    .A2(_06241_),
    .ZN(_06242_)
  );
  INV_X1 _40637_ (
    .A(_06242_),
    .ZN(_06243_)
  );
  AND2_X1 _40638_ (
    .A1(_06206_),
    .A2(_06243_),
    .ZN(_06244_)
  );
  AND2_X1 _40639_ (
    .A1(_21894_),
    .A2(_00007_[2]),
    .ZN(_06245_)
  );
  INV_X1 _40640_ (
    .A(_06245_),
    .ZN(_06246_)
  );
  AND2_X1 _40641_ (
    .A1(_21838_),
    .A2(_22077_),
    .ZN(_06247_)
  );
  INV_X1 _40642_ (
    .A(_06247_),
    .ZN(_06248_)
  );
  AND2_X1 _40643_ (
    .A1(_00007_[0]),
    .A2(_06248_),
    .ZN(_06249_)
  );
  AND2_X1 _40644_ (
    .A1(_06246_),
    .A2(_06249_),
    .ZN(_06250_)
  );
  INV_X1 _40645_ (
    .A(_06250_),
    .ZN(_06251_)
  );
  AND2_X1 _40646_ (
    .A1(_21572_),
    .A2(_22077_),
    .ZN(_06252_)
  );
  INV_X1 _40647_ (
    .A(_06252_),
    .ZN(_06253_)
  );
  AND2_X1 _40648_ (
    .A1(_21910_),
    .A2(_00007_[2]),
    .ZN(_06254_)
  );
  INV_X1 _40649_ (
    .A(_06254_),
    .ZN(_06255_)
  );
  AND2_X1 _40650_ (
    .A1(_06253_),
    .A2(_06255_),
    .ZN(_06256_)
  );
  AND2_X1 _40651_ (
    .A1(_22152_),
    .A2(_06256_),
    .ZN(_06257_)
  );
  INV_X1 _40652_ (
    .A(_06257_),
    .ZN(_06258_)
  );
  AND2_X1 _40653_ (
    .A1(_06251_),
    .A2(_06258_),
    .ZN(_06259_)
  );
  AND2_X1 _40654_ (
    .A1(_22078_),
    .A2(_06259_),
    .ZN(_06260_)
  );
  INV_X1 _40655_ (
    .A(_06260_),
    .ZN(_06261_)
  );
  AND2_X1 _40656_ (
    .A1(_21870_),
    .A2(_22077_),
    .ZN(_06262_)
  );
  INV_X1 _40657_ (
    .A(_06262_),
    .ZN(_06263_)
  );
  AND2_X1 _40658_ (
    .A1(_21854_),
    .A2(_00007_[2]),
    .ZN(_06264_)
  );
  INV_X1 _40659_ (
    .A(_06264_),
    .ZN(_06265_)
  );
  AND2_X1 _40660_ (
    .A1(_06263_),
    .A2(_06265_),
    .ZN(_06266_)
  );
  AND2_X1 _40661_ (
    .A1(_22152_),
    .A2(_06266_),
    .ZN(_06267_)
  );
  INV_X1 _40662_ (
    .A(_06267_),
    .ZN(_06268_)
  );
  AND2_X1 _40663_ (
    .A1(_21942_),
    .A2(_00007_[2]),
    .ZN(_06269_)
  );
  INV_X1 _40664_ (
    .A(_06269_),
    .ZN(_06270_)
  );
  AND2_X1 _40665_ (
    .A1(_21926_),
    .A2(_22077_),
    .ZN(_06271_)
  );
  INV_X1 _40666_ (
    .A(_06271_),
    .ZN(_06272_)
  );
  AND2_X1 _40667_ (
    .A1(_00007_[0]),
    .A2(_06272_),
    .ZN(_06273_)
  );
  AND2_X1 _40668_ (
    .A1(_06270_),
    .A2(_06273_),
    .ZN(_06274_)
  );
  INV_X1 _40669_ (
    .A(_06274_),
    .ZN(_06275_)
  );
  AND2_X1 _40670_ (
    .A1(_06268_),
    .A2(_06275_),
    .ZN(_06276_)
  );
  AND2_X1 _40671_ (
    .A1(_00007_[1]),
    .A2(_06276_),
    .ZN(_06277_)
  );
  INV_X1 _40672_ (
    .A(_06277_),
    .ZN(_06278_)
  );
  AND2_X1 _40673_ (
    .A1(_00007_[3]),
    .A2(_06261_),
    .ZN(_06279_)
  );
  AND2_X1 _40674_ (
    .A1(_06278_),
    .A2(_06279_),
    .ZN(_06280_)
  );
  INV_X1 _40675_ (
    .A(_06280_),
    .ZN(_06281_)
  );
  AND2_X1 _40676_ (
    .A1(_21596_),
    .A2(_22077_),
    .ZN(_06282_)
  );
  INV_X1 _40677_ (
    .A(_06282_),
    .ZN(_06283_)
  );
  AND2_X1 _40678_ (
    .A1(_21415_),
    .A2(_00007_[2]),
    .ZN(_06284_)
  );
  INV_X1 _40679_ (
    .A(_06284_),
    .ZN(_06285_)
  );
  AND2_X1 _40680_ (
    .A1(_21442_),
    .A2(_22077_),
    .ZN(_06286_)
  );
  INV_X1 _40681_ (
    .A(_06286_),
    .ZN(_06287_)
  );
  AND2_X1 _40682_ (
    .A1(_21653_),
    .A2(_00007_[2]),
    .ZN(_06288_)
  );
  INV_X1 _40683_ (
    .A(_06288_),
    .ZN(_06289_)
  );
  AND2_X1 _40684_ (
    .A1(_06287_),
    .A2(_06289_),
    .ZN(_06290_)
  );
  AND2_X1 _40685_ (
    .A1(_21376_),
    .A2(_00007_[2]),
    .ZN(_06291_)
  );
  INV_X1 _40686_ (
    .A(_06291_),
    .ZN(_06292_)
  );
  AND2_X1 _40687_ (
    .A1(_21622_),
    .A2(_22077_),
    .ZN(_06293_)
  );
  INV_X1 _40688_ (
    .A(_06293_),
    .ZN(_06294_)
  );
  AND2_X1 _40689_ (
    .A1(_21464_),
    .A2(_22077_),
    .ZN(_06295_)
  );
  INV_X1 _40690_ (
    .A(_06295_),
    .ZN(_06296_)
  );
  AND2_X1 _40691_ (
    .A1(_21763_),
    .A2(_00007_[2]),
    .ZN(_06297_)
  );
  INV_X1 _40692_ (
    .A(_06297_),
    .ZN(_06298_)
  );
  AND2_X1 _40693_ (
    .A1(_00007_[0]),
    .A2(_06294_),
    .ZN(_06299_)
  );
  AND2_X1 _40694_ (
    .A1(_06292_),
    .A2(_06299_),
    .ZN(_06300_)
  );
  INV_X1 _40695_ (
    .A(_06300_),
    .ZN(_06301_)
  );
  AND2_X1 _40696_ (
    .A1(_22152_),
    .A2(_06283_),
    .ZN(_06302_)
  );
  AND2_X1 _40697_ (
    .A1(_06285_),
    .A2(_06302_),
    .ZN(_06303_)
  );
  INV_X1 _40698_ (
    .A(_06303_),
    .ZN(_06304_)
  );
  AND2_X1 _40699_ (
    .A1(_06301_),
    .A2(_06304_),
    .ZN(_06305_)
  );
  AND2_X1 _40700_ (
    .A1(_00007_[1]),
    .A2(_06305_),
    .ZN(_06306_)
  );
  INV_X1 _40701_ (
    .A(_06306_),
    .ZN(_06307_)
  );
  AND2_X1 _40702_ (
    .A1(_00007_[0]),
    .A2(_06296_),
    .ZN(_06308_)
  );
  AND2_X1 _40703_ (
    .A1(_06298_),
    .A2(_06308_),
    .ZN(_06309_)
  );
  INV_X1 _40704_ (
    .A(_06309_),
    .ZN(_06310_)
  );
  AND2_X1 _40705_ (
    .A1(_22152_),
    .A2(_06290_),
    .ZN(_06311_)
  );
  INV_X1 _40706_ (
    .A(_06311_),
    .ZN(_06312_)
  );
  AND2_X1 _40707_ (
    .A1(_06310_),
    .A2(_06312_),
    .ZN(_06313_)
  );
  AND2_X1 _40708_ (
    .A1(_22078_),
    .A2(_06313_),
    .ZN(_06314_)
  );
  INV_X1 _40709_ (
    .A(_06314_),
    .ZN(_06315_)
  );
  AND2_X1 _40710_ (
    .A1(_06307_),
    .A2(_06315_),
    .ZN(_06316_)
  );
  AND2_X1 _40711_ (
    .A1(_22109_),
    .A2(_06316_),
    .ZN(_06317_)
  );
  INV_X1 _40712_ (
    .A(_06317_),
    .ZN(_06318_)
  );
  AND2_X1 _40713_ (
    .A1(_06281_),
    .A2(_06318_),
    .ZN(_06319_)
  );
  AND2_X1 _40714_ (
    .A1(_22144_),
    .A2(_06244_),
    .ZN(_06320_)
  );
  INV_X1 _40715_ (
    .A(_06320_),
    .ZN(_06321_)
  );
  AND2_X1 _40716_ (
    .A1(_00007_[4]),
    .A2(_06319_),
    .ZN(_06322_)
  );
  INV_X1 _40717_ (
    .A(_06322_),
    .ZN(_06323_)
  );
  AND2_X1 _40718_ (
    .A1(_06321_),
    .A2(_06323_),
    .ZN(_06324_)
  );
  AND2_X1 _40719_ (
    .A1(_05842_),
    .A2(_06324_),
    .ZN(_06325_)
  );
  INV_X1 _40720_ (
    .A(_06325_),
    .ZN(_06326_)
  );
  AND2_X1 _40721_ (
    .A1(decoded_imm[7]),
    .A2(_04966_),
    .ZN(_06327_)
  );
  INV_X1 _40722_ (
    .A(_06327_),
    .ZN(_06328_)
  );
  AND2_X1 _40723_ (
    .A1(_04962_),
    .A2(_06328_),
    .ZN(_06329_)
  );
  AND2_X1 _40724_ (
    .A1(_06326_),
    .A2(_06329_),
    .ZN(_06330_)
  );
  INV_X1 _40725_ (
    .A(_06330_),
    .ZN(_06331_)
  );
  AND2_X1 _40726_ (
    .A1(_21207_),
    .A2(_04963_),
    .ZN(_06332_)
  );
  INV_X1 _40727_ (
    .A(_06332_),
    .ZN(_06333_)
  );
  AND2_X1 _40728_ (
    .A1(_06331_),
    .A2(_06333_),
    .ZN(_00288_)
  );
  AND2_X1 _40729_ (
    .A1(decoded_imm[8]),
    .A2(_04966_),
    .ZN(_06334_)
  );
  INV_X1 _40730_ (
    .A(_06334_),
    .ZN(_06335_)
  );
  AND2_X1 _40731_ (
    .A1(\cpuregs[28] [8]),
    .A2(_00007_[2]),
    .ZN(_06336_)
  );
  INV_X1 _40732_ (
    .A(_06336_),
    .ZN(_06337_)
  );
  AND2_X1 _40733_ (
    .A1(\cpuregs[24] [8]),
    .A2(_22077_),
    .ZN(_06338_)
  );
  INV_X1 _40734_ (
    .A(_06338_),
    .ZN(_06339_)
  );
  AND2_X1 _40735_ (
    .A1(_22152_),
    .A2(_06339_),
    .ZN(_06340_)
  );
  AND2_X1 _40736_ (
    .A1(_06337_),
    .A2(_06340_),
    .ZN(_06341_)
  );
  INV_X1 _40737_ (
    .A(_06341_),
    .ZN(_06342_)
  );
  AND2_X1 _40738_ (
    .A1(\cpuregs[29] [8]),
    .A2(_00007_[2]),
    .ZN(_06343_)
  );
  INV_X1 _40739_ (
    .A(_06343_),
    .ZN(_06344_)
  );
  AND2_X1 _40740_ (
    .A1(\cpuregs[25] [8]),
    .A2(_22077_),
    .ZN(_06345_)
  );
  INV_X1 _40741_ (
    .A(_06345_),
    .ZN(_06346_)
  );
  AND2_X1 _40742_ (
    .A1(_00007_[0]),
    .A2(_06346_),
    .ZN(_06347_)
  );
  AND2_X1 _40743_ (
    .A1(_06344_),
    .A2(_06347_),
    .ZN(_06348_)
  );
  INV_X1 _40744_ (
    .A(_06348_),
    .ZN(_06349_)
  );
  AND2_X1 _40745_ (
    .A1(_06342_),
    .A2(_06349_),
    .ZN(_06350_)
  );
  INV_X1 _40746_ (
    .A(_06350_),
    .ZN(_06351_)
  );
  AND2_X1 _40747_ (
    .A1(_22078_),
    .A2(_06351_),
    .ZN(_06352_)
  );
  INV_X1 _40748_ (
    .A(_06352_),
    .ZN(_06353_)
  );
  AND2_X1 _40749_ (
    .A1(\cpuregs[26] [8]),
    .A2(_22077_),
    .ZN(_06354_)
  );
  INV_X1 _40750_ (
    .A(_06354_),
    .ZN(_06355_)
  );
  AND2_X1 _40751_ (
    .A1(\cpuregs[30] [8]),
    .A2(_00007_[2]),
    .ZN(_06356_)
  );
  INV_X1 _40752_ (
    .A(_06356_),
    .ZN(_06357_)
  );
  AND2_X1 _40753_ (
    .A1(_22152_),
    .A2(_06357_),
    .ZN(_06358_)
  );
  AND2_X1 _40754_ (
    .A1(_06355_),
    .A2(_06358_),
    .ZN(_06359_)
  );
  INV_X1 _40755_ (
    .A(_06359_),
    .ZN(_06360_)
  );
  AND2_X1 _40756_ (
    .A1(\cpuregs[27] [8]),
    .A2(_22077_),
    .ZN(_06361_)
  );
  INV_X1 _40757_ (
    .A(_06361_),
    .ZN(_06362_)
  );
  AND2_X1 _40758_ (
    .A1(\cpuregs[31] [8]),
    .A2(_00007_[2]),
    .ZN(_06363_)
  );
  INV_X1 _40759_ (
    .A(_06363_),
    .ZN(_06364_)
  );
  AND2_X1 _40760_ (
    .A1(_00007_[0]),
    .A2(_06364_),
    .ZN(_06365_)
  );
  AND2_X1 _40761_ (
    .A1(_06362_),
    .A2(_06365_),
    .ZN(_06366_)
  );
  INV_X1 _40762_ (
    .A(_06366_),
    .ZN(_06367_)
  );
  AND2_X1 _40763_ (
    .A1(_06360_),
    .A2(_06367_),
    .ZN(_06368_)
  );
  INV_X1 _40764_ (
    .A(_06368_),
    .ZN(_06369_)
  );
  AND2_X1 _40765_ (
    .A1(_00007_[1]),
    .A2(_06369_),
    .ZN(_06370_)
  );
  INV_X1 _40766_ (
    .A(_06370_),
    .ZN(_06371_)
  );
  AND2_X1 _40767_ (
    .A1(_00007_[3]),
    .A2(_06371_),
    .ZN(_06372_)
  );
  AND2_X1 _40768_ (
    .A1(_06353_),
    .A2(_06372_),
    .ZN(_06373_)
  );
  INV_X1 _40769_ (
    .A(_06373_),
    .ZN(_06374_)
  );
  AND2_X1 _40770_ (
    .A1(\cpuregs[19] [8]),
    .A2(_00007_[1]),
    .ZN(_06375_)
  );
  INV_X1 _40771_ (
    .A(_06375_),
    .ZN(_06376_)
  );
  AND2_X1 _40772_ (
    .A1(\cpuregs[17] [8]),
    .A2(_22078_),
    .ZN(_06377_)
  );
  INV_X1 _40773_ (
    .A(_06377_),
    .ZN(_06378_)
  );
  AND2_X1 _40774_ (
    .A1(_06376_),
    .A2(_06378_),
    .ZN(_06379_)
  );
  INV_X1 _40775_ (
    .A(_06379_),
    .ZN(_06380_)
  );
  AND2_X1 _40776_ (
    .A1(_22077_),
    .A2(_06380_),
    .ZN(_06381_)
  );
  INV_X1 _40777_ (
    .A(_06381_),
    .ZN(_06382_)
  );
  AND2_X1 _40778_ (
    .A1(\cpuregs[23] [8]),
    .A2(_00007_[1]),
    .ZN(_06383_)
  );
  INV_X1 _40779_ (
    .A(_06383_),
    .ZN(_06384_)
  );
  AND2_X1 _40780_ (
    .A1(\cpuregs[21] [8]),
    .A2(_22078_),
    .ZN(_06385_)
  );
  INV_X1 _40781_ (
    .A(_06385_),
    .ZN(_06386_)
  );
  AND2_X1 _40782_ (
    .A1(_06384_),
    .A2(_06386_),
    .ZN(_06387_)
  );
  INV_X1 _40783_ (
    .A(_06387_),
    .ZN(_06388_)
  );
  AND2_X1 _40784_ (
    .A1(_00007_[2]),
    .A2(_06388_),
    .ZN(_06389_)
  );
  INV_X1 _40785_ (
    .A(_06389_),
    .ZN(_06390_)
  );
  AND2_X1 _40786_ (
    .A1(_00007_[0]),
    .A2(_06390_),
    .ZN(_06391_)
  );
  AND2_X1 _40787_ (
    .A1(_06382_),
    .A2(_06391_),
    .ZN(_06392_)
  );
  INV_X1 _40788_ (
    .A(_06392_),
    .ZN(_06393_)
  );
  AND2_X1 _40789_ (
    .A1(\cpuregs[18] [8]),
    .A2(_00007_[1]),
    .ZN(_06394_)
  );
  INV_X1 _40790_ (
    .A(_06394_),
    .ZN(_06395_)
  );
  AND2_X1 _40791_ (
    .A1(\cpuregs[16] [8]),
    .A2(_22078_),
    .ZN(_06396_)
  );
  INV_X1 _40792_ (
    .A(_06396_),
    .ZN(_06397_)
  );
  AND2_X1 _40793_ (
    .A1(_06395_),
    .A2(_06397_),
    .ZN(_06398_)
  );
  INV_X1 _40794_ (
    .A(_06398_),
    .ZN(_06399_)
  );
  AND2_X1 _40795_ (
    .A1(_22077_),
    .A2(_06399_),
    .ZN(_06400_)
  );
  INV_X1 _40796_ (
    .A(_06400_),
    .ZN(_06401_)
  );
  AND2_X1 _40797_ (
    .A1(\cpuregs[22] [8]),
    .A2(_00007_[1]),
    .ZN(_06402_)
  );
  INV_X1 _40798_ (
    .A(_06402_),
    .ZN(_06403_)
  );
  AND2_X1 _40799_ (
    .A1(\cpuregs[20] [8]),
    .A2(_22078_),
    .ZN(_06404_)
  );
  INV_X1 _40800_ (
    .A(_06404_),
    .ZN(_06405_)
  );
  AND2_X1 _40801_ (
    .A1(_06403_),
    .A2(_06405_),
    .ZN(_06406_)
  );
  INV_X1 _40802_ (
    .A(_06406_),
    .ZN(_06407_)
  );
  AND2_X1 _40803_ (
    .A1(_00007_[2]),
    .A2(_06407_),
    .ZN(_06408_)
  );
  INV_X1 _40804_ (
    .A(_06408_),
    .ZN(_06409_)
  );
  AND2_X1 _40805_ (
    .A1(_22152_),
    .A2(_06409_),
    .ZN(_06410_)
  );
  AND2_X1 _40806_ (
    .A1(_06401_),
    .A2(_06410_),
    .ZN(_06411_)
  );
  INV_X1 _40807_ (
    .A(_06411_),
    .ZN(_06412_)
  );
  AND2_X1 _40808_ (
    .A1(_22109_),
    .A2(_06412_),
    .ZN(_06413_)
  );
  AND2_X1 _40809_ (
    .A1(_06393_),
    .A2(_06413_),
    .ZN(_06414_)
  );
  INV_X1 _40810_ (
    .A(_06414_),
    .ZN(_06415_)
  );
  AND2_X1 _40811_ (
    .A1(_06374_),
    .A2(_06415_),
    .ZN(_06416_)
  );
  AND2_X1 _40812_ (
    .A1(\cpuregs[8] [8]),
    .A2(_22078_),
    .ZN(_06417_)
  );
  INV_X1 _40813_ (
    .A(_06417_),
    .ZN(_06418_)
  );
  AND2_X1 _40814_ (
    .A1(\cpuregs[10] [8]),
    .A2(_00007_[1]),
    .ZN(_06419_)
  );
  INV_X1 _40815_ (
    .A(_06419_),
    .ZN(_06420_)
  );
  AND2_X1 _40816_ (
    .A1(_22077_),
    .A2(_06420_),
    .ZN(_06421_)
  );
  AND2_X1 _40817_ (
    .A1(_06418_),
    .A2(_06421_),
    .ZN(_06422_)
  );
  INV_X1 _40818_ (
    .A(_06422_),
    .ZN(_06423_)
  );
  AND2_X1 _40819_ (
    .A1(\cpuregs[12] [8]),
    .A2(_22078_),
    .ZN(_06424_)
  );
  INV_X1 _40820_ (
    .A(_06424_),
    .ZN(_06425_)
  );
  AND2_X1 _40821_ (
    .A1(\cpuregs[14] [8]),
    .A2(_00007_[1]),
    .ZN(_06426_)
  );
  INV_X1 _40822_ (
    .A(_06426_),
    .ZN(_06427_)
  );
  AND2_X1 _40823_ (
    .A1(_00007_[2]),
    .A2(_06427_),
    .ZN(_06428_)
  );
  AND2_X1 _40824_ (
    .A1(_06425_),
    .A2(_06428_),
    .ZN(_06429_)
  );
  INV_X1 _40825_ (
    .A(_06429_),
    .ZN(_06430_)
  );
  AND2_X1 _40826_ (
    .A1(_06423_),
    .A2(_06430_),
    .ZN(_06431_)
  );
  INV_X1 _40827_ (
    .A(_06431_),
    .ZN(_06432_)
  );
  AND2_X1 _40828_ (
    .A1(_22152_),
    .A2(_06432_),
    .ZN(_06433_)
  );
  INV_X1 _40829_ (
    .A(_06433_),
    .ZN(_06434_)
  );
  AND2_X1 _40830_ (
    .A1(\cpuregs[9] [8]),
    .A2(_22078_),
    .ZN(_06435_)
  );
  INV_X1 _40831_ (
    .A(_06435_),
    .ZN(_06436_)
  );
  AND2_X1 _40832_ (
    .A1(\cpuregs[11] [8]),
    .A2(_00007_[1]),
    .ZN(_06437_)
  );
  INV_X1 _40833_ (
    .A(_06437_),
    .ZN(_06438_)
  );
  AND2_X1 _40834_ (
    .A1(_22077_),
    .A2(_06438_),
    .ZN(_06439_)
  );
  AND2_X1 _40835_ (
    .A1(_06436_),
    .A2(_06439_),
    .ZN(_06440_)
  );
  INV_X1 _40836_ (
    .A(_06440_),
    .ZN(_06441_)
  );
  AND2_X1 _40837_ (
    .A1(\cpuregs[13] [8]),
    .A2(_22078_),
    .ZN(_06442_)
  );
  INV_X1 _40838_ (
    .A(_06442_),
    .ZN(_06443_)
  );
  AND2_X1 _40839_ (
    .A1(\cpuregs[15] [8]),
    .A2(_00007_[1]),
    .ZN(_06444_)
  );
  INV_X1 _40840_ (
    .A(_06444_),
    .ZN(_06445_)
  );
  AND2_X1 _40841_ (
    .A1(_00007_[2]),
    .A2(_06445_),
    .ZN(_06446_)
  );
  AND2_X1 _40842_ (
    .A1(_06443_),
    .A2(_06446_),
    .ZN(_06447_)
  );
  INV_X1 _40843_ (
    .A(_06447_),
    .ZN(_06448_)
  );
  AND2_X1 _40844_ (
    .A1(_06441_),
    .A2(_06448_),
    .ZN(_06449_)
  );
  INV_X1 _40845_ (
    .A(_06449_),
    .ZN(_06450_)
  );
  AND2_X1 _40846_ (
    .A1(_00007_[0]),
    .A2(_06450_),
    .ZN(_06451_)
  );
  INV_X1 _40847_ (
    .A(_06451_),
    .ZN(_06452_)
  );
  AND2_X1 _40848_ (
    .A1(_00007_[3]),
    .A2(_06452_),
    .ZN(_06453_)
  );
  AND2_X1 _40849_ (
    .A1(_06434_),
    .A2(_06453_),
    .ZN(_06454_)
  );
  INV_X1 _40850_ (
    .A(_06454_),
    .ZN(_06455_)
  );
  AND2_X1 _40851_ (
    .A1(_21520_),
    .A2(_22077_),
    .ZN(_06456_)
  );
  INV_X1 _40852_ (
    .A(_06456_),
    .ZN(_06457_)
  );
  AND2_X1 _40853_ (
    .A1(_21740_),
    .A2(_00007_[2]),
    .ZN(_06458_)
  );
  INV_X1 _40854_ (
    .A(_06458_),
    .ZN(_06459_)
  );
  AND2_X1 _40855_ (
    .A1(_21961_),
    .A2(_22077_),
    .ZN(_06460_)
  );
  INV_X1 _40856_ (
    .A(_06460_),
    .ZN(_06461_)
  );
  AND2_X1 _40857_ (
    .A1(_21677_),
    .A2(_00007_[2]),
    .ZN(_06462_)
  );
  INV_X1 _40858_ (
    .A(_06462_),
    .ZN(_06463_)
  );
  AND2_X1 _40859_ (
    .A1(_06461_),
    .A2(_06463_),
    .ZN(_06464_)
  );
  AND2_X1 _40860_ (
    .A1(_00007_[0]),
    .A2(_06457_),
    .ZN(_06465_)
  );
  AND2_X1 _40861_ (
    .A1(_06459_),
    .A2(_06465_),
    .ZN(_06466_)
  );
  INV_X1 _40862_ (
    .A(_06466_),
    .ZN(_06467_)
  );
  AND2_X1 _40863_ (
    .A1(_22152_),
    .A2(_06464_),
    .ZN(_06468_)
  );
  INV_X1 _40864_ (
    .A(_06468_),
    .ZN(_06469_)
  );
  AND2_X1 _40865_ (
    .A1(_06467_),
    .A2(_06469_),
    .ZN(_06470_)
  );
  AND2_X1 _40866_ (
    .A1(_22078_),
    .A2(_06470_),
    .ZN(_06471_)
  );
  INV_X1 _40867_ (
    .A(_06471_),
    .ZN(_06472_)
  );
  AND2_X1 _40868_ (
    .A1(_21787_),
    .A2(_00007_[2]),
    .ZN(_06473_)
  );
  INV_X1 _40869_ (
    .A(_06473_),
    .ZN(_06474_)
  );
  AND2_X1 _40870_ (
    .A1(_21495_),
    .A2(_22077_),
    .ZN(_06475_)
  );
  INV_X1 _40871_ (
    .A(_06475_),
    .ZN(_06476_)
  );
  AND2_X1 _40872_ (
    .A1(_21545_),
    .A2(_22077_),
    .ZN(_06477_)
  );
  INV_X1 _40873_ (
    .A(_06477_),
    .ZN(_06478_)
  );
  AND2_X1 _40874_ (
    .A1(_21812_),
    .A2(_00007_[2]),
    .ZN(_06479_)
  );
  INV_X1 _40875_ (
    .A(_06479_),
    .ZN(_06480_)
  );
  AND2_X1 _40876_ (
    .A1(_00007_[0]),
    .A2(_06476_),
    .ZN(_06481_)
  );
  AND2_X1 _40877_ (
    .A1(_06474_),
    .A2(_06481_),
    .ZN(_06482_)
  );
  INV_X1 _40878_ (
    .A(_06482_),
    .ZN(_06483_)
  );
  AND2_X1 _40879_ (
    .A1(_22152_),
    .A2(_06478_),
    .ZN(_06484_)
  );
  AND2_X1 _40880_ (
    .A1(_06480_),
    .A2(_06484_),
    .ZN(_06485_)
  );
  INV_X1 _40881_ (
    .A(_06485_),
    .ZN(_06486_)
  );
  AND2_X1 _40882_ (
    .A1(_06483_),
    .A2(_06486_),
    .ZN(_06487_)
  );
  AND2_X1 _40883_ (
    .A1(_00007_[1]),
    .A2(_06487_),
    .ZN(_06488_)
  );
  INV_X1 _40884_ (
    .A(_06488_),
    .ZN(_06489_)
  );
  AND2_X1 _40885_ (
    .A1(_06472_),
    .A2(_06489_),
    .ZN(_06490_)
  );
  AND2_X1 _40886_ (
    .A1(_22109_),
    .A2(_06490_),
    .ZN(_06491_)
  );
  INV_X1 _40887_ (
    .A(_06491_),
    .ZN(_06492_)
  );
  AND2_X1 _40888_ (
    .A1(_06455_),
    .A2(_06492_),
    .ZN(_06493_)
  );
  AND2_X1 _40889_ (
    .A1(_22144_),
    .A2(_06493_),
    .ZN(_06494_)
  );
  INV_X1 _40890_ (
    .A(_06494_),
    .ZN(_06495_)
  );
  AND2_X1 _40891_ (
    .A1(_00007_[4]),
    .A2(_06416_),
    .ZN(_06496_)
  );
  INV_X1 _40892_ (
    .A(_06496_),
    .ZN(_06497_)
  );
  AND2_X1 _40893_ (
    .A1(_21208_),
    .A2(_04963_),
    .ZN(_06498_)
  );
  INV_X1 _40894_ (
    .A(_06498_),
    .ZN(_06499_)
  );
  AND2_X1 _40895_ (
    .A1(_05842_),
    .A2(_06497_),
    .ZN(_06500_)
  );
  AND2_X1 _40896_ (
    .A1(_06495_),
    .A2(_06500_),
    .ZN(_06501_)
  );
  INV_X1 _40897_ (
    .A(_06501_),
    .ZN(_06502_)
  );
  AND2_X1 _40898_ (
    .A1(_04962_),
    .A2(_06335_),
    .ZN(_06503_)
  );
  AND2_X1 _40899_ (
    .A1(_06502_),
    .A2(_06503_),
    .ZN(_06504_)
  );
  INV_X1 _40900_ (
    .A(_06504_),
    .ZN(_06505_)
  );
  AND2_X1 _40901_ (
    .A1(_06499_),
    .A2(_06505_),
    .ZN(_00289_)
  );
  AND2_X1 _40902_ (
    .A1(decoded_imm[9]),
    .A2(_04966_),
    .ZN(_06506_)
  );
  INV_X1 _40903_ (
    .A(_06506_),
    .ZN(_06507_)
  );
  AND2_X1 _40904_ (
    .A1(\cpuregs[9] [9]),
    .A2(_22077_),
    .ZN(_06508_)
  );
  INV_X1 _40905_ (
    .A(_06508_),
    .ZN(_06509_)
  );
  AND2_X1 _40906_ (
    .A1(\cpuregs[13] [9]),
    .A2(_00007_[2]),
    .ZN(_06510_)
  );
  INV_X1 _40907_ (
    .A(_06510_),
    .ZN(_06511_)
  );
  AND2_X1 _40908_ (
    .A1(_00007_[0]),
    .A2(_06511_),
    .ZN(_06512_)
  );
  AND2_X1 _40909_ (
    .A1(_06509_),
    .A2(_06512_),
    .ZN(_06513_)
  );
  INV_X1 _40910_ (
    .A(_06513_),
    .ZN(_06514_)
  );
  AND2_X1 _40911_ (
    .A1(\cpuregs[8] [9]),
    .A2(_22077_),
    .ZN(_06515_)
  );
  INV_X1 _40912_ (
    .A(_06515_),
    .ZN(_06516_)
  );
  AND2_X1 _40913_ (
    .A1(\cpuregs[12] [9]),
    .A2(_00007_[2]),
    .ZN(_06517_)
  );
  INV_X1 _40914_ (
    .A(_06517_),
    .ZN(_06518_)
  );
  AND2_X1 _40915_ (
    .A1(_22152_),
    .A2(_06518_),
    .ZN(_06519_)
  );
  AND2_X1 _40916_ (
    .A1(_06516_),
    .A2(_06519_),
    .ZN(_06520_)
  );
  INV_X1 _40917_ (
    .A(_06520_),
    .ZN(_06521_)
  );
  AND2_X1 _40918_ (
    .A1(_22078_),
    .A2(_06521_),
    .ZN(_06522_)
  );
  AND2_X1 _40919_ (
    .A1(_06514_),
    .A2(_06522_),
    .ZN(_06523_)
  );
  INV_X1 _40920_ (
    .A(_06523_),
    .ZN(_06524_)
  );
  AND2_X1 _40921_ (
    .A1(\cpuregs[15] [9]),
    .A2(_00007_[2]),
    .ZN(_06525_)
  );
  INV_X1 _40922_ (
    .A(_06525_),
    .ZN(_06526_)
  );
  AND2_X1 _40923_ (
    .A1(\cpuregs[11] [9]),
    .A2(_22077_),
    .ZN(_06527_)
  );
  INV_X1 _40924_ (
    .A(_06527_),
    .ZN(_06528_)
  );
  AND2_X1 _40925_ (
    .A1(_00007_[0]),
    .A2(_06528_),
    .ZN(_06529_)
  );
  AND2_X1 _40926_ (
    .A1(_06526_),
    .A2(_06529_),
    .ZN(_06530_)
  );
  INV_X1 _40927_ (
    .A(_06530_),
    .ZN(_06531_)
  );
  AND2_X1 _40928_ (
    .A1(\cpuregs[14] [9]),
    .A2(_00007_[2]),
    .ZN(_06532_)
  );
  INV_X1 _40929_ (
    .A(_06532_),
    .ZN(_06533_)
  );
  AND2_X1 _40930_ (
    .A1(\cpuregs[10] [9]),
    .A2(_22077_),
    .ZN(_06534_)
  );
  INV_X1 _40931_ (
    .A(_06534_),
    .ZN(_06535_)
  );
  AND2_X1 _40932_ (
    .A1(_22152_),
    .A2(_06535_),
    .ZN(_06536_)
  );
  AND2_X1 _40933_ (
    .A1(_06533_),
    .A2(_06536_),
    .ZN(_06537_)
  );
  INV_X1 _40934_ (
    .A(_06537_),
    .ZN(_06538_)
  );
  AND2_X1 _40935_ (
    .A1(_00007_[1]),
    .A2(_06538_),
    .ZN(_06539_)
  );
  AND2_X1 _40936_ (
    .A1(_06531_),
    .A2(_06539_),
    .ZN(_06540_)
  );
  INV_X1 _40937_ (
    .A(_06540_),
    .ZN(_06541_)
  );
  AND2_X1 _40938_ (
    .A1(_06524_),
    .A2(_06541_),
    .ZN(_06542_)
  );
  INV_X1 _40939_ (
    .A(_06542_),
    .ZN(_06543_)
  );
  AND2_X1 _40940_ (
    .A1(_00007_[3]),
    .A2(_06543_),
    .ZN(_06544_)
  );
  INV_X1 _40941_ (
    .A(_06544_),
    .ZN(_06545_)
  );
  AND2_X1 _40942_ (
    .A1(\cpuregs[1] [9]),
    .A2(_22077_),
    .ZN(_06546_)
  );
  INV_X1 _40943_ (
    .A(_06546_),
    .ZN(_06547_)
  );
  AND2_X1 _40944_ (
    .A1(\cpuregs[5] [9]),
    .A2(_00007_[2]),
    .ZN(_06548_)
  );
  INV_X1 _40945_ (
    .A(_06548_),
    .ZN(_06549_)
  );
  AND2_X1 _40946_ (
    .A1(_00007_[0]),
    .A2(_06549_),
    .ZN(_06550_)
  );
  AND2_X1 _40947_ (
    .A1(_06547_),
    .A2(_06550_),
    .ZN(_06551_)
  );
  INV_X1 _40948_ (
    .A(_06551_),
    .ZN(_06552_)
  );
  AND2_X1 _40949_ (
    .A1(\cpuregs[0] [9]),
    .A2(_22077_),
    .ZN(_06553_)
  );
  INV_X1 _40950_ (
    .A(_06553_),
    .ZN(_06554_)
  );
  AND2_X1 _40951_ (
    .A1(\cpuregs[4] [9]),
    .A2(_00007_[2]),
    .ZN(_06555_)
  );
  INV_X1 _40952_ (
    .A(_06555_),
    .ZN(_06556_)
  );
  AND2_X1 _40953_ (
    .A1(_22152_),
    .A2(_06556_),
    .ZN(_06557_)
  );
  AND2_X1 _40954_ (
    .A1(_06554_),
    .A2(_06557_),
    .ZN(_06558_)
  );
  INV_X1 _40955_ (
    .A(_06558_),
    .ZN(_06559_)
  );
  AND2_X1 _40956_ (
    .A1(_22078_),
    .A2(_06559_),
    .ZN(_06560_)
  );
  AND2_X1 _40957_ (
    .A1(_06552_),
    .A2(_06560_),
    .ZN(_06561_)
  );
  INV_X1 _40958_ (
    .A(_06561_),
    .ZN(_06562_)
  );
  AND2_X1 _40959_ (
    .A1(\cpuregs[3] [9]),
    .A2(_22077_),
    .ZN(_06563_)
  );
  INV_X1 _40960_ (
    .A(_06563_),
    .ZN(_06564_)
  );
  AND2_X1 _40961_ (
    .A1(\cpuregs[7] [9]),
    .A2(_00007_[2]),
    .ZN(_06565_)
  );
  INV_X1 _40962_ (
    .A(_06565_),
    .ZN(_06566_)
  );
  AND2_X1 _40963_ (
    .A1(_00007_[0]),
    .A2(_06566_),
    .ZN(_06567_)
  );
  AND2_X1 _40964_ (
    .A1(_06564_),
    .A2(_06567_),
    .ZN(_06568_)
  );
  INV_X1 _40965_ (
    .A(_06568_),
    .ZN(_06569_)
  );
  AND2_X1 _40966_ (
    .A1(\cpuregs[6] [9]),
    .A2(_00007_[2]),
    .ZN(_06570_)
  );
  INV_X1 _40967_ (
    .A(_06570_),
    .ZN(_06571_)
  );
  AND2_X1 _40968_ (
    .A1(\cpuregs[2] [9]),
    .A2(_22077_),
    .ZN(_06572_)
  );
  INV_X1 _40969_ (
    .A(_06572_),
    .ZN(_06573_)
  );
  AND2_X1 _40970_ (
    .A1(_22152_),
    .A2(_06573_),
    .ZN(_06574_)
  );
  AND2_X1 _40971_ (
    .A1(_06571_),
    .A2(_06574_),
    .ZN(_06575_)
  );
  INV_X1 _40972_ (
    .A(_06575_),
    .ZN(_06576_)
  );
  AND2_X1 _40973_ (
    .A1(_00007_[1]),
    .A2(_06576_),
    .ZN(_06577_)
  );
  AND2_X1 _40974_ (
    .A1(_06569_),
    .A2(_06577_),
    .ZN(_06578_)
  );
  INV_X1 _40975_ (
    .A(_06578_),
    .ZN(_06579_)
  );
  AND2_X1 _40976_ (
    .A1(_06562_),
    .A2(_06579_),
    .ZN(_06580_)
  );
  INV_X1 _40977_ (
    .A(_06580_),
    .ZN(_06581_)
  );
  AND2_X1 _40978_ (
    .A1(_22109_),
    .A2(_06581_),
    .ZN(_06582_)
  );
  INV_X1 _40979_ (
    .A(_06582_),
    .ZN(_06583_)
  );
  AND2_X1 _40980_ (
    .A1(_06545_),
    .A2(_06583_),
    .ZN(_06584_)
  );
  AND2_X1 _40981_ (
    .A1(_21895_),
    .A2(_00007_[2]),
    .ZN(_06585_)
  );
  INV_X1 _40982_ (
    .A(_06585_),
    .ZN(_06586_)
  );
  AND2_X1 _40983_ (
    .A1(_21839_),
    .A2(_22077_),
    .ZN(_06587_)
  );
  INV_X1 _40984_ (
    .A(_06587_),
    .ZN(_06588_)
  );
  AND2_X1 _40985_ (
    .A1(_00007_[0]),
    .A2(_06588_),
    .ZN(_06589_)
  );
  AND2_X1 _40986_ (
    .A1(_06586_),
    .A2(_06589_),
    .ZN(_06590_)
  );
  INV_X1 _40987_ (
    .A(_06590_),
    .ZN(_06591_)
  );
  AND2_X1 _40988_ (
    .A1(_21573_),
    .A2(_22077_),
    .ZN(_06592_)
  );
  INV_X1 _40989_ (
    .A(_06592_),
    .ZN(_06593_)
  );
  AND2_X1 _40990_ (
    .A1(_21911_),
    .A2(_00007_[2]),
    .ZN(_06594_)
  );
  INV_X1 _40991_ (
    .A(_06594_),
    .ZN(_06595_)
  );
  AND2_X1 _40992_ (
    .A1(_06593_),
    .A2(_06595_),
    .ZN(_06596_)
  );
  AND2_X1 _40993_ (
    .A1(_22152_),
    .A2(_06596_),
    .ZN(_06597_)
  );
  INV_X1 _40994_ (
    .A(_06597_),
    .ZN(_06598_)
  );
  AND2_X1 _40995_ (
    .A1(_06591_),
    .A2(_06598_),
    .ZN(_06599_)
  );
  AND2_X1 _40996_ (
    .A1(_22078_),
    .A2(_06599_),
    .ZN(_06600_)
  );
  INV_X1 _40997_ (
    .A(_06600_),
    .ZN(_06601_)
  );
  AND2_X1 _40998_ (
    .A1(_21872_),
    .A2(_22077_),
    .ZN(_06602_)
  );
  INV_X1 _40999_ (
    .A(_06602_),
    .ZN(_06603_)
  );
  AND2_X1 _41000_ (
    .A1(_21855_),
    .A2(_00007_[2]),
    .ZN(_06604_)
  );
  INV_X1 _41001_ (
    .A(_06604_),
    .ZN(_06605_)
  );
  AND2_X1 _41002_ (
    .A1(_06603_),
    .A2(_06605_),
    .ZN(_06606_)
  );
  AND2_X1 _41003_ (
    .A1(_22152_),
    .A2(_06606_),
    .ZN(_06607_)
  );
  INV_X1 _41004_ (
    .A(_06607_),
    .ZN(_06608_)
  );
  AND2_X1 _41005_ (
    .A1(_21943_),
    .A2(_00007_[2]),
    .ZN(_06609_)
  );
  INV_X1 _41006_ (
    .A(_06609_),
    .ZN(_06610_)
  );
  AND2_X1 _41007_ (
    .A1(_21927_),
    .A2(_22077_),
    .ZN(_06611_)
  );
  INV_X1 _41008_ (
    .A(_06611_),
    .ZN(_06612_)
  );
  AND2_X1 _41009_ (
    .A1(_00007_[0]),
    .A2(_06612_),
    .ZN(_06613_)
  );
  AND2_X1 _41010_ (
    .A1(_06610_),
    .A2(_06613_),
    .ZN(_06614_)
  );
  INV_X1 _41011_ (
    .A(_06614_),
    .ZN(_06615_)
  );
  AND2_X1 _41012_ (
    .A1(_06608_),
    .A2(_06615_),
    .ZN(_06616_)
  );
  AND2_X1 _41013_ (
    .A1(_00007_[1]),
    .A2(_06616_),
    .ZN(_06617_)
  );
  INV_X1 _41014_ (
    .A(_06617_),
    .ZN(_06618_)
  );
  AND2_X1 _41015_ (
    .A1(_00007_[3]),
    .A2(_06601_),
    .ZN(_06619_)
  );
  AND2_X1 _41016_ (
    .A1(_06618_),
    .A2(_06619_),
    .ZN(_06620_)
  );
  INV_X1 _41017_ (
    .A(_06620_),
    .ZN(_06621_)
  );
  AND2_X1 _41018_ (
    .A1(_21597_),
    .A2(_22077_),
    .ZN(_06622_)
  );
  INV_X1 _41019_ (
    .A(_06622_),
    .ZN(_06623_)
  );
  AND2_X1 _41020_ (
    .A1(_21417_),
    .A2(_00007_[2]),
    .ZN(_06624_)
  );
  INV_X1 _41021_ (
    .A(_06624_),
    .ZN(_06625_)
  );
  AND2_X1 _41022_ (
    .A1(_21443_),
    .A2(_22077_),
    .ZN(_06626_)
  );
  INV_X1 _41023_ (
    .A(_06626_),
    .ZN(_06627_)
  );
  AND2_X1 _41024_ (
    .A1(_21654_),
    .A2(_00007_[2]),
    .ZN(_06628_)
  );
  INV_X1 _41025_ (
    .A(_06628_),
    .ZN(_06629_)
  );
  AND2_X1 _41026_ (
    .A1(_06627_),
    .A2(_06629_),
    .ZN(_06630_)
  );
  AND2_X1 _41027_ (
    .A1(_21377_),
    .A2(_00007_[2]),
    .ZN(_06631_)
  );
  INV_X1 _41028_ (
    .A(_06631_),
    .ZN(_06632_)
  );
  AND2_X1 _41029_ (
    .A1(_21623_),
    .A2(_22077_),
    .ZN(_06633_)
  );
  INV_X1 _41030_ (
    .A(_06633_),
    .ZN(_06634_)
  );
  AND2_X1 _41031_ (
    .A1(_21465_),
    .A2(_22077_),
    .ZN(_06635_)
  );
  INV_X1 _41032_ (
    .A(_06635_),
    .ZN(_06636_)
  );
  AND2_X1 _41033_ (
    .A1(_21764_),
    .A2(_00007_[2]),
    .ZN(_06637_)
  );
  INV_X1 _41034_ (
    .A(_06637_),
    .ZN(_06638_)
  );
  AND2_X1 _41035_ (
    .A1(_00007_[0]),
    .A2(_06634_),
    .ZN(_06639_)
  );
  AND2_X1 _41036_ (
    .A1(_06632_),
    .A2(_06639_),
    .ZN(_06640_)
  );
  INV_X1 _41037_ (
    .A(_06640_),
    .ZN(_06641_)
  );
  AND2_X1 _41038_ (
    .A1(_22152_),
    .A2(_06623_),
    .ZN(_06642_)
  );
  AND2_X1 _41039_ (
    .A1(_06625_),
    .A2(_06642_),
    .ZN(_06643_)
  );
  INV_X1 _41040_ (
    .A(_06643_),
    .ZN(_06644_)
  );
  AND2_X1 _41041_ (
    .A1(_06641_),
    .A2(_06644_),
    .ZN(_06645_)
  );
  AND2_X1 _41042_ (
    .A1(_00007_[1]),
    .A2(_06645_),
    .ZN(_06646_)
  );
  INV_X1 _41043_ (
    .A(_06646_),
    .ZN(_06647_)
  );
  AND2_X1 _41044_ (
    .A1(_00007_[0]),
    .A2(_06636_),
    .ZN(_06648_)
  );
  AND2_X1 _41045_ (
    .A1(_06638_),
    .A2(_06648_),
    .ZN(_06649_)
  );
  INV_X1 _41046_ (
    .A(_06649_),
    .ZN(_06650_)
  );
  AND2_X1 _41047_ (
    .A1(_22152_),
    .A2(_06630_),
    .ZN(_06651_)
  );
  INV_X1 _41048_ (
    .A(_06651_),
    .ZN(_06652_)
  );
  AND2_X1 _41049_ (
    .A1(_06650_),
    .A2(_06652_),
    .ZN(_06653_)
  );
  AND2_X1 _41050_ (
    .A1(_22078_),
    .A2(_06653_),
    .ZN(_06654_)
  );
  INV_X1 _41051_ (
    .A(_06654_),
    .ZN(_06655_)
  );
  AND2_X1 _41052_ (
    .A1(_06647_),
    .A2(_06655_),
    .ZN(_06656_)
  );
  AND2_X1 _41053_ (
    .A1(_22109_),
    .A2(_06656_),
    .ZN(_06657_)
  );
  INV_X1 _41054_ (
    .A(_06657_),
    .ZN(_06658_)
  );
  AND2_X1 _41055_ (
    .A1(_06621_),
    .A2(_06658_),
    .ZN(_06659_)
  );
  AND2_X1 _41056_ (
    .A1(_22144_),
    .A2(_06584_),
    .ZN(_06660_)
  );
  INV_X1 _41057_ (
    .A(_06660_),
    .ZN(_06661_)
  );
  AND2_X1 _41058_ (
    .A1(_00007_[4]),
    .A2(_06659_),
    .ZN(_06662_)
  );
  INV_X1 _41059_ (
    .A(_06662_),
    .ZN(_06663_)
  );
  AND2_X1 _41060_ (
    .A1(_21209_),
    .A2(_04963_),
    .ZN(_06664_)
  );
  INV_X1 _41061_ (
    .A(_06664_),
    .ZN(_06665_)
  );
  AND2_X1 _41062_ (
    .A1(_05842_),
    .A2(_06663_),
    .ZN(_06666_)
  );
  AND2_X1 _41063_ (
    .A1(_06661_),
    .A2(_06666_),
    .ZN(_06667_)
  );
  INV_X1 _41064_ (
    .A(_06667_),
    .ZN(_06668_)
  );
  AND2_X1 _41065_ (
    .A1(_04962_),
    .A2(_06507_),
    .ZN(_06669_)
  );
  AND2_X1 _41066_ (
    .A1(_06668_),
    .A2(_06669_),
    .ZN(_06670_)
  );
  INV_X1 _41067_ (
    .A(_06670_),
    .ZN(_06671_)
  );
  AND2_X1 _41068_ (
    .A1(_06665_),
    .A2(_06671_),
    .ZN(_00290_)
  );
  AND2_X1 _41069_ (
    .A1(\cpuregs[9] [10]),
    .A2(_22077_),
    .ZN(_06672_)
  );
  INV_X1 _41070_ (
    .A(_06672_),
    .ZN(_06673_)
  );
  AND2_X1 _41071_ (
    .A1(\cpuregs[13] [10]),
    .A2(_00007_[2]),
    .ZN(_06674_)
  );
  INV_X1 _41072_ (
    .A(_06674_),
    .ZN(_06675_)
  );
  AND2_X1 _41073_ (
    .A1(_00007_[0]),
    .A2(_06675_),
    .ZN(_06676_)
  );
  AND2_X1 _41074_ (
    .A1(_06673_),
    .A2(_06676_),
    .ZN(_06677_)
  );
  INV_X1 _41075_ (
    .A(_06677_),
    .ZN(_06678_)
  );
  AND2_X1 _41076_ (
    .A1(\cpuregs[8] [10]),
    .A2(_22077_),
    .ZN(_06679_)
  );
  INV_X1 _41077_ (
    .A(_06679_),
    .ZN(_06680_)
  );
  AND2_X1 _41078_ (
    .A1(\cpuregs[12] [10]),
    .A2(_00007_[2]),
    .ZN(_06681_)
  );
  INV_X1 _41079_ (
    .A(_06681_),
    .ZN(_06682_)
  );
  AND2_X1 _41080_ (
    .A1(_22152_),
    .A2(_06682_),
    .ZN(_06683_)
  );
  AND2_X1 _41081_ (
    .A1(_06680_),
    .A2(_06683_),
    .ZN(_06684_)
  );
  INV_X1 _41082_ (
    .A(_06684_),
    .ZN(_06685_)
  );
  AND2_X1 _41083_ (
    .A1(_22078_),
    .A2(_06685_),
    .ZN(_06686_)
  );
  AND2_X1 _41084_ (
    .A1(_06678_),
    .A2(_06686_),
    .ZN(_06687_)
  );
  INV_X1 _41085_ (
    .A(_06687_),
    .ZN(_06688_)
  );
  AND2_X1 _41086_ (
    .A1(\cpuregs[15] [10]),
    .A2(_00007_[2]),
    .ZN(_06689_)
  );
  INV_X1 _41087_ (
    .A(_06689_),
    .ZN(_06690_)
  );
  AND2_X1 _41088_ (
    .A1(\cpuregs[11] [10]),
    .A2(_22077_),
    .ZN(_06691_)
  );
  INV_X1 _41089_ (
    .A(_06691_),
    .ZN(_06692_)
  );
  AND2_X1 _41090_ (
    .A1(_00007_[0]),
    .A2(_06692_),
    .ZN(_06693_)
  );
  AND2_X1 _41091_ (
    .A1(_06690_),
    .A2(_06693_),
    .ZN(_06694_)
  );
  INV_X1 _41092_ (
    .A(_06694_),
    .ZN(_06695_)
  );
  AND2_X1 _41093_ (
    .A1(\cpuregs[14] [10]),
    .A2(_00007_[2]),
    .ZN(_06696_)
  );
  INV_X1 _41094_ (
    .A(_06696_),
    .ZN(_06697_)
  );
  AND2_X1 _41095_ (
    .A1(\cpuregs[10] [10]),
    .A2(_22077_),
    .ZN(_06698_)
  );
  INV_X1 _41096_ (
    .A(_06698_),
    .ZN(_06699_)
  );
  AND2_X1 _41097_ (
    .A1(_22152_),
    .A2(_06699_),
    .ZN(_06700_)
  );
  AND2_X1 _41098_ (
    .A1(_06697_),
    .A2(_06700_),
    .ZN(_06701_)
  );
  INV_X1 _41099_ (
    .A(_06701_),
    .ZN(_06702_)
  );
  AND2_X1 _41100_ (
    .A1(_00007_[1]),
    .A2(_06702_),
    .ZN(_06703_)
  );
  AND2_X1 _41101_ (
    .A1(_06695_),
    .A2(_06703_),
    .ZN(_06704_)
  );
  INV_X1 _41102_ (
    .A(_06704_),
    .ZN(_06705_)
  );
  AND2_X1 _41103_ (
    .A1(_06688_),
    .A2(_06705_),
    .ZN(_06706_)
  );
  INV_X1 _41104_ (
    .A(_06706_),
    .ZN(_06707_)
  );
  AND2_X1 _41105_ (
    .A1(_00007_[3]),
    .A2(_06707_),
    .ZN(_06708_)
  );
  INV_X1 _41106_ (
    .A(_06708_),
    .ZN(_06709_)
  );
  AND2_X1 _41107_ (
    .A1(\cpuregs[1] [10]),
    .A2(_22077_),
    .ZN(_06710_)
  );
  INV_X1 _41108_ (
    .A(_06710_),
    .ZN(_06711_)
  );
  AND2_X1 _41109_ (
    .A1(\cpuregs[5] [10]),
    .A2(_00007_[2]),
    .ZN(_06712_)
  );
  INV_X1 _41110_ (
    .A(_06712_),
    .ZN(_06713_)
  );
  AND2_X1 _41111_ (
    .A1(_00007_[0]),
    .A2(_06713_),
    .ZN(_06714_)
  );
  AND2_X1 _41112_ (
    .A1(_06711_),
    .A2(_06714_),
    .ZN(_06715_)
  );
  INV_X1 _41113_ (
    .A(_06715_),
    .ZN(_06716_)
  );
  AND2_X1 _41114_ (
    .A1(\cpuregs[0] [10]),
    .A2(_22077_),
    .ZN(_06717_)
  );
  INV_X1 _41115_ (
    .A(_06717_),
    .ZN(_06718_)
  );
  AND2_X1 _41116_ (
    .A1(\cpuregs[4] [10]),
    .A2(_00007_[2]),
    .ZN(_06719_)
  );
  INV_X1 _41117_ (
    .A(_06719_),
    .ZN(_06720_)
  );
  AND2_X1 _41118_ (
    .A1(_22152_),
    .A2(_06720_),
    .ZN(_06721_)
  );
  AND2_X1 _41119_ (
    .A1(_06718_),
    .A2(_06721_),
    .ZN(_06722_)
  );
  INV_X1 _41120_ (
    .A(_06722_),
    .ZN(_06723_)
  );
  AND2_X1 _41121_ (
    .A1(_22078_),
    .A2(_06723_),
    .ZN(_06724_)
  );
  AND2_X1 _41122_ (
    .A1(_06716_),
    .A2(_06724_),
    .ZN(_06725_)
  );
  INV_X1 _41123_ (
    .A(_06725_),
    .ZN(_06726_)
  );
  AND2_X1 _41124_ (
    .A1(\cpuregs[3] [10]),
    .A2(_22077_),
    .ZN(_06727_)
  );
  INV_X1 _41125_ (
    .A(_06727_),
    .ZN(_06728_)
  );
  AND2_X1 _41126_ (
    .A1(\cpuregs[7] [10]),
    .A2(_00007_[2]),
    .ZN(_06729_)
  );
  INV_X1 _41127_ (
    .A(_06729_),
    .ZN(_06730_)
  );
  AND2_X1 _41128_ (
    .A1(_00007_[0]),
    .A2(_06730_),
    .ZN(_06731_)
  );
  AND2_X1 _41129_ (
    .A1(_06728_),
    .A2(_06731_),
    .ZN(_06732_)
  );
  INV_X1 _41130_ (
    .A(_06732_),
    .ZN(_06733_)
  );
  AND2_X1 _41131_ (
    .A1(\cpuregs[6] [10]),
    .A2(_00007_[2]),
    .ZN(_06734_)
  );
  INV_X1 _41132_ (
    .A(_06734_),
    .ZN(_06735_)
  );
  AND2_X1 _41133_ (
    .A1(\cpuregs[2] [10]),
    .A2(_22077_),
    .ZN(_06736_)
  );
  INV_X1 _41134_ (
    .A(_06736_),
    .ZN(_06737_)
  );
  AND2_X1 _41135_ (
    .A1(_22152_),
    .A2(_06737_),
    .ZN(_06738_)
  );
  AND2_X1 _41136_ (
    .A1(_06735_),
    .A2(_06738_),
    .ZN(_06739_)
  );
  INV_X1 _41137_ (
    .A(_06739_),
    .ZN(_06740_)
  );
  AND2_X1 _41138_ (
    .A1(_00007_[1]),
    .A2(_06740_),
    .ZN(_06741_)
  );
  AND2_X1 _41139_ (
    .A1(_06733_),
    .A2(_06741_),
    .ZN(_06742_)
  );
  INV_X1 _41140_ (
    .A(_06742_),
    .ZN(_06743_)
  );
  AND2_X1 _41141_ (
    .A1(_06726_),
    .A2(_06743_),
    .ZN(_06744_)
  );
  INV_X1 _41142_ (
    .A(_06744_),
    .ZN(_06745_)
  );
  AND2_X1 _41143_ (
    .A1(_22109_),
    .A2(_06745_),
    .ZN(_06746_)
  );
  INV_X1 _41144_ (
    .A(_06746_),
    .ZN(_06747_)
  );
  AND2_X1 _41145_ (
    .A1(_06709_),
    .A2(_06747_),
    .ZN(_06748_)
  );
  AND2_X1 _41146_ (
    .A1(\cpuregs[29] [10]),
    .A2(_00007_[2]),
    .ZN(_06749_)
  );
  INV_X1 _41147_ (
    .A(_06749_),
    .ZN(_06750_)
  );
  AND2_X1 _41148_ (
    .A1(\cpuregs[25] [10]),
    .A2(_22077_),
    .ZN(_06751_)
  );
  INV_X1 _41149_ (
    .A(_06751_),
    .ZN(_06752_)
  );
  AND2_X1 _41150_ (
    .A1(_00007_[0]),
    .A2(_06752_),
    .ZN(_06753_)
  );
  AND2_X1 _41151_ (
    .A1(_06750_),
    .A2(_06753_),
    .ZN(_06754_)
  );
  INV_X1 _41152_ (
    .A(_06754_),
    .ZN(_06755_)
  );
  AND2_X1 _41153_ (
    .A1(\cpuregs[28] [10]),
    .A2(_00007_[2]),
    .ZN(_06756_)
  );
  INV_X1 _41154_ (
    .A(_06756_),
    .ZN(_06757_)
  );
  AND2_X1 _41155_ (
    .A1(\cpuregs[24] [10]),
    .A2(_22077_),
    .ZN(_06758_)
  );
  INV_X1 _41156_ (
    .A(_06758_),
    .ZN(_06759_)
  );
  AND2_X1 _41157_ (
    .A1(_22152_),
    .A2(_06759_),
    .ZN(_06760_)
  );
  AND2_X1 _41158_ (
    .A1(_06757_),
    .A2(_06760_),
    .ZN(_06761_)
  );
  INV_X1 _41159_ (
    .A(_06761_),
    .ZN(_06762_)
  );
  AND2_X1 _41160_ (
    .A1(_22078_),
    .A2(_06762_),
    .ZN(_06763_)
  );
  AND2_X1 _41161_ (
    .A1(_06755_),
    .A2(_06763_),
    .ZN(_06764_)
  );
  INV_X1 _41162_ (
    .A(_06764_),
    .ZN(_06765_)
  );
  AND2_X1 _41163_ (
    .A1(\cpuregs[27] [10]),
    .A2(_22077_),
    .ZN(_06766_)
  );
  INV_X1 _41164_ (
    .A(_06766_),
    .ZN(_06767_)
  );
  AND2_X1 _41165_ (
    .A1(\cpuregs[31] [10]),
    .A2(_00007_[2]),
    .ZN(_06768_)
  );
  INV_X1 _41166_ (
    .A(_06768_),
    .ZN(_06769_)
  );
  AND2_X1 _41167_ (
    .A1(_00007_[0]),
    .A2(_06769_),
    .ZN(_06770_)
  );
  AND2_X1 _41168_ (
    .A1(_06767_),
    .A2(_06770_),
    .ZN(_06771_)
  );
  INV_X1 _41169_ (
    .A(_06771_),
    .ZN(_06772_)
  );
  AND2_X1 _41170_ (
    .A1(\cpuregs[26] [10]),
    .A2(_22077_),
    .ZN(_06773_)
  );
  INV_X1 _41171_ (
    .A(_06773_),
    .ZN(_06774_)
  );
  AND2_X1 _41172_ (
    .A1(\cpuregs[30] [10]),
    .A2(_00007_[2]),
    .ZN(_06775_)
  );
  INV_X1 _41173_ (
    .A(_06775_),
    .ZN(_06776_)
  );
  AND2_X1 _41174_ (
    .A1(_22152_),
    .A2(_06776_),
    .ZN(_06777_)
  );
  AND2_X1 _41175_ (
    .A1(_06774_),
    .A2(_06777_),
    .ZN(_06778_)
  );
  INV_X1 _41176_ (
    .A(_06778_),
    .ZN(_06779_)
  );
  AND2_X1 _41177_ (
    .A1(_00007_[1]),
    .A2(_06779_),
    .ZN(_06780_)
  );
  AND2_X1 _41178_ (
    .A1(_06772_),
    .A2(_06780_),
    .ZN(_06781_)
  );
  INV_X1 _41179_ (
    .A(_06781_),
    .ZN(_06782_)
  );
  AND2_X1 _41180_ (
    .A1(_06765_),
    .A2(_06782_),
    .ZN(_06783_)
  );
  INV_X1 _41181_ (
    .A(_06783_),
    .ZN(_06784_)
  );
  AND2_X1 _41182_ (
    .A1(_00007_[3]),
    .A2(_06784_),
    .ZN(_06785_)
  );
  INV_X1 _41183_ (
    .A(_06785_),
    .ZN(_06786_)
  );
  AND2_X1 _41184_ (
    .A1(_21378_),
    .A2(_00007_[2]),
    .ZN(_06787_)
  );
  INV_X1 _41185_ (
    .A(_06787_),
    .ZN(_06788_)
  );
  AND2_X1 _41186_ (
    .A1(_21624_),
    .A2(_22077_),
    .ZN(_06789_)
  );
  INV_X1 _41187_ (
    .A(_06789_),
    .ZN(_06790_)
  );
  AND2_X1 _41188_ (
    .A1(_00007_[0]),
    .A2(_06790_),
    .ZN(_06791_)
  );
  AND2_X1 _41189_ (
    .A1(_06788_),
    .A2(_06791_),
    .ZN(_06792_)
  );
  INV_X1 _41190_ (
    .A(_06792_),
    .ZN(_06793_)
  );
  AND2_X1 _41191_ (
    .A1(_21418_),
    .A2(_00007_[2]),
    .ZN(_06794_)
  );
  INV_X1 _41192_ (
    .A(_06794_),
    .ZN(_06795_)
  );
  AND2_X1 _41193_ (
    .A1(_21598_),
    .A2(_22077_),
    .ZN(_06796_)
  );
  INV_X1 _41194_ (
    .A(_06796_),
    .ZN(_06797_)
  );
  AND2_X1 _41195_ (
    .A1(_22152_),
    .A2(_06797_),
    .ZN(_06798_)
  );
  AND2_X1 _41196_ (
    .A1(_06795_),
    .A2(_06798_),
    .ZN(_06799_)
  );
  INV_X1 _41197_ (
    .A(_06799_),
    .ZN(_06800_)
  );
  AND2_X1 _41198_ (
    .A1(_06793_),
    .A2(_06800_),
    .ZN(_06801_)
  );
  AND2_X1 _41199_ (
    .A1(_00007_[1]),
    .A2(_06801_),
    .ZN(_06802_)
  );
  INV_X1 _41200_ (
    .A(_06802_),
    .ZN(_06803_)
  );
  AND2_X1 _41201_ (
    .A1(_21765_),
    .A2(_00007_[2]),
    .ZN(_06804_)
  );
  INV_X1 _41202_ (
    .A(_06804_),
    .ZN(_06805_)
  );
  AND2_X1 _41203_ (
    .A1(_21466_),
    .A2(_22077_),
    .ZN(_06806_)
  );
  INV_X1 _41204_ (
    .A(_06806_),
    .ZN(_06807_)
  );
  AND2_X1 _41205_ (
    .A1(_00007_[0]),
    .A2(_06807_),
    .ZN(_06808_)
  );
  AND2_X1 _41206_ (
    .A1(_06805_),
    .A2(_06808_),
    .ZN(_06809_)
  );
  INV_X1 _41207_ (
    .A(_06809_),
    .ZN(_06810_)
  );
  AND2_X1 _41208_ (
    .A1(_21444_),
    .A2(_22077_),
    .ZN(_06811_)
  );
  INV_X1 _41209_ (
    .A(_06811_),
    .ZN(_06812_)
  );
  AND2_X1 _41210_ (
    .A1(_21655_),
    .A2(_00007_[2]),
    .ZN(_06813_)
  );
  INV_X1 _41211_ (
    .A(_06813_),
    .ZN(_06814_)
  );
  AND2_X1 _41212_ (
    .A1(_06812_),
    .A2(_06814_),
    .ZN(_06815_)
  );
  AND2_X1 _41213_ (
    .A1(_22152_),
    .A2(_06815_),
    .ZN(_06816_)
  );
  INV_X1 _41214_ (
    .A(_06816_),
    .ZN(_06817_)
  );
  AND2_X1 _41215_ (
    .A1(_06810_),
    .A2(_06817_),
    .ZN(_06818_)
  );
  AND2_X1 _41216_ (
    .A1(_22078_),
    .A2(_06818_),
    .ZN(_06819_)
  );
  INV_X1 _41217_ (
    .A(_06819_),
    .ZN(_06820_)
  );
  AND2_X1 _41218_ (
    .A1(_06803_),
    .A2(_06820_),
    .ZN(_06821_)
  );
  AND2_X1 _41219_ (
    .A1(_22109_),
    .A2(_06821_),
    .ZN(_06822_)
  );
  INV_X1 _41220_ (
    .A(_06822_),
    .ZN(_06823_)
  );
  AND2_X1 _41221_ (
    .A1(_22144_),
    .A2(_06748_),
    .ZN(_06824_)
  );
  INV_X1 _41222_ (
    .A(_06824_),
    .ZN(_06825_)
  );
  AND2_X1 _41223_ (
    .A1(_00007_[4]),
    .A2(_06823_),
    .ZN(_06826_)
  );
  AND2_X1 _41224_ (
    .A1(_06786_),
    .A2(_06826_),
    .ZN(_06827_)
  );
  INV_X1 _41225_ (
    .A(_06827_),
    .ZN(_06828_)
  );
  AND2_X1 _41226_ (
    .A1(decoded_imm[10]),
    .A2(_04966_),
    .ZN(_06829_)
  );
  INV_X1 _41227_ (
    .A(_06829_),
    .ZN(_06830_)
  );
  AND2_X1 _41228_ (
    .A1(_04962_),
    .A2(_06830_),
    .ZN(_06831_)
  );
  AND2_X1 _41229_ (
    .A1(_05842_),
    .A2(_06828_),
    .ZN(_06832_)
  );
  AND2_X1 _41230_ (
    .A1(_06825_),
    .A2(_06832_),
    .ZN(_06833_)
  );
  INV_X1 _41231_ (
    .A(_06833_),
    .ZN(_06834_)
  );
  AND2_X1 _41232_ (
    .A1(_06831_),
    .A2(_06834_),
    .ZN(_06835_)
  );
  INV_X1 _41233_ (
    .A(_06835_),
    .ZN(_06836_)
  );
  AND2_X1 _41234_ (
    .A1(_21210_),
    .A2(_04963_),
    .ZN(_06837_)
  );
  INV_X1 _41235_ (
    .A(_06837_),
    .ZN(_06838_)
  );
  AND2_X1 _41236_ (
    .A1(_06836_),
    .A2(_06838_),
    .ZN(_00291_)
  );
  AND2_X1 _41237_ (
    .A1(decoded_imm[11]),
    .A2(_04966_),
    .ZN(_06839_)
  );
  INV_X1 _41238_ (
    .A(_06839_),
    .ZN(_06840_)
  );
  AND2_X1 _41239_ (
    .A1(\cpuregs[19] [11]),
    .A2(_22077_),
    .ZN(_06841_)
  );
  INV_X1 _41240_ (
    .A(_06841_),
    .ZN(_06842_)
  );
  AND2_X1 _41241_ (
    .A1(\cpuregs[23] [11]),
    .A2(_00007_[2]),
    .ZN(_06843_)
  );
  INV_X1 _41242_ (
    .A(_06843_),
    .ZN(_06844_)
  );
  AND2_X1 _41243_ (
    .A1(_06842_),
    .A2(_06844_),
    .ZN(_06845_)
  );
  INV_X1 _41244_ (
    .A(_06845_),
    .ZN(_06846_)
  );
  AND2_X1 _41245_ (
    .A1(_00007_[0]),
    .A2(_06846_),
    .ZN(_06847_)
  );
  INV_X1 _41246_ (
    .A(_06847_),
    .ZN(_06848_)
  );
  AND2_X1 _41247_ (
    .A1(\cpuregs[22] [11]),
    .A2(_00007_[2]),
    .ZN(_06849_)
  );
  INV_X1 _41248_ (
    .A(_06849_),
    .ZN(_06850_)
  );
  AND2_X1 _41249_ (
    .A1(\cpuregs[18] [11]),
    .A2(_22077_),
    .ZN(_06851_)
  );
  INV_X1 _41250_ (
    .A(_06851_),
    .ZN(_06852_)
  );
  AND2_X1 _41251_ (
    .A1(_06850_),
    .A2(_06852_),
    .ZN(_06853_)
  );
  INV_X1 _41252_ (
    .A(_06853_),
    .ZN(_06854_)
  );
  AND2_X1 _41253_ (
    .A1(_22152_),
    .A2(_06854_),
    .ZN(_06855_)
  );
  INV_X1 _41254_ (
    .A(_06855_),
    .ZN(_06856_)
  );
  AND2_X1 _41255_ (
    .A1(_21496_),
    .A2(_22077_),
    .ZN(_06857_)
  );
  INV_X1 _41256_ (
    .A(_06857_),
    .ZN(_06858_)
  );
  AND2_X1 _41257_ (
    .A1(_21788_),
    .A2(_00007_[2]),
    .ZN(_06859_)
  );
  INV_X1 _41258_ (
    .A(_06859_),
    .ZN(_06860_)
  );
  AND2_X1 _41259_ (
    .A1(_00007_[0]),
    .A2(_06860_),
    .ZN(_06861_)
  );
  AND2_X1 _41260_ (
    .A1(_06858_),
    .A2(_06861_),
    .ZN(_06862_)
  );
  INV_X1 _41261_ (
    .A(_06862_),
    .ZN(_06863_)
  );
  AND2_X1 _41262_ (
    .A1(_21814_),
    .A2(_00007_[2]),
    .ZN(_06864_)
  );
  INV_X1 _41263_ (
    .A(_06864_),
    .ZN(_06865_)
  );
  AND2_X1 _41264_ (
    .A1(_21548_),
    .A2(_22077_),
    .ZN(_06866_)
  );
  INV_X1 _41265_ (
    .A(_06866_),
    .ZN(_06867_)
  );
  AND2_X1 _41266_ (
    .A1(_22152_),
    .A2(_06867_),
    .ZN(_06868_)
  );
  AND2_X1 _41267_ (
    .A1(_06865_),
    .A2(_06868_),
    .ZN(_06869_)
  );
  INV_X1 _41268_ (
    .A(_06869_),
    .ZN(_06870_)
  );
  AND2_X1 _41269_ (
    .A1(\cpuregs[17] [11]),
    .A2(_22077_),
    .ZN(_06871_)
  );
  INV_X1 _41270_ (
    .A(_06871_),
    .ZN(_06872_)
  );
  AND2_X1 _41271_ (
    .A1(\cpuregs[21] [11]),
    .A2(_00007_[2]),
    .ZN(_06873_)
  );
  INV_X1 _41272_ (
    .A(_06873_),
    .ZN(_06874_)
  );
  AND2_X1 _41273_ (
    .A1(_06872_),
    .A2(_06874_),
    .ZN(_06875_)
  );
  INV_X1 _41274_ (
    .A(_06875_),
    .ZN(_06876_)
  );
  AND2_X1 _41275_ (
    .A1(_00007_[0]),
    .A2(_06876_),
    .ZN(_06877_)
  );
  INV_X1 _41276_ (
    .A(_06877_),
    .ZN(_06878_)
  );
  AND2_X1 _41277_ (
    .A1(\cpuregs[16] [11]),
    .A2(_22077_),
    .ZN(_06879_)
  );
  INV_X1 _41278_ (
    .A(_06879_),
    .ZN(_06880_)
  );
  AND2_X1 _41279_ (
    .A1(\cpuregs[20] [11]),
    .A2(_00007_[2]),
    .ZN(_06881_)
  );
  INV_X1 _41280_ (
    .A(_06881_),
    .ZN(_06882_)
  );
  AND2_X1 _41281_ (
    .A1(_06880_),
    .A2(_06882_),
    .ZN(_06883_)
  );
  INV_X1 _41282_ (
    .A(_06883_),
    .ZN(_06884_)
  );
  AND2_X1 _41283_ (
    .A1(_22152_),
    .A2(_06884_),
    .ZN(_06885_)
  );
  INV_X1 _41284_ (
    .A(_06885_),
    .ZN(_06886_)
  );
  AND2_X1 _41285_ (
    .A1(_06878_),
    .A2(_06886_),
    .ZN(_06887_)
  );
  AND2_X1 _41286_ (
    .A1(_21521_),
    .A2(_22077_),
    .ZN(_06888_)
  );
  INV_X1 _41287_ (
    .A(_06888_),
    .ZN(_06889_)
  );
  AND2_X1 _41288_ (
    .A1(_21741_),
    .A2(_00007_[2]),
    .ZN(_06890_)
  );
  INV_X1 _41289_ (
    .A(_06890_),
    .ZN(_06891_)
  );
  AND2_X1 _41290_ (
    .A1(_00007_[0]),
    .A2(_06891_),
    .ZN(_06892_)
  );
  AND2_X1 _41291_ (
    .A1(_06889_),
    .A2(_06892_),
    .ZN(_06893_)
  );
  INV_X1 _41292_ (
    .A(_06893_),
    .ZN(_06894_)
  );
  AND2_X1 _41293_ (
    .A1(_21962_),
    .A2(_22077_),
    .ZN(_06895_)
  );
  INV_X1 _41294_ (
    .A(_06895_),
    .ZN(_06896_)
  );
  AND2_X1 _41295_ (
    .A1(_21678_),
    .A2(_00007_[2]),
    .ZN(_06897_)
  );
  INV_X1 _41296_ (
    .A(_06897_),
    .ZN(_06898_)
  );
  AND2_X1 _41297_ (
    .A1(_06896_),
    .A2(_06898_),
    .ZN(_06899_)
  );
  AND2_X1 _41298_ (
    .A1(_22152_),
    .A2(_06899_),
    .ZN(_06900_)
  );
  INV_X1 _41299_ (
    .A(_06900_),
    .ZN(_06901_)
  );
  AND2_X1 _41300_ (
    .A1(_06894_),
    .A2(_06901_),
    .ZN(_06902_)
  );
  AND2_X1 _41301_ (
    .A1(_22078_),
    .A2(_06902_),
    .ZN(_06903_)
  );
  INV_X1 _41302_ (
    .A(_06903_),
    .ZN(_06904_)
  );
  AND2_X1 _41303_ (
    .A1(_00007_[1]),
    .A2(_06870_),
    .ZN(_06905_)
  );
  AND2_X1 _41304_ (
    .A1(_06863_),
    .A2(_06905_),
    .ZN(_06906_)
  );
  INV_X1 _41305_ (
    .A(_06906_),
    .ZN(_06907_)
  );
  AND2_X1 _41306_ (
    .A1(_06904_),
    .A2(_06907_),
    .ZN(_06908_)
  );
  AND2_X1 _41307_ (
    .A1(_22144_),
    .A2(_06908_),
    .ZN(_06909_)
  );
  INV_X1 _41308_ (
    .A(_06909_),
    .ZN(_06910_)
  );
  AND2_X1 _41309_ (
    .A1(_00007_[1]),
    .A2(_06856_),
    .ZN(_06911_)
  );
  AND2_X1 _41310_ (
    .A1(_06848_),
    .A2(_06911_),
    .ZN(_06912_)
  );
  INV_X1 _41311_ (
    .A(_06912_),
    .ZN(_06913_)
  );
  AND2_X1 _41312_ (
    .A1(_22078_),
    .A2(_06887_),
    .ZN(_06914_)
  );
  INV_X1 _41313_ (
    .A(_06914_),
    .ZN(_06915_)
  );
  AND2_X1 _41314_ (
    .A1(_06913_),
    .A2(_06915_),
    .ZN(_06916_)
  );
  AND2_X1 _41315_ (
    .A1(_00007_[4]),
    .A2(_06916_),
    .ZN(_06917_)
  );
  INV_X1 _41316_ (
    .A(_06917_),
    .ZN(_06918_)
  );
  AND2_X1 _41317_ (
    .A1(_06910_),
    .A2(_06918_),
    .ZN(_06919_)
  );
  AND2_X1 _41318_ (
    .A1(\cpuregs[26] [11]),
    .A2(_22077_),
    .ZN(_06920_)
  );
  INV_X1 _41319_ (
    .A(_06920_),
    .ZN(_06921_)
  );
  AND2_X1 _41320_ (
    .A1(\cpuregs[30] [11]),
    .A2(_00007_[2]),
    .ZN(_06922_)
  );
  INV_X1 _41321_ (
    .A(_06922_),
    .ZN(_06923_)
  );
  AND2_X1 _41322_ (
    .A1(_00007_[1]),
    .A2(_06923_),
    .ZN(_06924_)
  );
  AND2_X1 _41323_ (
    .A1(_06921_),
    .A2(_06924_),
    .ZN(_06925_)
  );
  INV_X1 _41324_ (
    .A(_06925_),
    .ZN(_06926_)
  );
  AND2_X1 _41325_ (
    .A1(\cpuregs[28] [11]),
    .A2(_00007_[2]),
    .ZN(_06927_)
  );
  INV_X1 _41326_ (
    .A(_06927_),
    .ZN(_06928_)
  );
  AND2_X1 _41327_ (
    .A1(\cpuregs[24] [11]),
    .A2(_22077_),
    .ZN(_06929_)
  );
  INV_X1 _41328_ (
    .A(_06929_),
    .ZN(_06930_)
  );
  AND2_X1 _41329_ (
    .A1(_22078_),
    .A2(_06930_),
    .ZN(_06931_)
  );
  AND2_X1 _41330_ (
    .A1(_06928_),
    .A2(_06931_),
    .ZN(_06932_)
  );
  INV_X1 _41331_ (
    .A(_06932_),
    .ZN(_06933_)
  );
  AND2_X1 _41332_ (
    .A1(_22152_),
    .A2(_06933_),
    .ZN(_06934_)
  );
  AND2_X1 _41333_ (
    .A1(_06926_),
    .A2(_06934_),
    .ZN(_06935_)
  );
  INV_X1 _41334_ (
    .A(_06935_),
    .ZN(_06936_)
  );
  AND2_X1 _41335_ (
    .A1(\cpuregs[27] [11]),
    .A2(_22077_),
    .ZN(_06937_)
  );
  INV_X1 _41336_ (
    .A(_06937_),
    .ZN(_06938_)
  );
  AND2_X1 _41337_ (
    .A1(\cpuregs[31] [11]),
    .A2(_00007_[2]),
    .ZN(_06939_)
  );
  INV_X1 _41338_ (
    .A(_06939_),
    .ZN(_06940_)
  );
  AND2_X1 _41339_ (
    .A1(_00007_[1]),
    .A2(_06940_),
    .ZN(_06941_)
  );
  AND2_X1 _41340_ (
    .A1(_06938_),
    .A2(_06941_),
    .ZN(_06942_)
  );
  INV_X1 _41341_ (
    .A(_06942_),
    .ZN(_06943_)
  );
  AND2_X1 _41342_ (
    .A1(\cpuregs[29] [11]),
    .A2(_00007_[2]),
    .ZN(_06944_)
  );
  INV_X1 _41343_ (
    .A(_06944_),
    .ZN(_06945_)
  );
  AND2_X1 _41344_ (
    .A1(\cpuregs[25] [11]),
    .A2(_22077_),
    .ZN(_06946_)
  );
  INV_X1 _41345_ (
    .A(_06946_),
    .ZN(_06947_)
  );
  AND2_X1 _41346_ (
    .A1(_22078_),
    .A2(_06947_),
    .ZN(_06948_)
  );
  AND2_X1 _41347_ (
    .A1(_06945_),
    .A2(_06948_),
    .ZN(_06949_)
  );
  INV_X1 _41348_ (
    .A(_06949_),
    .ZN(_06950_)
  );
  AND2_X1 _41349_ (
    .A1(_00007_[0]),
    .A2(_06950_),
    .ZN(_06951_)
  );
  AND2_X1 _41350_ (
    .A1(_06943_),
    .A2(_06951_),
    .ZN(_06952_)
  );
  INV_X1 _41351_ (
    .A(_06952_),
    .ZN(_06953_)
  );
  AND2_X1 _41352_ (
    .A1(_06936_),
    .A2(_06953_),
    .ZN(_06954_)
  );
  INV_X1 _41353_ (
    .A(_06954_),
    .ZN(_06955_)
  );
  AND2_X1 _41354_ (
    .A1(_00007_[4]),
    .A2(_06955_),
    .ZN(_06956_)
  );
  INV_X1 _41355_ (
    .A(_06956_),
    .ZN(_06957_)
  );
  AND2_X1 _41356_ (
    .A1(\cpuregs[12] [11]),
    .A2(_22078_),
    .ZN(_06958_)
  );
  INV_X1 _41357_ (
    .A(_06958_),
    .ZN(_06959_)
  );
  AND2_X1 _41358_ (
    .A1(\cpuregs[14] [11]),
    .A2(_00007_[1]),
    .ZN(_06960_)
  );
  INV_X1 _41359_ (
    .A(_06960_),
    .ZN(_06961_)
  );
  AND2_X1 _41360_ (
    .A1(_00007_[2]),
    .A2(_06961_),
    .ZN(_06962_)
  );
  AND2_X1 _41361_ (
    .A1(_06959_),
    .A2(_06962_),
    .ZN(_06963_)
  );
  INV_X1 _41362_ (
    .A(_06963_),
    .ZN(_06964_)
  );
  AND2_X1 _41363_ (
    .A1(\cpuregs[8] [11]),
    .A2(_22078_),
    .ZN(_06965_)
  );
  INV_X1 _41364_ (
    .A(_06965_),
    .ZN(_06966_)
  );
  AND2_X1 _41365_ (
    .A1(\cpuregs[10] [11]),
    .A2(_00007_[1]),
    .ZN(_06967_)
  );
  INV_X1 _41366_ (
    .A(_06967_),
    .ZN(_06968_)
  );
  AND2_X1 _41367_ (
    .A1(_22077_),
    .A2(_06968_),
    .ZN(_06969_)
  );
  AND2_X1 _41368_ (
    .A1(_06966_),
    .A2(_06969_),
    .ZN(_06970_)
  );
  INV_X1 _41369_ (
    .A(_06970_),
    .ZN(_06971_)
  );
  AND2_X1 _41370_ (
    .A1(_22152_),
    .A2(_06971_),
    .ZN(_06972_)
  );
  AND2_X1 _41371_ (
    .A1(_06964_),
    .A2(_06972_),
    .ZN(_06973_)
  );
  INV_X1 _41372_ (
    .A(_06973_),
    .ZN(_06974_)
  );
  AND2_X1 _41373_ (
    .A1(\cpuregs[13] [11]),
    .A2(_22078_),
    .ZN(_06975_)
  );
  INV_X1 _41374_ (
    .A(_06975_),
    .ZN(_06976_)
  );
  AND2_X1 _41375_ (
    .A1(\cpuregs[15] [11]),
    .A2(_00007_[1]),
    .ZN(_06977_)
  );
  INV_X1 _41376_ (
    .A(_06977_),
    .ZN(_06978_)
  );
  AND2_X1 _41377_ (
    .A1(_00007_[2]),
    .A2(_06978_),
    .ZN(_06979_)
  );
  AND2_X1 _41378_ (
    .A1(_06976_),
    .A2(_06979_),
    .ZN(_06980_)
  );
  INV_X1 _41379_ (
    .A(_06980_),
    .ZN(_06981_)
  );
  AND2_X1 _41380_ (
    .A1(\cpuregs[9] [11]),
    .A2(_22078_),
    .ZN(_06982_)
  );
  INV_X1 _41381_ (
    .A(_06982_),
    .ZN(_06983_)
  );
  AND2_X1 _41382_ (
    .A1(\cpuregs[11] [11]),
    .A2(_00007_[1]),
    .ZN(_06984_)
  );
  INV_X1 _41383_ (
    .A(_06984_),
    .ZN(_06985_)
  );
  AND2_X1 _41384_ (
    .A1(_22077_),
    .A2(_06985_),
    .ZN(_06986_)
  );
  AND2_X1 _41385_ (
    .A1(_06983_),
    .A2(_06986_),
    .ZN(_06987_)
  );
  INV_X1 _41386_ (
    .A(_06987_),
    .ZN(_06988_)
  );
  AND2_X1 _41387_ (
    .A1(_00007_[0]),
    .A2(_06988_),
    .ZN(_06989_)
  );
  AND2_X1 _41388_ (
    .A1(_06981_),
    .A2(_06989_),
    .ZN(_06990_)
  );
  INV_X1 _41389_ (
    .A(_06990_),
    .ZN(_06991_)
  );
  AND2_X1 _41390_ (
    .A1(_06974_),
    .A2(_06991_),
    .ZN(_06992_)
  );
  INV_X1 _41391_ (
    .A(_06992_),
    .ZN(_06993_)
  );
  AND2_X1 _41392_ (
    .A1(_22144_),
    .A2(_06993_),
    .ZN(_06994_)
  );
  INV_X1 _41393_ (
    .A(_06994_),
    .ZN(_06995_)
  );
  AND2_X1 _41394_ (
    .A1(_00007_[3]),
    .A2(_06995_),
    .ZN(_06996_)
  );
  AND2_X1 _41395_ (
    .A1(_06957_),
    .A2(_06996_),
    .ZN(_06997_)
  );
  INV_X1 _41396_ (
    .A(_06997_),
    .ZN(_06998_)
  );
  AND2_X1 _41397_ (
    .A1(_22109_),
    .A2(_06919_),
    .ZN(_06999_)
  );
  INV_X1 _41398_ (
    .A(_06999_),
    .ZN(_07000_)
  );
  AND2_X1 _41399_ (
    .A1(_06998_),
    .A2(_07000_),
    .ZN(_07001_)
  );
  AND2_X1 _41400_ (
    .A1(_05842_),
    .A2(_07001_),
    .ZN(_07002_)
  );
  INV_X1 _41401_ (
    .A(_07002_),
    .ZN(_07003_)
  );
  AND2_X1 _41402_ (
    .A1(_21211_),
    .A2(_04963_),
    .ZN(_07004_)
  );
  INV_X1 _41403_ (
    .A(_07004_),
    .ZN(_07005_)
  );
  AND2_X1 _41404_ (
    .A1(_04962_),
    .A2(_07003_),
    .ZN(_07006_)
  );
  AND2_X1 _41405_ (
    .A1(_06840_),
    .A2(_07006_),
    .ZN(_07007_)
  );
  INV_X1 _41406_ (
    .A(_07007_),
    .ZN(_07008_)
  );
  AND2_X1 _41407_ (
    .A1(_07005_),
    .A2(_07008_),
    .ZN(_00292_)
  );
  AND2_X1 _41408_ (
    .A1(decoded_imm[12]),
    .A2(_04966_),
    .ZN(_07009_)
  );
  INV_X1 _41409_ (
    .A(_07009_),
    .ZN(_07010_)
  );
  AND2_X1 _41410_ (
    .A1(\cpuregs[29] [12]),
    .A2(_00007_[2]),
    .ZN(_07011_)
  );
  INV_X1 _41411_ (
    .A(_07011_),
    .ZN(_07012_)
  );
  AND2_X1 _41412_ (
    .A1(\cpuregs[25] [12]),
    .A2(_22077_),
    .ZN(_07013_)
  );
  INV_X1 _41413_ (
    .A(_07013_),
    .ZN(_07014_)
  );
  AND2_X1 _41414_ (
    .A1(_00007_[0]),
    .A2(_07014_),
    .ZN(_07015_)
  );
  AND2_X1 _41415_ (
    .A1(_07012_),
    .A2(_07015_),
    .ZN(_07016_)
  );
  INV_X1 _41416_ (
    .A(_07016_),
    .ZN(_07017_)
  );
  AND2_X1 _41417_ (
    .A1(\cpuregs[24] [12]),
    .A2(_22077_),
    .ZN(_07018_)
  );
  INV_X1 _41418_ (
    .A(_07018_),
    .ZN(_07019_)
  );
  AND2_X1 _41419_ (
    .A1(\cpuregs[28] [12]),
    .A2(_00007_[2]),
    .ZN(_07020_)
  );
  INV_X1 _41420_ (
    .A(_07020_),
    .ZN(_07021_)
  );
  AND2_X1 _41421_ (
    .A1(_22152_),
    .A2(_07021_),
    .ZN(_07022_)
  );
  AND2_X1 _41422_ (
    .A1(_07019_),
    .A2(_07022_),
    .ZN(_07023_)
  );
  INV_X1 _41423_ (
    .A(_07023_),
    .ZN(_07024_)
  );
  AND2_X1 _41424_ (
    .A1(_22078_),
    .A2(_07024_),
    .ZN(_07025_)
  );
  AND2_X1 _41425_ (
    .A1(_07017_),
    .A2(_07025_),
    .ZN(_07026_)
  );
  INV_X1 _41426_ (
    .A(_07026_),
    .ZN(_07027_)
  );
  AND2_X1 _41427_ (
    .A1(\cpuregs[31] [12]),
    .A2(_00007_[2]),
    .ZN(_07028_)
  );
  INV_X1 _41428_ (
    .A(_07028_),
    .ZN(_07029_)
  );
  AND2_X1 _41429_ (
    .A1(\cpuregs[27] [12]),
    .A2(_22077_),
    .ZN(_07030_)
  );
  INV_X1 _41430_ (
    .A(_07030_),
    .ZN(_07031_)
  );
  AND2_X1 _41431_ (
    .A1(_00007_[0]),
    .A2(_07031_),
    .ZN(_07032_)
  );
  AND2_X1 _41432_ (
    .A1(_07029_),
    .A2(_07032_),
    .ZN(_07033_)
  );
  INV_X1 _41433_ (
    .A(_07033_),
    .ZN(_07034_)
  );
  AND2_X1 _41434_ (
    .A1(\cpuregs[26] [12]),
    .A2(_22077_),
    .ZN(_07035_)
  );
  INV_X1 _41435_ (
    .A(_07035_),
    .ZN(_07036_)
  );
  AND2_X1 _41436_ (
    .A1(\cpuregs[30] [12]),
    .A2(_00007_[2]),
    .ZN(_07037_)
  );
  INV_X1 _41437_ (
    .A(_07037_),
    .ZN(_07038_)
  );
  AND2_X1 _41438_ (
    .A1(_22152_),
    .A2(_07038_),
    .ZN(_07039_)
  );
  AND2_X1 _41439_ (
    .A1(_07036_),
    .A2(_07039_),
    .ZN(_07040_)
  );
  INV_X1 _41440_ (
    .A(_07040_),
    .ZN(_07041_)
  );
  AND2_X1 _41441_ (
    .A1(_00007_[1]),
    .A2(_07041_),
    .ZN(_07042_)
  );
  AND2_X1 _41442_ (
    .A1(_07034_),
    .A2(_07042_),
    .ZN(_07043_)
  );
  INV_X1 _41443_ (
    .A(_07043_),
    .ZN(_07044_)
  );
  AND2_X1 _41444_ (
    .A1(_07027_),
    .A2(_07044_),
    .ZN(_07045_)
  );
  INV_X1 _41445_ (
    .A(_07045_),
    .ZN(_07046_)
  );
  AND2_X1 _41446_ (
    .A1(\cpuregs[11] [12]),
    .A2(_22077_),
    .ZN(_07047_)
  );
  INV_X1 _41447_ (
    .A(_07047_),
    .ZN(_07048_)
  );
  AND2_X1 _41448_ (
    .A1(\cpuregs[15] [12]),
    .A2(_00007_[2]),
    .ZN(_07049_)
  );
  INV_X1 _41449_ (
    .A(_07049_),
    .ZN(_07050_)
  );
  AND2_X1 _41450_ (
    .A1(_07048_),
    .A2(_07050_),
    .ZN(_07051_)
  );
  INV_X1 _41451_ (
    .A(_07051_),
    .ZN(_07052_)
  );
  AND2_X1 _41452_ (
    .A1(_00007_[0]),
    .A2(_07052_),
    .ZN(_07053_)
  );
  INV_X1 _41453_ (
    .A(_07053_),
    .ZN(_07054_)
  );
  AND2_X1 _41454_ (
    .A1(\cpuregs[14] [12]),
    .A2(_00007_[2]),
    .ZN(_07055_)
  );
  INV_X1 _41455_ (
    .A(_07055_),
    .ZN(_07056_)
  );
  AND2_X1 _41456_ (
    .A1(\cpuregs[10] [12]),
    .A2(_22077_),
    .ZN(_07057_)
  );
  INV_X1 _41457_ (
    .A(_07057_),
    .ZN(_07058_)
  );
  AND2_X1 _41458_ (
    .A1(_07056_),
    .A2(_07058_),
    .ZN(_07059_)
  );
  INV_X1 _41459_ (
    .A(_07059_),
    .ZN(_07060_)
  );
  AND2_X1 _41460_ (
    .A1(_22152_),
    .A2(_07060_),
    .ZN(_07061_)
  );
  INV_X1 _41461_ (
    .A(_07061_),
    .ZN(_07062_)
  );
  AND2_X1 _41462_ (
    .A1(_07054_),
    .A2(_07062_),
    .ZN(_07063_)
  );
  AND2_X1 _41463_ (
    .A1(\cpuregs[9] [12]),
    .A2(_22077_),
    .ZN(_07064_)
  );
  INV_X1 _41464_ (
    .A(_07064_),
    .ZN(_07065_)
  );
  AND2_X1 _41465_ (
    .A1(\cpuregs[13] [12]),
    .A2(_00007_[2]),
    .ZN(_07066_)
  );
  INV_X1 _41466_ (
    .A(_07066_),
    .ZN(_07067_)
  );
  AND2_X1 _41467_ (
    .A1(_07065_),
    .A2(_07067_),
    .ZN(_07068_)
  );
  INV_X1 _41468_ (
    .A(_07068_),
    .ZN(_07069_)
  );
  AND2_X1 _41469_ (
    .A1(_00007_[0]),
    .A2(_07069_),
    .ZN(_07070_)
  );
  INV_X1 _41470_ (
    .A(_07070_),
    .ZN(_07071_)
  );
  AND2_X1 _41471_ (
    .A1(\cpuregs[12] [12]),
    .A2(_00007_[2]),
    .ZN(_07072_)
  );
  INV_X1 _41472_ (
    .A(_07072_),
    .ZN(_07073_)
  );
  AND2_X1 _41473_ (
    .A1(\cpuregs[8] [12]),
    .A2(_22077_),
    .ZN(_07074_)
  );
  INV_X1 _41474_ (
    .A(_07074_),
    .ZN(_07075_)
  );
  AND2_X1 _41475_ (
    .A1(_07073_),
    .A2(_07075_),
    .ZN(_07076_)
  );
  INV_X1 _41476_ (
    .A(_07076_),
    .ZN(_07077_)
  );
  AND2_X1 _41477_ (
    .A1(_22152_),
    .A2(_07077_),
    .ZN(_07078_)
  );
  INV_X1 _41478_ (
    .A(_07078_),
    .ZN(_07079_)
  );
  AND2_X1 _41479_ (
    .A1(_07071_),
    .A2(_07079_),
    .ZN(_07080_)
  );
  AND2_X1 _41480_ (
    .A1(_21445_),
    .A2(_22077_),
    .ZN(_07081_)
  );
  INV_X1 _41481_ (
    .A(_07081_),
    .ZN(_07082_)
  );
  AND2_X1 _41482_ (
    .A1(_21656_),
    .A2(_00007_[2]),
    .ZN(_07083_)
  );
  INV_X1 _41483_ (
    .A(_07083_),
    .ZN(_07084_)
  );
  AND2_X1 _41484_ (
    .A1(_07082_),
    .A2(_07084_),
    .ZN(_07085_)
  );
  AND2_X1 _41485_ (
    .A1(_21467_),
    .A2(_22077_),
    .ZN(_07086_)
  );
  INV_X1 _41486_ (
    .A(_07086_),
    .ZN(_07087_)
  );
  AND2_X1 _41487_ (
    .A1(_21766_),
    .A2(_00007_[2]),
    .ZN(_07088_)
  );
  INV_X1 _41488_ (
    .A(_07088_),
    .ZN(_07089_)
  );
  AND2_X1 _41489_ (
    .A1(_00007_[0]),
    .A2(_07089_),
    .ZN(_07090_)
  );
  AND2_X1 _41490_ (
    .A1(_07087_),
    .A2(_07090_),
    .ZN(_07091_)
  );
  INV_X1 _41491_ (
    .A(_07091_),
    .ZN(_07092_)
  );
  AND2_X1 _41492_ (
    .A1(_22152_),
    .A2(_07085_),
    .ZN(_07093_)
  );
  INV_X1 _41493_ (
    .A(_07093_),
    .ZN(_07094_)
  );
  AND2_X1 _41494_ (
    .A1(_07092_),
    .A2(_07094_),
    .ZN(_07095_)
  );
  AND2_X1 _41495_ (
    .A1(_21599_),
    .A2(_22077_),
    .ZN(_07096_)
  );
  INV_X1 _41496_ (
    .A(_07096_),
    .ZN(_07097_)
  );
  AND2_X1 _41497_ (
    .A1(_21419_),
    .A2(_00007_[2]),
    .ZN(_07098_)
  );
  INV_X1 _41498_ (
    .A(_07098_),
    .ZN(_07099_)
  );
  AND2_X1 _41499_ (
    .A1(_21379_),
    .A2(_00007_[2]),
    .ZN(_07100_)
  );
  INV_X1 _41500_ (
    .A(_07100_),
    .ZN(_07101_)
  );
  AND2_X1 _41501_ (
    .A1(_21625_),
    .A2(_22077_),
    .ZN(_07102_)
  );
  INV_X1 _41502_ (
    .A(_07102_),
    .ZN(_07103_)
  );
  AND2_X1 _41503_ (
    .A1(_22152_),
    .A2(_07099_),
    .ZN(_07104_)
  );
  AND2_X1 _41504_ (
    .A1(_07097_),
    .A2(_07104_),
    .ZN(_07105_)
  );
  INV_X1 _41505_ (
    .A(_07105_),
    .ZN(_07106_)
  );
  AND2_X1 _41506_ (
    .A1(_00007_[0]),
    .A2(_07101_),
    .ZN(_07107_)
  );
  AND2_X1 _41507_ (
    .A1(_07103_),
    .A2(_07107_),
    .ZN(_07108_)
  );
  INV_X1 _41508_ (
    .A(_07108_),
    .ZN(_07109_)
  );
  AND2_X1 _41509_ (
    .A1(_07106_),
    .A2(_07109_),
    .ZN(_07110_)
  );
  AND2_X1 _41510_ (
    .A1(_21549_),
    .A2(_22077_),
    .ZN(_07111_)
  );
  INV_X1 _41511_ (
    .A(_07111_),
    .ZN(_07112_)
  );
  AND2_X1 _41512_ (
    .A1(_21815_),
    .A2(_00007_[2]),
    .ZN(_07113_)
  );
  INV_X1 _41513_ (
    .A(_07113_),
    .ZN(_07114_)
  );
  AND2_X1 _41514_ (
    .A1(_22152_),
    .A2(_07114_),
    .ZN(_07115_)
  );
  AND2_X1 _41515_ (
    .A1(_07112_),
    .A2(_07115_),
    .ZN(_07116_)
  );
  INV_X1 _41516_ (
    .A(_07116_),
    .ZN(_07117_)
  );
  AND2_X1 _41517_ (
    .A1(\cpuregs[7] [12]),
    .A2(_00007_[2]),
    .ZN(_07118_)
  );
  INV_X1 _41518_ (
    .A(_07118_),
    .ZN(_07119_)
  );
  AND2_X1 _41519_ (
    .A1(\cpuregs[3] [12]),
    .A2(_22077_),
    .ZN(_07120_)
  );
  INV_X1 _41520_ (
    .A(_07120_),
    .ZN(_07121_)
  );
  AND2_X1 _41521_ (
    .A1(_07119_),
    .A2(_07121_),
    .ZN(_07122_)
  );
  INV_X1 _41522_ (
    .A(_07122_),
    .ZN(_07123_)
  );
  AND2_X1 _41523_ (
    .A1(_00007_[0]),
    .A2(_07123_),
    .ZN(_07124_)
  );
  INV_X1 _41524_ (
    .A(_07124_),
    .ZN(_07125_)
  );
  AND2_X1 _41525_ (
    .A1(_07117_),
    .A2(_07125_),
    .ZN(_07126_)
  );
  AND2_X1 _41526_ (
    .A1(\cpuregs[1] [12]),
    .A2(_22077_),
    .ZN(_07127_)
  );
  INV_X1 _41527_ (
    .A(_07127_),
    .ZN(_07128_)
  );
  AND2_X1 _41528_ (
    .A1(\cpuregs[5] [12]),
    .A2(_00007_[2]),
    .ZN(_07129_)
  );
  INV_X1 _41529_ (
    .A(_07129_),
    .ZN(_07130_)
  );
  AND2_X1 _41530_ (
    .A1(_07128_),
    .A2(_07130_),
    .ZN(_07131_)
  );
  INV_X1 _41531_ (
    .A(_07131_),
    .ZN(_07132_)
  );
  AND2_X1 _41532_ (
    .A1(_00007_[0]),
    .A2(_07132_),
    .ZN(_07133_)
  );
  INV_X1 _41533_ (
    .A(_07133_),
    .ZN(_07134_)
  );
  AND2_X1 _41534_ (
    .A1(\cpuregs[4] [12]),
    .A2(_00007_[2]),
    .ZN(_07135_)
  );
  INV_X1 _41535_ (
    .A(_07135_),
    .ZN(_07136_)
  );
  AND2_X1 _41536_ (
    .A1(\cpuregs[0] [12]),
    .A2(_22077_),
    .ZN(_07137_)
  );
  INV_X1 _41537_ (
    .A(_07137_),
    .ZN(_07138_)
  );
  AND2_X1 _41538_ (
    .A1(_07136_),
    .A2(_07138_),
    .ZN(_07139_)
  );
  INV_X1 _41539_ (
    .A(_07139_),
    .ZN(_07140_)
  );
  AND2_X1 _41540_ (
    .A1(_22152_),
    .A2(_07140_),
    .ZN(_07141_)
  );
  INV_X1 _41541_ (
    .A(_07141_),
    .ZN(_07142_)
  );
  AND2_X1 _41542_ (
    .A1(_07134_),
    .A2(_07142_),
    .ZN(_07143_)
  );
  AND2_X1 _41543_ (
    .A1(_00007_[1]),
    .A2(_07126_),
    .ZN(_07144_)
  );
  INV_X1 _41544_ (
    .A(_07144_),
    .ZN(_07145_)
  );
  AND2_X1 _41545_ (
    .A1(_22078_),
    .A2(_07143_),
    .ZN(_07146_)
  );
  INV_X1 _41546_ (
    .A(_07146_),
    .ZN(_07147_)
  );
  AND2_X1 _41547_ (
    .A1(_07145_),
    .A2(_07147_),
    .ZN(_07148_)
  );
  AND2_X1 _41548_ (
    .A1(_00007_[1]),
    .A2(_07110_),
    .ZN(_07149_)
  );
  INV_X1 _41549_ (
    .A(_07149_),
    .ZN(_07150_)
  );
  AND2_X1 _41550_ (
    .A1(_22078_),
    .A2(_07095_),
    .ZN(_07151_)
  );
  INV_X1 _41551_ (
    .A(_07151_),
    .ZN(_07152_)
  );
  AND2_X1 _41552_ (
    .A1(_22109_),
    .A2(_07152_),
    .ZN(_07153_)
  );
  AND2_X1 _41553_ (
    .A1(_07150_),
    .A2(_07153_),
    .ZN(_07154_)
  );
  INV_X1 _41554_ (
    .A(_07154_),
    .ZN(_07155_)
  );
  AND2_X1 _41555_ (
    .A1(_00007_[3]),
    .A2(_07046_),
    .ZN(_07156_)
  );
  INV_X1 _41556_ (
    .A(_07156_),
    .ZN(_07157_)
  );
  AND2_X1 _41557_ (
    .A1(_00007_[4]),
    .A2(_07157_),
    .ZN(_07158_)
  );
  AND2_X1 _41558_ (
    .A1(_07155_),
    .A2(_07158_),
    .ZN(_07159_)
  );
  INV_X1 _41559_ (
    .A(_07159_),
    .ZN(_07160_)
  );
  AND2_X1 _41560_ (
    .A1(_22109_),
    .A2(_07148_),
    .ZN(_07161_)
  );
  INV_X1 _41561_ (
    .A(_07161_),
    .ZN(_07162_)
  );
  AND2_X1 _41562_ (
    .A1(_00007_[1]),
    .A2(_07063_),
    .ZN(_07163_)
  );
  INV_X1 _41563_ (
    .A(_07163_),
    .ZN(_07164_)
  );
  AND2_X1 _41564_ (
    .A1(_22078_),
    .A2(_07080_),
    .ZN(_07165_)
  );
  INV_X1 _41565_ (
    .A(_07165_),
    .ZN(_07166_)
  );
  AND2_X1 _41566_ (
    .A1(_00007_[3]),
    .A2(_07166_),
    .ZN(_07167_)
  );
  AND2_X1 _41567_ (
    .A1(_07164_),
    .A2(_07167_),
    .ZN(_07168_)
  );
  INV_X1 _41568_ (
    .A(_07168_),
    .ZN(_07169_)
  );
  AND2_X1 _41569_ (
    .A1(_07162_),
    .A2(_07169_),
    .ZN(_07170_)
  );
  AND2_X1 _41570_ (
    .A1(_22144_),
    .A2(_07170_),
    .ZN(_07171_)
  );
  INV_X1 _41571_ (
    .A(_07171_),
    .ZN(_07172_)
  );
  AND2_X1 _41572_ (
    .A1(_07160_),
    .A2(_07172_),
    .ZN(_07173_)
  );
  AND2_X1 _41573_ (
    .A1(_05842_),
    .A2(_07173_),
    .ZN(_07174_)
  );
  INV_X1 _41574_ (
    .A(_07174_),
    .ZN(_07175_)
  );
  AND2_X1 _41575_ (
    .A1(_21212_),
    .A2(_04963_),
    .ZN(_07176_)
  );
  INV_X1 _41576_ (
    .A(_07176_),
    .ZN(_07177_)
  );
  AND2_X1 _41577_ (
    .A1(_04962_),
    .A2(_07175_),
    .ZN(_07178_)
  );
  AND2_X1 _41578_ (
    .A1(_07010_),
    .A2(_07178_),
    .ZN(_07179_)
  );
  INV_X1 _41579_ (
    .A(_07179_),
    .ZN(_07180_)
  );
  AND2_X1 _41580_ (
    .A1(_07177_),
    .A2(_07180_),
    .ZN(_00293_)
  );
  AND2_X1 _41581_ (
    .A1(_21600_),
    .A2(_22077_),
    .ZN(_07181_)
  );
  INV_X1 _41582_ (
    .A(_07181_),
    .ZN(_07182_)
  );
  AND2_X1 _41583_ (
    .A1(_21420_),
    .A2(_00007_[2]),
    .ZN(_07183_)
  );
  INV_X1 _41584_ (
    .A(_07183_),
    .ZN(_07184_)
  );
  AND2_X1 _41585_ (
    .A1(_21380_),
    .A2(_00007_[2]),
    .ZN(_07185_)
  );
  INV_X1 _41586_ (
    .A(_07185_),
    .ZN(_07186_)
  );
  AND2_X1 _41587_ (
    .A1(_21626_),
    .A2(_22077_),
    .ZN(_07187_)
  );
  INV_X1 _41588_ (
    .A(_07187_),
    .ZN(_07188_)
  );
  AND2_X1 _41589_ (
    .A1(\cpuregs[11] [13]),
    .A2(_22077_),
    .ZN(_07189_)
  );
  INV_X1 _41590_ (
    .A(_07189_),
    .ZN(_07190_)
  );
  AND2_X1 _41591_ (
    .A1(\cpuregs[15] [13]),
    .A2(_00007_[2]),
    .ZN(_07191_)
  );
  INV_X1 _41592_ (
    .A(_07191_),
    .ZN(_07192_)
  );
  AND2_X1 _41593_ (
    .A1(_07190_),
    .A2(_07192_),
    .ZN(_07193_)
  );
  INV_X1 _41594_ (
    .A(_07193_),
    .ZN(_07194_)
  );
  AND2_X1 _41595_ (
    .A1(_00007_[0]),
    .A2(_07194_),
    .ZN(_07195_)
  );
  INV_X1 _41596_ (
    .A(_07195_),
    .ZN(_07196_)
  );
  AND2_X1 _41597_ (
    .A1(\cpuregs[14] [13]),
    .A2(_00007_[2]),
    .ZN(_07197_)
  );
  INV_X1 _41598_ (
    .A(_07197_),
    .ZN(_07198_)
  );
  AND2_X1 _41599_ (
    .A1(\cpuregs[10] [13]),
    .A2(_22077_),
    .ZN(_07199_)
  );
  INV_X1 _41600_ (
    .A(_07199_),
    .ZN(_07200_)
  );
  AND2_X1 _41601_ (
    .A1(_07198_),
    .A2(_07200_),
    .ZN(_07201_)
  );
  INV_X1 _41602_ (
    .A(_07201_),
    .ZN(_07202_)
  );
  AND2_X1 _41603_ (
    .A1(_22152_),
    .A2(_07202_),
    .ZN(_07203_)
  );
  INV_X1 _41604_ (
    .A(_07203_),
    .ZN(_07204_)
  );
  AND2_X1 _41605_ (
    .A1(_07196_),
    .A2(_07204_),
    .ZN(_07205_)
  );
  AND2_X1 _41606_ (
    .A1(_21550_),
    .A2(_22077_),
    .ZN(_07206_)
  );
  INV_X1 _41607_ (
    .A(_07206_),
    .ZN(_07207_)
  );
  AND2_X1 _41608_ (
    .A1(_21816_),
    .A2(_00007_[2]),
    .ZN(_07208_)
  );
  INV_X1 _41609_ (
    .A(_07208_),
    .ZN(_07209_)
  );
  AND2_X1 _41610_ (
    .A1(_22152_),
    .A2(_07209_),
    .ZN(_07210_)
  );
  AND2_X1 _41611_ (
    .A1(_07207_),
    .A2(_07210_),
    .ZN(_07211_)
  );
  INV_X1 _41612_ (
    .A(_07211_),
    .ZN(_07212_)
  );
  AND2_X1 _41613_ (
    .A1(_21789_),
    .A2(_00007_[2]),
    .ZN(_07213_)
  );
  INV_X1 _41614_ (
    .A(_07213_),
    .ZN(_07214_)
  );
  AND2_X1 _41615_ (
    .A1(_21497_),
    .A2(_22077_),
    .ZN(_07215_)
  );
  INV_X1 _41616_ (
    .A(_07215_),
    .ZN(_07216_)
  );
  AND2_X1 _41617_ (
    .A1(_00007_[0]),
    .A2(_07216_),
    .ZN(_07217_)
  );
  AND2_X1 _41618_ (
    .A1(_07214_),
    .A2(_07217_),
    .ZN(_07218_)
  );
  INV_X1 _41619_ (
    .A(_07218_),
    .ZN(_07219_)
  );
  AND2_X1 _41620_ (
    .A1(_07212_),
    .A2(_07219_),
    .ZN(_07220_)
  );
  AND2_X1 _41621_ (
    .A1(_21446_),
    .A2(_22077_),
    .ZN(_07221_)
  );
  INV_X1 _41622_ (
    .A(_07221_),
    .ZN(_07222_)
  );
  AND2_X1 _41623_ (
    .A1(_21657_),
    .A2(_00007_[2]),
    .ZN(_07223_)
  );
  INV_X1 _41624_ (
    .A(_07223_),
    .ZN(_07224_)
  );
  AND2_X1 _41625_ (
    .A1(_07222_),
    .A2(_07224_),
    .ZN(_07225_)
  );
  AND2_X1 _41626_ (
    .A1(_21468_),
    .A2(_22077_),
    .ZN(_07226_)
  );
  INV_X1 _41627_ (
    .A(_07226_),
    .ZN(_07227_)
  );
  AND2_X1 _41628_ (
    .A1(_21767_),
    .A2(_00007_[2]),
    .ZN(_07228_)
  );
  INV_X1 _41629_ (
    .A(_07228_),
    .ZN(_07229_)
  );
  AND2_X1 _41630_ (
    .A1(\cpuregs[9] [13]),
    .A2(_22077_),
    .ZN(_07230_)
  );
  INV_X1 _41631_ (
    .A(_07230_),
    .ZN(_07231_)
  );
  AND2_X1 _41632_ (
    .A1(\cpuregs[13] [13]),
    .A2(_00007_[2]),
    .ZN(_07232_)
  );
  INV_X1 _41633_ (
    .A(_07232_),
    .ZN(_07233_)
  );
  AND2_X1 _41634_ (
    .A1(_07231_),
    .A2(_07233_),
    .ZN(_07234_)
  );
  INV_X1 _41635_ (
    .A(_07234_),
    .ZN(_07235_)
  );
  AND2_X1 _41636_ (
    .A1(_00007_[0]),
    .A2(_07235_),
    .ZN(_07236_)
  );
  INV_X1 _41637_ (
    .A(_07236_),
    .ZN(_07237_)
  );
  AND2_X1 _41638_ (
    .A1(\cpuregs[12] [13]),
    .A2(_00007_[2]),
    .ZN(_07238_)
  );
  INV_X1 _41639_ (
    .A(_07238_),
    .ZN(_07239_)
  );
  AND2_X1 _41640_ (
    .A1(\cpuregs[8] [13]),
    .A2(_22077_),
    .ZN(_07240_)
  );
  INV_X1 _41641_ (
    .A(_07240_),
    .ZN(_07241_)
  );
  AND2_X1 _41642_ (
    .A1(_07239_),
    .A2(_07241_),
    .ZN(_07242_)
  );
  INV_X1 _41643_ (
    .A(_07242_),
    .ZN(_07243_)
  );
  AND2_X1 _41644_ (
    .A1(_22152_),
    .A2(_07243_),
    .ZN(_07244_)
  );
  INV_X1 _41645_ (
    .A(_07244_),
    .ZN(_07245_)
  );
  AND2_X1 _41646_ (
    .A1(_07237_),
    .A2(_07245_),
    .ZN(_07246_)
  );
  AND2_X1 _41647_ (
    .A1(_21679_),
    .A2(_00007_[2]),
    .ZN(_07247_)
  );
  INV_X1 _41648_ (
    .A(_07247_),
    .ZN(_07248_)
  );
  AND2_X1 _41649_ (
    .A1(_21963_),
    .A2(_22077_),
    .ZN(_07249_)
  );
  INV_X1 _41650_ (
    .A(_07249_),
    .ZN(_07250_)
  );
  AND2_X1 _41651_ (
    .A1(_07248_),
    .A2(_07250_),
    .ZN(_07251_)
  );
  AND2_X1 _41652_ (
    .A1(_22152_),
    .A2(_07251_),
    .ZN(_07252_)
  );
  INV_X1 _41653_ (
    .A(_07252_),
    .ZN(_07253_)
  );
  AND2_X1 _41654_ (
    .A1(_21522_),
    .A2(_22077_),
    .ZN(_07254_)
  );
  INV_X1 _41655_ (
    .A(_07254_),
    .ZN(_07255_)
  );
  AND2_X1 _41656_ (
    .A1(_21742_),
    .A2(_00007_[2]),
    .ZN(_07256_)
  );
  INV_X1 _41657_ (
    .A(_07256_),
    .ZN(_07257_)
  );
  AND2_X1 _41658_ (
    .A1(_00007_[0]),
    .A2(_07257_),
    .ZN(_07258_)
  );
  AND2_X1 _41659_ (
    .A1(_07255_),
    .A2(_07258_),
    .ZN(_07259_)
  );
  INV_X1 _41660_ (
    .A(_07259_),
    .ZN(_07260_)
  );
  AND2_X1 _41661_ (
    .A1(_07253_),
    .A2(_07260_),
    .ZN(_07261_)
  );
  AND2_X1 _41662_ (
    .A1(_22152_),
    .A2(_07184_),
    .ZN(_07262_)
  );
  AND2_X1 _41663_ (
    .A1(_07182_),
    .A2(_07262_),
    .ZN(_07263_)
  );
  INV_X1 _41664_ (
    .A(_07263_),
    .ZN(_07264_)
  );
  AND2_X1 _41665_ (
    .A1(_00007_[0]),
    .A2(_07186_),
    .ZN(_07265_)
  );
  AND2_X1 _41666_ (
    .A1(_07188_),
    .A2(_07265_),
    .ZN(_07266_)
  );
  INV_X1 _41667_ (
    .A(_07266_),
    .ZN(_07267_)
  );
  AND2_X1 _41668_ (
    .A1(_07264_),
    .A2(_07267_),
    .ZN(_07268_)
  );
  AND2_X1 _41669_ (
    .A1(_00007_[1]),
    .A2(_07268_),
    .ZN(_07269_)
  );
  INV_X1 _41670_ (
    .A(_07269_),
    .ZN(_07270_)
  );
  AND2_X1 _41671_ (
    .A1(_00007_[0]),
    .A2(_07229_),
    .ZN(_07271_)
  );
  AND2_X1 _41672_ (
    .A1(_07227_),
    .A2(_07271_),
    .ZN(_07272_)
  );
  INV_X1 _41673_ (
    .A(_07272_),
    .ZN(_07273_)
  );
  AND2_X1 _41674_ (
    .A1(_22152_),
    .A2(_07225_),
    .ZN(_07274_)
  );
  INV_X1 _41675_ (
    .A(_07274_),
    .ZN(_07275_)
  );
  AND2_X1 _41676_ (
    .A1(_07273_),
    .A2(_07275_),
    .ZN(_07276_)
  );
  AND2_X1 _41677_ (
    .A1(_22078_),
    .A2(_07276_),
    .ZN(_07277_)
  );
  INV_X1 _41678_ (
    .A(_07277_),
    .ZN(_07278_)
  );
  AND2_X1 _41679_ (
    .A1(_22109_),
    .A2(_07278_),
    .ZN(_07279_)
  );
  AND2_X1 _41680_ (
    .A1(_07270_),
    .A2(_07279_),
    .ZN(_07280_)
  );
  INV_X1 _41681_ (
    .A(_07280_),
    .ZN(_07281_)
  );
  AND2_X1 _41682_ (
    .A1(_21928_),
    .A2(_22077_),
    .ZN(_07282_)
  );
  INV_X1 _41683_ (
    .A(_07282_),
    .ZN(_07283_)
  );
  AND2_X1 _41684_ (
    .A1(_21944_),
    .A2(_00007_[2]),
    .ZN(_07284_)
  );
  INV_X1 _41685_ (
    .A(_07284_),
    .ZN(_07285_)
  );
  AND2_X1 _41686_ (
    .A1(_00007_[0]),
    .A2(_07285_),
    .ZN(_07286_)
  );
  AND2_X1 _41687_ (
    .A1(_07283_),
    .A2(_07286_),
    .ZN(_07287_)
  );
  INV_X1 _41688_ (
    .A(_07287_),
    .ZN(_07288_)
  );
  AND2_X1 _41689_ (
    .A1(_21876_),
    .A2(_22077_),
    .ZN(_07289_)
  );
  INV_X1 _41690_ (
    .A(_07289_),
    .ZN(_07290_)
  );
  AND2_X1 _41691_ (
    .A1(_21856_),
    .A2(_00007_[2]),
    .ZN(_07291_)
  );
  INV_X1 _41692_ (
    .A(_07291_),
    .ZN(_07292_)
  );
  AND2_X1 _41693_ (
    .A1(_07290_),
    .A2(_07292_),
    .ZN(_07293_)
  );
  AND2_X1 _41694_ (
    .A1(_22152_),
    .A2(_07293_),
    .ZN(_07294_)
  );
  INV_X1 _41695_ (
    .A(_07294_),
    .ZN(_07295_)
  );
  AND2_X1 _41696_ (
    .A1(_07288_),
    .A2(_07295_),
    .ZN(_07296_)
  );
  AND2_X1 _41697_ (
    .A1(_00007_[1]),
    .A2(_07296_),
    .ZN(_07297_)
  );
  INV_X1 _41698_ (
    .A(_07297_),
    .ZN(_07298_)
  );
  AND2_X1 _41699_ (
    .A1(_21840_),
    .A2(_22077_),
    .ZN(_07299_)
  );
  INV_X1 _41700_ (
    .A(_07299_),
    .ZN(_07300_)
  );
  AND2_X1 _41701_ (
    .A1(_21896_),
    .A2(_00007_[2]),
    .ZN(_07301_)
  );
  INV_X1 _41702_ (
    .A(_07301_),
    .ZN(_07302_)
  );
  AND2_X1 _41703_ (
    .A1(_00007_[0]),
    .A2(_07302_),
    .ZN(_07303_)
  );
  AND2_X1 _41704_ (
    .A1(_07300_),
    .A2(_07303_),
    .ZN(_07304_)
  );
  INV_X1 _41705_ (
    .A(_07304_),
    .ZN(_07305_)
  );
  AND2_X1 _41706_ (
    .A1(_21574_),
    .A2(_22077_),
    .ZN(_07306_)
  );
  INV_X1 _41707_ (
    .A(_07306_),
    .ZN(_07307_)
  );
  AND2_X1 _41708_ (
    .A1(_21912_),
    .A2(_00007_[2]),
    .ZN(_07308_)
  );
  INV_X1 _41709_ (
    .A(_07308_),
    .ZN(_07309_)
  );
  AND2_X1 _41710_ (
    .A1(_07307_),
    .A2(_07309_),
    .ZN(_07310_)
  );
  AND2_X1 _41711_ (
    .A1(_22152_),
    .A2(_07310_),
    .ZN(_07311_)
  );
  INV_X1 _41712_ (
    .A(_07311_),
    .ZN(_07312_)
  );
  AND2_X1 _41713_ (
    .A1(_07305_),
    .A2(_07312_),
    .ZN(_07313_)
  );
  AND2_X1 _41714_ (
    .A1(_22078_),
    .A2(_07313_),
    .ZN(_07314_)
  );
  INV_X1 _41715_ (
    .A(_07314_),
    .ZN(_07315_)
  );
  AND2_X1 _41716_ (
    .A1(_00007_[3]),
    .A2(_07315_),
    .ZN(_07316_)
  );
  AND2_X1 _41717_ (
    .A1(_07298_),
    .A2(_07316_),
    .ZN(_07317_)
  );
  INV_X1 _41718_ (
    .A(_07317_),
    .ZN(_07318_)
  );
  AND2_X1 _41719_ (
    .A1(_00007_[4]),
    .A2(_07318_),
    .ZN(_07319_)
  );
  AND2_X1 _41720_ (
    .A1(_07281_),
    .A2(_07319_),
    .ZN(_07320_)
  );
  INV_X1 _41721_ (
    .A(_07320_),
    .ZN(_07321_)
  );
  AND2_X1 _41722_ (
    .A1(_00007_[1]),
    .A2(_07220_),
    .ZN(_07322_)
  );
  INV_X1 _41723_ (
    .A(_07322_),
    .ZN(_07323_)
  );
  AND2_X1 _41724_ (
    .A1(_22078_),
    .A2(_07261_),
    .ZN(_07324_)
  );
  INV_X1 _41725_ (
    .A(_07324_),
    .ZN(_07325_)
  );
  AND2_X1 _41726_ (
    .A1(_22109_),
    .A2(_07325_),
    .ZN(_07326_)
  );
  AND2_X1 _41727_ (
    .A1(_07323_),
    .A2(_07326_),
    .ZN(_07327_)
  );
  INV_X1 _41728_ (
    .A(_07327_),
    .ZN(_07328_)
  );
  AND2_X1 _41729_ (
    .A1(_00007_[1]),
    .A2(_07205_),
    .ZN(_07329_)
  );
  INV_X1 _41730_ (
    .A(_07329_),
    .ZN(_07330_)
  );
  AND2_X1 _41731_ (
    .A1(_22078_),
    .A2(_07246_),
    .ZN(_07331_)
  );
  INV_X1 _41732_ (
    .A(_07331_),
    .ZN(_07332_)
  );
  AND2_X1 _41733_ (
    .A1(_00007_[3]),
    .A2(_07332_),
    .ZN(_07333_)
  );
  AND2_X1 _41734_ (
    .A1(_07330_),
    .A2(_07333_),
    .ZN(_07334_)
  );
  INV_X1 _41735_ (
    .A(_07334_),
    .ZN(_07335_)
  );
  AND2_X1 _41736_ (
    .A1(_07328_),
    .A2(_07335_),
    .ZN(_07336_)
  );
  AND2_X1 _41737_ (
    .A1(_22144_),
    .A2(_07336_),
    .ZN(_07337_)
  );
  INV_X1 _41738_ (
    .A(_07337_),
    .ZN(_07338_)
  );
  AND2_X1 _41739_ (
    .A1(_07321_),
    .A2(_07338_),
    .ZN(_07339_)
  );
  AND2_X1 _41740_ (
    .A1(_05842_),
    .A2(_07339_),
    .ZN(_07340_)
  );
  INV_X1 _41741_ (
    .A(_07340_),
    .ZN(_07341_)
  );
  AND2_X1 _41742_ (
    .A1(decoded_imm[13]),
    .A2(_04966_),
    .ZN(_07342_)
  );
  INV_X1 _41743_ (
    .A(_07342_),
    .ZN(_07343_)
  );
  AND2_X1 _41744_ (
    .A1(_21213_),
    .A2(_04963_),
    .ZN(_07344_)
  );
  INV_X1 _41745_ (
    .A(_07344_),
    .ZN(_07345_)
  );
  AND2_X1 _41746_ (
    .A1(_04962_),
    .A2(_07343_),
    .ZN(_07346_)
  );
  AND2_X1 _41747_ (
    .A1(_07341_),
    .A2(_07346_),
    .ZN(_07347_)
  );
  INV_X1 _41748_ (
    .A(_07347_),
    .ZN(_07348_)
  );
  AND2_X1 _41749_ (
    .A1(_07345_),
    .A2(_07348_),
    .ZN(_00294_)
  );
  AND2_X1 _41750_ (
    .A1(decoded_imm[14]),
    .A2(_04966_),
    .ZN(_07349_)
  );
  INV_X1 _41751_ (
    .A(_07349_),
    .ZN(_07350_)
  );
  AND2_X1 _41752_ (
    .A1(\cpuregs[19] [14]),
    .A2(_22077_),
    .ZN(_07351_)
  );
  INV_X1 _41753_ (
    .A(_07351_),
    .ZN(_07352_)
  );
  AND2_X1 _41754_ (
    .A1(\cpuregs[23] [14]),
    .A2(_00007_[2]),
    .ZN(_07353_)
  );
  INV_X1 _41755_ (
    .A(_07353_),
    .ZN(_07354_)
  );
  AND2_X1 _41756_ (
    .A1(_07352_),
    .A2(_07354_),
    .ZN(_07355_)
  );
  INV_X1 _41757_ (
    .A(_07355_),
    .ZN(_07356_)
  );
  AND2_X1 _41758_ (
    .A1(_00007_[0]),
    .A2(_07356_),
    .ZN(_07357_)
  );
  INV_X1 _41759_ (
    .A(_07357_),
    .ZN(_07358_)
  );
  AND2_X1 _41760_ (
    .A1(_21601_),
    .A2(_22077_),
    .ZN(_07359_)
  );
  INV_X1 _41761_ (
    .A(_07359_),
    .ZN(_07360_)
  );
  AND2_X1 _41762_ (
    .A1(_21421_),
    .A2(_00007_[2]),
    .ZN(_07361_)
  );
  INV_X1 _41763_ (
    .A(_07361_),
    .ZN(_07362_)
  );
  AND2_X1 _41764_ (
    .A1(_22152_),
    .A2(_07362_),
    .ZN(_07363_)
  );
  AND2_X1 _41765_ (
    .A1(_07360_),
    .A2(_07363_),
    .ZN(_07364_)
  );
  INV_X1 _41766_ (
    .A(_07364_),
    .ZN(_07365_)
  );
  AND2_X1 _41767_ (
    .A1(_21498_),
    .A2(_22077_),
    .ZN(_07366_)
  );
  INV_X1 _41768_ (
    .A(_07366_),
    .ZN(_07367_)
  );
  AND2_X1 _41769_ (
    .A1(_21790_),
    .A2(_00007_[2]),
    .ZN(_07368_)
  );
  INV_X1 _41770_ (
    .A(_07368_),
    .ZN(_07369_)
  );
  AND2_X1 _41771_ (
    .A1(_00007_[0]),
    .A2(_07369_),
    .ZN(_07370_)
  );
  AND2_X1 _41772_ (
    .A1(_07367_),
    .A2(_07370_),
    .ZN(_07371_)
  );
  INV_X1 _41773_ (
    .A(_07371_),
    .ZN(_07372_)
  );
  AND2_X1 _41774_ (
    .A1(_21817_),
    .A2(_00007_[2]),
    .ZN(_07373_)
  );
  INV_X1 _41775_ (
    .A(_07373_),
    .ZN(_07374_)
  );
  AND2_X1 _41776_ (
    .A1(_21551_),
    .A2(_22077_),
    .ZN(_07375_)
  );
  INV_X1 _41777_ (
    .A(_07375_),
    .ZN(_07376_)
  );
  AND2_X1 _41778_ (
    .A1(_22152_),
    .A2(_07376_),
    .ZN(_07377_)
  );
  AND2_X1 _41779_ (
    .A1(_07374_),
    .A2(_07377_),
    .ZN(_07378_)
  );
  INV_X1 _41780_ (
    .A(_07378_),
    .ZN(_07379_)
  );
  AND2_X1 _41781_ (
    .A1(\cpuregs[17] [14]),
    .A2(_22077_),
    .ZN(_07380_)
  );
  INV_X1 _41782_ (
    .A(_07380_),
    .ZN(_07381_)
  );
  AND2_X1 _41783_ (
    .A1(\cpuregs[21] [14]),
    .A2(_00007_[2]),
    .ZN(_07382_)
  );
  INV_X1 _41784_ (
    .A(_07382_),
    .ZN(_07383_)
  );
  AND2_X1 _41785_ (
    .A1(_07381_),
    .A2(_07383_),
    .ZN(_07384_)
  );
  INV_X1 _41786_ (
    .A(_07384_),
    .ZN(_07385_)
  );
  AND2_X1 _41787_ (
    .A1(_00007_[0]),
    .A2(_07385_),
    .ZN(_07386_)
  );
  INV_X1 _41788_ (
    .A(_07386_),
    .ZN(_07387_)
  );
  AND2_X1 _41789_ (
    .A1(\cpuregs[16] [14]),
    .A2(_22077_),
    .ZN(_07388_)
  );
  INV_X1 _41790_ (
    .A(_07388_),
    .ZN(_07389_)
  );
  AND2_X1 _41791_ (
    .A1(\cpuregs[20] [14]),
    .A2(_00007_[2]),
    .ZN(_07390_)
  );
  INV_X1 _41792_ (
    .A(_07390_),
    .ZN(_07391_)
  );
  AND2_X1 _41793_ (
    .A1(_07389_),
    .A2(_07391_),
    .ZN(_07392_)
  );
  INV_X1 _41794_ (
    .A(_07392_),
    .ZN(_07393_)
  );
  AND2_X1 _41795_ (
    .A1(_22152_),
    .A2(_07393_),
    .ZN(_07394_)
  );
  INV_X1 _41796_ (
    .A(_07394_),
    .ZN(_07395_)
  );
  AND2_X1 _41797_ (
    .A1(_07387_),
    .A2(_07395_),
    .ZN(_07396_)
  );
  AND2_X1 _41798_ (
    .A1(_21523_),
    .A2(_22077_),
    .ZN(_07397_)
  );
  INV_X1 _41799_ (
    .A(_07397_),
    .ZN(_07398_)
  );
  AND2_X1 _41800_ (
    .A1(_21743_),
    .A2(_00007_[2]),
    .ZN(_07399_)
  );
  INV_X1 _41801_ (
    .A(_07399_),
    .ZN(_07400_)
  );
  AND2_X1 _41802_ (
    .A1(_00007_[0]),
    .A2(_07400_),
    .ZN(_07401_)
  );
  AND2_X1 _41803_ (
    .A1(_07398_),
    .A2(_07401_),
    .ZN(_07402_)
  );
  INV_X1 _41804_ (
    .A(_07402_),
    .ZN(_07403_)
  );
  AND2_X1 _41805_ (
    .A1(_21964_),
    .A2(_22077_),
    .ZN(_07404_)
  );
  INV_X1 _41806_ (
    .A(_07404_),
    .ZN(_07405_)
  );
  AND2_X1 _41807_ (
    .A1(_21680_),
    .A2(_00007_[2]),
    .ZN(_07406_)
  );
  INV_X1 _41808_ (
    .A(_07406_),
    .ZN(_07407_)
  );
  AND2_X1 _41809_ (
    .A1(_07405_),
    .A2(_07407_),
    .ZN(_07408_)
  );
  AND2_X1 _41810_ (
    .A1(_22152_),
    .A2(_07408_),
    .ZN(_07409_)
  );
  INV_X1 _41811_ (
    .A(_07409_),
    .ZN(_07410_)
  );
  AND2_X1 _41812_ (
    .A1(_07403_),
    .A2(_07410_),
    .ZN(_07411_)
  );
  AND2_X1 _41813_ (
    .A1(_22078_),
    .A2(_07411_),
    .ZN(_07412_)
  );
  INV_X1 _41814_ (
    .A(_07412_),
    .ZN(_07413_)
  );
  AND2_X1 _41815_ (
    .A1(_00007_[1]),
    .A2(_07379_),
    .ZN(_07414_)
  );
  AND2_X1 _41816_ (
    .A1(_07372_),
    .A2(_07414_),
    .ZN(_07415_)
  );
  INV_X1 _41817_ (
    .A(_07415_),
    .ZN(_07416_)
  );
  AND2_X1 _41818_ (
    .A1(_07413_),
    .A2(_07416_),
    .ZN(_07417_)
  );
  AND2_X1 _41819_ (
    .A1(_22144_),
    .A2(_07417_),
    .ZN(_07418_)
  );
  INV_X1 _41820_ (
    .A(_07418_),
    .ZN(_07419_)
  );
  AND2_X1 _41821_ (
    .A1(_00007_[1]),
    .A2(_07365_),
    .ZN(_07420_)
  );
  AND2_X1 _41822_ (
    .A1(_07358_),
    .A2(_07420_),
    .ZN(_07421_)
  );
  INV_X1 _41823_ (
    .A(_07421_),
    .ZN(_07422_)
  );
  AND2_X1 _41824_ (
    .A1(_22078_),
    .A2(_07396_),
    .ZN(_07423_)
  );
  INV_X1 _41825_ (
    .A(_07423_),
    .ZN(_07424_)
  );
  AND2_X1 _41826_ (
    .A1(_07422_),
    .A2(_07424_),
    .ZN(_07425_)
  );
  AND2_X1 _41827_ (
    .A1(_00007_[4]),
    .A2(_07425_),
    .ZN(_07426_)
  );
  INV_X1 _41828_ (
    .A(_07426_),
    .ZN(_07427_)
  );
  AND2_X1 _41829_ (
    .A1(_07419_),
    .A2(_07427_),
    .ZN(_07428_)
  );
  AND2_X1 _41830_ (
    .A1(\cpuregs[26] [14]),
    .A2(_22077_),
    .ZN(_07429_)
  );
  INV_X1 _41831_ (
    .A(_07429_),
    .ZN(_07430_)
  );
  AND2_X1 _41832_ (
    .A1(\cpuregs[30] [14]),
    .A2(_00007_[2]),
    .ZN(_07431_)
  );
  INV_X1 _41833_ (
    .A(_07431_),
    .ZN(_07432_)
  );
  AND2_X1 _41834_ (
    .A1(_00007_[1]),
    .A2(_07432_),
    .ZN(_07433_)
  );
  AND2_X1 _41835_ (
    .A1(_07430_),
    .A2(_07433_),
    .ZN(_07434_)
  );
  INV_X1 _41836_ (
    .A(_07434_),
    .ZN(_07435_)
  );
  AND2_X1 _41837_ (
    .A1(\cpuregs[28] [14]),
    .A2(_00007_[2]),
    .ZN(_07436_)
  );
  INV_X1 _41838_ (
    .A(_07436_),
    .ZN(_07437_)
  );
  AND2_X1 _41839_ (
    .A1(\cpuregs[24] [14]),
    .A2(_22077_),
    .ZN(_07438_)
  );
  INV_X1 _41840_ (
    .A(_07438_),
    .ZN(_07439_)
  );
  AND2_X1 _41841_ (
    .A1(_22078_),
    .A2(_07439_),
    .ZN(_07440_)
  );
  AND2_X1 _41842_ (
    .A1(_07437_),
    .A2(_07440_),
    .ZN(_07441_)
  );
  INV_X1 _41843_ (
    .A(_07441_),
    .ZN(_07442_)
  );
  AND2_X1 _41844_ (
    .A1(_22152_),
    .A2(_07442_),
    .ZN(_07443_)
  );
  AND2_X1 _41845_ (
    .A1(_07435_),
    .A2(_07443_),
    .ZN(_07444_)
  );
  INV_X1 _41846_ (
    .A(_07444_),
    .ZN(_07445_)
  );
  AND2_X1 _41847_ (
    .A1(\cpuregs[27] [14]),
    .A2(_22077_),
    .ZN(_07446_)
  );
  INV_X1 _41848_ (
    .A(_07446_),
    .ZN(_07447_)
  );
  AND2_X1 _41849_ (
    .A1(\cpuregs[31] [14]),
    .A2(_00007_[2]),
    .ZN(_07448_)
  );
  INV_X1 _41850_ (
    .A(_07448_),
    .ZN(_07449_)
  );
  AND2_X1 _41851_ (
    .A1(_00007_[1]),
    .A2(_07449_),
    .ZN(_07450_)
  );
  AND2_X1 _41852_ (
    .A1(_07447_),
    .A2(_07450_),
    .ZN(_07451_)
  );
  INV_X1 _41853_ (
    .A(_07451_),
    .ZN(_07452_)
  );
  AND2_X1 _41854_ (
    .A1(\cpuregs[29] [14]),
    .A2(_00007_[2]),
    .ZN(_07453_)
  );
  INV_X1 _41855_ (
    .A(_07453_),
    .ZN(_07454_)
  );
  AND2_X1 _41856_ (
    .A1(\cpuregs[25] [14]),
    .A2(_22077_),
    .ZN(_07455_)
  );
  INV_X1 _41857_ (
    .A(_07455_),
    .ZN(_07456_)
  );
  AND2_X1 _41858_ (
    .A1(_22078_),
    .A2(_07456_),
    .ZN(_07457_)
  );
  AND2_X1 _41859_ (
    .A1(_07454_),
    .A2(_07457_),
    .ZN(_07458_)
  );
  INV_X1 _41860_ (
    .A(_07458_),
    .ZN(_07459_)
  );
  AND2_X1 _41861_ (
    .A1(_00007_[0]),
    .A2(_07459_),
    .ZN(_07460_)
  );
  AND2_X1 _41862_ (
    .A1(_07452_),
    .A2(_07460_),
    .ZN(_07461_)
  );
  INV_X1 _41863_ (
    .A(_07461_),
    .ZN(_07462_)
  );
  AND2_X1 _41864_ (
    .A1(_07445_),
    .A2(_07462_),
    .ZN(_07463_)
  );
  INV_X1 _41865_ (
    .A(_07463_),
    .ZN(_07464_)
  );
  AND2_X1 _41866_ (
    .A1(_00007_[4]),
    .A2(_07464_),
    .ZN(_07465_)
  );
  INV_X1 _41867_ (
    .A(_07465_),
    .ZN(_07466_)
  );
  AND2_X1 _41868_ (
    .A1(\cpuregs[12] [14]),
    .A2(_22078_),
    .ZN(_07467_)
  );
  INV_X1 _41869_ (
    .A(_07467_),
    .ZN(_07468_)
  );
  AND2_X1 _41870_ (
    .A1(\cpuregs[14] [14]),
    .A2(_00007_[1]),
    .ZN(_07469_)
  );
  INV_X1 _41871_ (
    .A(_07469_),
    .ZN(_07470_)
  );
  AND2_X1 _41872_ (
    .A1(_00007_[2]),
    .A2(_07470_),
    .ZN(_07471_)
  );
  AND2_X1 _41873_ (
    .A1(_07468_),
    .A2(_07471_),
    .ZN(_07472_)
  );
  INV_X1 _41874_ (
    .A(_07472_),
    .ZN(_07473_)
  );
  AND2_X1 _41875_ (
    .A1(\cpuregs[8] [14]),
    .A2(_22078_),
    .ZN(_07474_)
  );
  INV_X1 _41876_ (
    .A(_07474_),
    .ZN(_07475_)
  );
  AND2_X1 _41877_ (
    .A1(\cpuregs[10] [14]),
    .A2(_00007_[1]),
    .ZN(_07476_)
  );
  INV_X1 _41878_ (
    .A(_07476_),
    .ZN(_07477_)
  );
  AND2_X1 _41879_ (
    .A1(_22077_),
    .A2(_07477_),
    .ZN(_07478_)
  );
  AND2_X1 _41880_ (
    .A1(_07475_),
    .A2(_07478_),
    .ZN(_07479_)
  );
  INV_X1 _41881_ (
    .A(_07479_),
    .ZN(_07480_)
  );
  AND2_X1 _41882_ (
    .A1(_22152_),
    .A2(_07480_),
    .ZN(_07481_)
  );
  AND2_X1 _41883_ (
    .A1(_07473_),
    .A2(_07481_),
    .ZN(_07482_)
  );
  INV_X1 _41884_ (
    .A(_07482_),
    .ZN(_07483_)
  );
  AND2_X1 _41885_ (
    .A1(\cpuregs[13] [14]),
    .A2(_22078_),
    .ZN(_07484_)
  );
  INV_X1 _41886_ (
    .A(_07484_),
    .ZN(_07485_)
  );
  AND2_X1 _41887_ (
    .A1(\cpuregs[15] [14]),
    .A2(_00007_[1]),
    .ZN(_07486_)
  );
  INV_X1 _41888_ (
    .A(_07486_),
    .ZN(_07487_)
  );
  AND2_X1 _41889_ (
    .A1(_00007_[2]),
    .A2(_07487_),
    .ZN(_07488_)
  );
  AND2_X1 _41890_ (
    .A1(_07485_),
    .A2(_07488_),
    .ZN(_07489_)
  );
  INV_X1 _41891_ (
    .A(_07489_),
    .ZN(_07490_)
  );
  AND2_X1 _41892_ (
    .A1(\cpuregs[9] [14]),
    .A2(_22078_),
    .ZN(_07491_)
  );
  INV_X1 _41893_ (
    .A(_07491_),
    .ZN(_07492_)
  );
  AND2_X1 _41894_ (
    .A1(\cpuregs[11] [14]),
    .A2(_00007_[1]),
    .ZN(_07493_)
  );
  INV_X1 _41895_ (
    .A(_07493_),
    .ZN(_07494_)
  );
  AND2_X1 _41896_ (
    .A1(_22077_),
    .A2(_07494_),
    .ZN(_07495_)
  );
  AND2_X1 _41897_ (
    .A1(_07492_),
    .A2(_07495_),
    .ZN(_07496_)
  );
  INV_X1 _41898_ (
    .A(_07496_),
    .ZN(_07497_)
  );
  AND2_X1 _41899_ (
    .A1(_00007_[0]),
    .A2(_07497_),
    .ZN(_07498_)
  );
  AND2_X1 _41900_ (
    .A1(_07490_),
    .A2(_07498_),
    .ZN(_07499_)
  );
  INV_X1 _41901_ (
    .A(_07499_),
    .ZN(_07500_)
  );
  AND2_X1 _41902_ (
    .A1(_07483_),
    .A2(_07500_),
    .ZN(_07501_)
  );
  INV_X1 _41903_ (
    .A(_07501_),
    .ZN(_07502_)
  );
  AND2_X1 _41904_ (
    .A1(_22144_),
    .A2(_07502_),
    .ZN(_07503_)
  );
  INV_X1 _41905_ (
    .A(_07503_),
    .ZN(_07504_)
  );
  AND2_X1 _41906_ (
    .A1(_00007_[3]),
    .A2(_07504_),
    .ZN(_07505_)
  );
  AND2_X1 _41907_ (
    .A1(_07466_),
    .A2(_07505_),
    .ZN(_07506_)
  );
  INV_X1 _41908_ (
    .A(_07506_),
    .ZN(_07507_)
  );
  AND2_X1 _41909_ (
    .A1(_22109_),
    .A2(_07428_),
    .ZN(_07508_)
  );
  INV_X1 _41910_ (
    .A(_07508_),
    .ZN(_07509_)
  );
  AND2_X1 _41911_ (
    .A1(_07507_),
    .A2(_07509_),
    .ZN(_07510_)
  );
  AND2_X1 _41912_ (
    .A1(_05842_),
    .A2(_07510_),
    .ZN(_07511_)
  );
  INV_X1 _41913_ (
    .A(_07511_),
    .ZN(_07512_)
  );
  AND2_X1 _41914_ (
    .A1(_21214_),
    .A2(_04963_),
    .ZN(_07513_)
  );
  INV_X1 _41915_ (
    .A(_07513_),
    .ZN(_07514_)
  );
  AND2_X1 _41916_ (
    .A1(_04962_),
    .A2(_07512_),
    .ZN(_07515_)
  );
  AND2_X1 _41917_ (
    .A1(_07350_),
    .A2(_07515_),
    .ZN(_07516_)
  );
  INV_X1 _41918_ (
    .A(_07516_),
    .ZN(_07517_)
  );
  AND2_X1 _41919_ (
    .A1(_07514_),
    .A2(_07517_),
    .ZN(_00295_)
  );
  AND2_X1 _41920_ (
    .A1(decoded_imm[15]),
    .A2(_04966_),
    .ZN(_07518_)
  );
  INV_X1 _41921_ (
    .A(_07518_),
    .ZN(_07519_)
  );
  AND2_X1 _41922_ (
    .A1(_21602_),
    .A2(_22077_),
    .ZN(_07520_)
  );
  INV_X1 _41923_ (
    .A(_07520_),
    .ZN(_07521_)
  );
  AND2_X1 _41924_ (
    .A1(_21422_),
    .A2(_00007_[2]),
    .ZN(_07522_)
  );
  INV_X1 _41925_ (
    .A(_07522_),
    .ZN(_07523_)
  );
  AND2_X1 _41926_ (
    .A1(_21381_),
    .A2(_00007_[2]),
    .ZN(_07524_)
  );
  INV_X1 _41927_ (
    .A(_07524_),
    .ZN(_07525_)
  );
  AND2_X1 _41928_ (
    .A1(_21627_),
    .A2(_22077_),
    .ZN(_07526_)
  );
  INV_X1 _41929_ (
    .A(_07526_),
    .ZN(_07527_)
  );
  AND2_X1 _41930_ (
    .A1(\cpuregs[11] [15]),
    .A2(_22077_),
    .ZN(_07528_)
  );
  INV_X1 _41931_ (
    .A(_07528_),
    .ZN(_07529_)
  );
  AND2_X1 _41932_ (
    .A1(\cpuregs[15] [15]),
    .A2(_00007_[2]),
    .ZN(_07530_)
  );
  INV_X1 _41933_ (
    .A(_07530_),
    .ZN(_07531_)
  );
  AND2_X1 _41934_ (
    .A1(_07529_),
    .A2(_07531_),
    .ZN(_07532_)
  );
  INV_X1 _41935_ (
    .A(_07532_),
    .ZN(_07533_)
  );
  AND2_X1 _41936_ (
    .A1(_00007_[0]),
    .A2(_07533_),
    .ZN(_07534_)
  );
  INV_X1 _41937_ (
    .A(_07534_),
    .ZN(_07535_)
  );
  AND2_X1 _41938_ (
    .A1(\cpuregs[14] [15]),
    .A2(_00007_[2]),
    .ZN(_07536_)
  );
  INV_X1 _41939_ (
    .A(_07536_),
    .ZN(_07537_)
  );
  AND2_X1 _41940_ (
    .A1(\cpuregs[10] [15]),
    .A2(_22077_),
    .ZN(_07538_)
  );
  INV_X1 _41941_ (
    .A(_07538_),
    .ZN(_07539_)
  );
  AND2_X1 _41942_ (
    .A1(_07537_),
    .A2(_07539_),
    .ZN(_07540_)
  );
  INV_X1 _41943_ (
    .A(_07540_),
    .ZN(_07541_)
  );
  AND2_X1 _41944_ (
    .A1(_22152_),
    .A2(_07541_),
    .ZN(_07542_)
  );
  INV_X1 _41945_ (
    .A(_07542_),
    .ZN(_07543_)
  );
  AND2_X1 _41946_ (
    .A1(_07535_),
    .A2(_07543_),
    .ZN(_07544_)
  );
  AND2_X1 _41947_ (
    .A1(_21552_),
    .A2(_22077_),
    .ZN(_07545_)
  );
  INV_X1 _41948_ (
    .A(_07545_),
    .ZN(_07546_)
  );
  AND2_X1 _41949_ (
    .A1(_21818_),
    .A2(_00007_[2]),
    .ZN(_07547_)
  );
  INV_X1 _41950_ (
    .A(_07547_),
    .ZN(_07548_)
  );
  AND2_X1 _41951_ (
    .A1(_22152_),
    .A2(_07548_),
    .ZN(_07549_)
  );
  AND2_X1 _41952_ (
    .A1(_07546_),
    .A2(_07549_),
    .ZN(_07550_)
  );
  INV_X1 _41953_ (
    .A(_07550_),
    .ZN(_07551_)
  );
  AND2_X1 _41954_ (
    .A1(_21791_),
    .A2(_00007_[2]),
    .ZN(_07552_)
  );
  INV_X1 _41955_ (
    .A(_07552_),
    .ZN(_07553_)
  );
  AND2_X1 _41956_ (
    .A1(_21499_),
    .A2(_22077_),
    .ZN(_07554_)
  );
  INV_X1 _41957_ (
    .A(_07554_),
    .ZN(_07555_)
  );
  AND2_X1 _41958_ (
    .A1(_00007_[0]),
    .A2(_07555_),
    .ZN(_07556_)
  );
  AND2_X1 _41959_ (
    .A1(_07553_),
    .A2(_07556_),
    .ZN(_07557_)
  );
  INV_X1 _41960_ (
    .A(_07557_),
    .ZN(_07558_)
  );
  AND2_X1 _41961_ (
    .A1(_07551_),
    .A2(_07558_),
    .ZN(_07559_)
  );
  AND2_X1 _41962_ (
    .A1(_21447_),
    .A2(_22077_),
    .ZN(_07560_)
  );
  INV_X1 _41963_ (
    .A(_07560_),
    .ZN(_07561_)
  );
  AND2_X1 _41964_ (
    .A1(_21658_),
    .A2(_00007_[2]),
    .ZN(_07562_)
  );
  INV_X1 _41965_ (
    .A(_07562_),
    .ZN(_07563_)
  );
  AND2_X1 _41966_ (
    .A1(_07561_),
    .A2(_07563_),
    .ZN(_07564_)
  );
  AND2_X1 _41967_ (
    .A1(_21469_),
    .A2(_22077_),
    .ZN(_07565_)
  );
  INV_X1 _41968_ (
    .A(_07565_),
    .ZN(_07566_)
  );
  AND2_X1 _41969_ (
    .A1(_21768_),
    .A2(_00007_[2]),
    .ZN(_07567_)
  );
  INV_X1 _41970_ (
    .A(_07567_),
    .ZN(_07568_)
  );
  AND2_X1 _41971_ (
    .A1(\cpuregs[9] [15]),
    .A2(_22077_),
    .ZN(_07569_)
  );
  INV_X1 _41972_ (
    .A(_07569_),
    .ZN(_07570_)
  );
  AND2_X1 _41973_ (
    .A1(\cpuregs[13] [15]),
    .A2(_00007_[2]),
    .ZN(_07571_)
  );
  INV_X1 _41974_ (
    .A(_07571_),
    .ZN(_07572_)
  );
  AND2_X1 _41975_ (
    .A1(_07570_),
    .A2(_07572_),
    .ZN(_07573_)
  );
  INV_X1 _41976_ (
    .A(_07573_),
    .ZN(_07574_)
  );
  AND2_X1 _41977_ (
    .A1(_00007_[0]),
    .A2(_07574_),
    .ZN(_07575_)
  );
  INV_X1 _41978_ (
    .A(_07575_),
    .ZN(_07576_)
  );
  AND2_X1 _41979_ (
    .A1(\cpuregs[12] [15]),
    .A2(_00007_[2]),
    .ZN(_07577_)
  );
  INV_X1 _41980_ (
    .A(_07577_),
    .ZN(_07578_)
  );
  AND2_X1 _41981_ (
    .A1(\cpuregs[8] [15]),
    .A2(_22077_),
    .ZN(_07579_)
  );
  INV_X1 _41982_ (
    .A(_07579_),
    .ZN(_07580_)
  );
  AND2_X1 _41983_ (
    .A1(_07578_),
    .A2(_07580_),
    .ZN(_07581_)
  );
  INV_X1 _41984_ (
    .A(_07581_),
    .ZN(_07582_)
  );
  AND2_X1 _41985_ (
    .A1(_22152_),
    .A2(_07582_),
    .ZN(_07583_)
  );
  INV_X1 _41986_ (
    .A(_07583_),
    .ZN(_07584_)
  );
  AND2_X1 _41987_ (
    .A1(_07576_),
    .A2(_07584_),
    .ZN(_07585_)
  );
  AND2_X1 _41988_ (
    .A1(_21681_),
    .A2(_00007_[2]),
    .ZN(_07586_)
  );
  INV_X1 _41989_ (
    .A(_07586_),
    .ZN(_07587_)
  );
  AND2_X1 _41990_ (
    .A1(_21965_),
    .A2(_22077_),
    .ZN(_07588_)
  );
  INV_X1 _41991_ (
    .A(_07588_),
    .ZN(_07589_)
  );
  AND2_X1 _41992_ (
    .A1(_07587_),
    .A2(_07589_),
    .ZN(_07590_)
  );
  AND2_X1 _41993_ (
    .A1(_22152_),
    .A2(_07590_),
    .ZN(_07591_)
  );
  INV_X1 _41994_ (
    .A(_07591_),
    .ZN(_07592_)
  );
  AND2_X1 _41995_ (
    .A1(_21524_),
    .A2(_22077_),
    .ZN(_07593_)
  );
  INV_X1 _41996_ (
    .A(_07593_),
    .ZN(_07594_)
  );
  AND2_X1 _41997_ (
    .A1(_21744_),
    .A2(_00007_[2]),
    .ZN(_07595_)
  );
  INV_X1 _41998_ (
    .A(_07595_),
    .ZN(_07596_)
  );
  AND2_X1 _41999_ (
    .A1(_00007_[0]),
    .A2(_07596_),
    .ZN(_07597_)
  );
  AND2_X1 _42000_ (
    .A1(_07594_),
    .A2(_07597_),
    .ZN(_07598_)
  );
  INV_X1 _42001_ (
    .A(_07598_),
    .ZN(_07599_)
  );
  AND2_X1 _42002_ (
    .A1(_07592_),
    .A2(_07599_),
    .ZN(_07600_)
  );
  AND2_X1 _42003_ (
    .A1(_22152_),
    .A2(_07523_),
    .ZN(_07601_)
  );
  AND2_X1 _42004_ (
    .A1(_07521_),
    .A2(_07601_),
    .ZN(_07602_)
  );
  INV_X1 _42005_ (
    .A(_07602_),
    .ZN(_07603_)
  );
  AND2_X1 _42006_ (
    .A1(_00007_[0]),
    .A2(_07525_),
    .ZN(_07604_)
  );
  AND2_X1 _42007_ (
    .A1(_07527_),
    .A2(_07604_),
    .ZN(_07605_)
  );
  INV_X1 _42008_ (
    .A(_07605_),
    .ZN(_07606_)
  );
  AND2_X1 _42009_ (
    .A1(_07603_),
    .A2(_07606_),
    .ZN(_07607_)
  );
  AND2_X1 _42010_ (
    .A1(_00007_[1]),
    .A2(_07607_),
    .ZN(_07608_)
  );
  INV_X1 _42011_ (
    .A(_07608_),
    .ZN(_07609_)
  );
  AND2_X1 _42012_ (
    .A1(_00007_[0]),
    .A2(_07568_),
    .ZN(_07610_)
  );
  AND2_X1 _42013_ (
    .A1(_07566_),
    .A2(_07610_),
    .ZN(_07611_)
  );
  INV_X1 _42014_ (
    .A(_07611_),
    .ZN(_07612_)
  );
  AND2_X1 _42015_ (
    .A1(_22152_),
    .A2(_07564_),
    .ZN(_07613_)
  );
  INV_X1 _42016_ (
    .A(_07613_),
    .ZN(_07614_)
  );
  AND2_X1 _42017_ (
    .A1(_07612_),
    .A2(_07614_),
    .ZN(_07615_)
  );
  AND2_X1 _42018_ (
    .A1(_22078_),
    .A2(_07615_),
    .ZN(_07616_)
  );
  INV_X1 _42019_ (
    .A(_07616_),
    .ZN(_07617_)
  );
  AND2_X1 _42020_ (
    .A1(_22109_),
    .A2(_07617_),
    .ZN(_07618_)
  );
  AND2_X1 _42021_ (
    .A1(_07609_),
    .A2(_07618_),
    .ZN(_07619_)
  );
  INV_X1 _42022_ (
    .A(_07619_),
    .ZN(_07620_)
  );
  AND2_X1 _42023_ (
    .A1(_21929_),
    .A2(_22077_),
    .ZN(_07621_)
  );
  INV_X1 _42024_ (
    .A(_07621_),
    .ZN(_07622_)
  );
  AND2_X1 _42025_ (
    .A1(_21945_),
    .A2(_00007_[2]),
    .ZN(_07623_)
  );
  INV_X1 _42026_ (
    .A(_07623_),
    .ZN(_07624_)
  );
  AND2_X1 _42027_ (
    .A1(_00007_[0]),
    .A2(_07624_),
    .ZN(_07625_)
  );
  AND2_X1 _42028_ (
    .A1(_07622_),
    .A2(_07625_),
    .ZN(_07626_)
  );
  INV_X1 _42029_ (
    .A(_07626_),
    .ZN(_07627_)
  );
  AND2_X1 _42030_ (
    .A1(_21877_),
    .A2(_22077_),
    .ZN(_07628_)
  );
  INV_X1 _42031_ (
    .A(_07628_),
    .ZN(_07629_)
  );
  AND2_X1 _42032_ (
    .A1(_21857_),
    .A2(_00007_[2]),
    .ZN(_07630_)
  );
  INV_X1 _42033_ (
    .A(_07630_),
    .ZN(_07631_)
  );
  AND2_X1 _42034_ (
    .A1(_07629_),
    .A2(_07631_),
    .ZN(_07632_)
  );
  AND2_X1 _42035_ (
    .A1(_22152_),
    .A2(_07632_),
    .ZN(_07633_)
  );
  INV_X1 _42036_ (
    .A(_07633_),
    .ZN(_07634_)
  );
  AND2_X1 _42037_ (
    .A1(_07627_),
    .A2(_07634_),
    .ZN(_07635_)
  );
  AND2_X1 _42038_ (
    .A1(_00007_[1]),
    .A2(_07635_),
    .ZN(_07636_)
  );
  INV_X1 _42039_ (
    .A(_07636_),
    .ZN(_07637_)
  );
  AND2_X1 _42040_ (
    .A1(_21841_),
    .A2(_22077_),
    .ZN(_07638_)
  );
  INV_X1 _42041_ (
    .A(_07638_),
    .ZN(_07639_)
  );
  AND2_X1 _42042_ (
    .A1(_21897_),
    .A2(_00007_[2]),
    .ZN(_07640_)
  );
  INV_X1 _42043_ (
    .A(_07640_),
    .ZN(_07641_)
  );
  AND2_X1 _42044_ (
    .A1(_00007_[0]),
    .A2(_07641_),
    .ZN(_07642_)
  );
  AND2_X1 _42045_ (
    .A1(_07639_),
    .A2(_07642_),
    .ZN(_07643_)
  );
  INV_X1 _42046_ (
    .A(_07643_),
    .ZN(_07644_)
  );
  AND2_X1 _42047_ (
    .A1(_21575_),
    .A2(_22077_),
    .ZN(_07645_)
  );
  INV_X1 _42048_ (
    .A(_07645_),
    .ZN(_07646_)
  );
  AND2_X1 _42049_ (
    .A1(_21913_),
    .A2(_00007_[2]),
    .ZN(_07647_)
  );
  INV_X1 _42050_ (
    .A(_07647_),
    .ZN(_07648_)
  );
  AND2_X1 _42051_ (
    .A1(_07646_),
    .A2(_07648_),
    .ZN(_07649_)
  );
  AND2_X1 _42052_ (
    .A1(_22152_),
    .A2(_07649_),
    .ZN(_07650_)
  );
  INV_X1 _42053_ (
    .A(_07650_),
    .ZN(_07651_)
  );
  AND2_X1 _42054_ (
    .A1(_07644_),
    .A2(_07651_),
    .ZN(_07652_)
  );
  AND2_X1 _42055_ (
    .A1(_22078_),
    .A2(_07652_),
    .ZN(_07653_)
  );
  INV_X1 _42056_ (
    .A(_07653_),
    .ZN(_07654_)
  );
  AND2_X1 _42057_ (
    .A1(_00007_[3]),
    .A2(_07654_),
    .ZN(_07655_)
  );
  AND2_X1 _42058_ (
    .A1(_07637_),
    .A2(_07655_),
    .ZN(_07656_)
  );
  INV_X1 _42059_ (
    .A(_07656_),
    .ZN(_07657_)
  );
  AND2_X1 _42060_ (
    .A1(_00007_[4]),
    .A2(_07657_),
    .ZN(_07658_)
  );
  AND2_X1 _42061_ (
    .A1(_07620_),
    .A2(_07658_),
    .ZN(_07659_)
  );
  INV_X1 _42062_ (
    .A(_07659_),
    .ZN(_07660_)
  );
  AND2_X1 _42063_ (
    .A1(_00007_[1]),
    .A2(_07559_),
    .ZN(_07661_)
  );
  INV_X1 _42064_ (
    .A(_07661_),
    .ZN(_07662_)
  );
  AND2_X1 _42065_ (
    .A1(_22078_),
    .A2(_07600_),
    .ZN(_07663_)
  );
  INV_X1 _42066_ (
    .A(_07663_),
    .ZN(_07664_)
  );
  AND2_X1 _42067_ (
    .A1(_22109_),
    .A2(_07664_),
    .ZN(_07665_)
  );
  AND2_X1 _42068_ (
    .A1(_07662_),
    .A2(_07665_),
    .ZN(_07666_)
  );
  INV_X1 _42069_ (
    .A(_07666_),
    .ZN(_07667_)
  );
  AND2_X1 _42070_ (
    .A1(_00007_[1]),
    .A2(_07544_),
    .ZN(_07668_)
  );
  INV_X1 _42071_ (
    .A(_07668_),
    .ZN(_07669_)
  );
  AND2_X1 _42072_ (
    .A1(_22078_),
    .A2(_07585_),
    .ZN(_07670_)
  );
  INV_X1 _42073_ (
    .A(_07670_),
    .ZN(_07671_)
  );
  AND2_X1 _42074_ (
    .A1(_00007_[3]),
    .A2(_07671_),
    .ZN(_07672_)
  );
  AND2_X1 _42075_ (
    .A1(_07669_),
    .A2(_07672_),
    .ZN(_07673_)
  );
  INV_X1 _42076_ (
    .A(_07673_),
    .ZN(_07674_)
  );
  AND2_X1 _42077_ (
    .A1(_07667_),
    .A2(_07674_),
    .ZN(_07675_)
  );
  AND2_X1 _42078_ (
    .A1(_22144_),
    .A2(_07675_),
    .ZN(_07676_)
  );
  INV_X1 _42079_ (
    .A(_07676_),
    .ZN(_07677_)
  );
  AND2_X1 _42080_ (
    .A1(_07660_),
    .A2(_07677_),
    .ZN(_07678_)
  );
  AND2_X1 _42081_ (
    .A1(_05842_),
    .A2(_07678_),
    .ZN(_07679_)
  );
  INV_X1 _42082_ (
    .A(_07679_),
    .ZN(_07680_)
  );
  AND2_X1 _42083_ (
    .A1(_21215_),
    .A2(_04963_),
    .ZN(_07681_)
  );
  INV_X1 _42084_ (
    .A(_07681_),
    .ZN(_07682_)
  );
  AND2_X1 _42085_ (
    .A1(_04962_),
    .A2(_07680_),
    .ZN(_07683_)
  );
  AND2_X1 _42086_ (
    .A1(_07519_),
    .A2(_07683_),
    .ZN(_07684_)
  );
  INV_X1 _42087_ (
    .A(_07684_),
    .ZN(_07685_)
  );
  AND2_X1 _42088_ (
    .A1(_07682_),
    .A2(_07685_),
    .ZN(_00296_)
  );
  AND2_X1 _42089_ (
    .A1(decoded_imm[16]),
    .A2(_04966_),
    .ZN(_07686_)
  );
  INV_X1 _42090_ (
    .A(_07686_),
    .ZN(_07687_)
  );
  AND2_X1 _42091_ (
    .A1(_21603_),
    .A2(_22077_),
    .ZN(_07688_)
  );
  INV_X1 _42092_ (
    .A(_07688_),
    .ZN(_07689_)
  );
  AND2_X1 _42093_ (
    .A1(_21423_),
    .A2(_00007_[2]),
    .ZN(_07690_)
  );
  INV_X1 _42094_ (
    .A(_07690_),
    .ZN(_07691_)
  );
  AND2_X1 _42095_ (
    .A1(_21382_),
    .A2(_00007_[2]),
    .ZN(_07692_)
  );
  INV_X1 _42096_ (
    .A(_07692_),
    .ZN(_07693_)
  );
  AND2_X1 _42097_ (
    .A1(_21628_),
    .A2(_22077_),
    .ZN(_07694_)
  );
  INV_X1 _42098_ (
    .A(_07694_),
    .ZN(_07695_)
  );
  AND2_X1 _42099_ (
    .A1(\cpuregs[11] [16]),
    .A2(_22077_),
    .ZN(_07696_)
  );
  INV_X1 _42100_ (
    .A(_07696_),
    .ZN(_07697_)
  );
  AND2_X1 _42101_ (
    .A1(\cpuregs[15] [16]),
    .A2(_00007_[2]),
    .ZN(_07698_)
  );
  INV_X1 _42102_ (
    .A(_07698_),
    .ZN(_07699_)
  );
  AND2_X1 _42103_ (
    .A1(_07697_),
    .A2(_07699_),
    .ZN(_07700_)
  );
  INV_X1 _42104_ (
    .A(_07700_),
    .ZN(_07701_)
  );
  AND2_X1 _42105_ (
    .A1(_00007_[0]),
    .A2(_07701_),
    .ZN(_07702_)
  );
  INV_X1 _42106_ (
    .A(_07702_),
    .ZN(_07703_)
  );
  AND2_X1 _42107_ (
    .A1(\cpuregs[14] [16]),
    .A2(_00007_[2]),
    .ZN(_07704_)
  );
  INV_X1 _42108_ (
    .A(_07704_),
    .ZN(_07705_)
  );
  AND2_X1 _42109_ (
    .A1(\cpuregs[10] [16]),
    .A2(_22077_),
    .ZN(_07706_)
  );
  INV_X1 _42110_ (
    .A(_07706_),
    .ZN(_07707_)
  );
  AND2_X1 _42111_ (
    .A1(_07705_),
    .A2(_07707_),
    .ZN(_07708_)
  );
  INV_X1 _42112_ (
    .A(_07708_),
    .ZN(_07709_)
  );
  AND2_X1 _42113_ (
    .A1(_22152_),
    .A2(_07709_),
    .ZN(_07710_)
  );
  INV_X1 _42114_ (
    .A(_07710_),
    .ZN(_07711_)
  );
  AND2_X1 _42115_ (
    .A1(_07703_),
    .A2(_07711_),
    .ZN(_07712_)
  );
  AND2_X1 _42116_ (
    .A1(_21553_),
    .A2(_22077_),
    .ZN(_07713_)
  );
  INV_X1 _42117_ (
    .A(_07713_),
    .ZN(_07714_)
  );
  AND2_X1 _42118_ (
    .A1(_21819_),
    .A2(_00007_[2]),
    .ZN(_07715_)
  );
  INV_X1 _42119_ (
    .A(_07715_),
    .ZN(_07716_)
  );
  AND2_X1 _42120_ (
    .A1(_22152_),
    .A2(_07716_),
    .ZN(_07717_)
  );
  AND2_X1 _42121_ (
    .A1(_07714_),
    .A2(_07717_),
    .ZN(_07718_)
  );
  INV_X1 _42122_ (
    .A(_07718_),
    .ZN(_07719_)
  );
  AND2_X1 _42123_ (
    .A1(_21792_),
    .A2(_00007_[2]),
    .ZN(_07720_)
  );
  INV_X1 _42124_ (
    .A(_07720_),
    .ZN(_07721_)
  );
  AND2_X1 _42125_ (
    .A1(_21500_),
    .A2(_22077_),
    .ZN(_07722_)
  );
  INV_X1 _42126_ (
    .A(_07722_),
    .ZN(_07723_)
  );
  AND2_X1 _42127_ (
    .A1(_00007_[0]),
    .A2(_07723_),
    .ZN(_07724_)
  );
  AND2_X1 _42128_ (
    .A1(_07721_),
    .A2(_07724_),
    .ZN(_07725_)
  );
  INV_X1 _42129_ (
    .A(_07725_),
    .ZN(_07726_)
  );
  AND2_X1 _42130_ (
    .A1(_07719_),
    .A2(_07726_),
    .ZN(_07727_)
  );
  AND2_X1 _42131_ (
    .A1(_21448_),
    .A2(_22077_),
    .ZN(_07728_)
  );
  INV_X1 _42132_ (
    .A(_07728_),
    .ZN(_07729_)
  );
  AND2_X1 _42133_ (
    .A1(_21659_),
    .A2(_00007_[2]),
    .ZN(_07730_)
  );
  INV_X1 _42134_ (
    .A(_07730_),
    .ZN(_07731_)
  );
  AND2_X1 _42135_ (
    .A1(_07729_),
    .A2(_07731_),
    .ZN(_07732_)
  );
  AND2_X1 _42136_ (
    .A1(_21470_),
    .A2(_22077_),
    .ZN(_07733_)
  );
  INV_X1 _42137_ (
    .A(_07733_),
    .ZN(_07734_)
  );
  AND2_X1 _42138_ (
    .A1(_21769_),
    .A2(_00007_[2]),
    .ZN(_07735_)
  );
  INV_X1 _42139_ (
    .A(_07735_),
    .ZN(_07736_)
  );
  AND2_X1 _42140_ (
    .A1(\cpuregs[9] [16]),
    .A2(_22077_),
    .ZN(_07737_)
  );
  INV_X1 _42141_ (
    .A(_07737_),
    .ZN(_07738_)
  );
  AND2_X1 _42142_ (
    .A1(\cpuregs[13] [16]),
    .A2(_00007_[2]),
    .ZN(_07739_)
  );
  INV_X1 _42143_ (
    .A(_07739_),
    .ZN(_07740_)
  );
  AND2_X1 _42144_ (
    .A1(_07738_),
    .A2(_07740_),
    .ZN(_07741_)
  );
  INV_X1 _42145_ (
    .A(_07741_),
    .ZN(_07742_)
  );
  AND2_X1 _42146_ (
    .A1(_00007_[0]),
    .A2(_07742_),
    .ZN(_07743_)
  );
  INV_X1 _42147_ (
    .A(_07743_),
    .ZN(_07744_)
  );
  AND2_X1 _42148_ (
    .A1(\cpuregs[12] [16]),
    .A2(_00007_[2]),
    .ZN(_07745_)
  );
  INV_X1 _42149_ (
    .A(_07745_),
    .ZN(_07746_)
  );
  AND2_X1 _42150_ (
    .A1(\cpuregs[8] [16]),
    .A2(_22077_),
    .ZN(_07747_)
  );
  INV_X1 _42151_ (
    .A(_07747_),
    .ZN(_07748_)
  );
  AND2_X1 _42152_ (
    .A1(_07746_),
    .A2(_07748_),
    .ZN(_07749_)
  );
  INV_X1 _42153_ (
    .A(_07749_),
    .ZN(_07750_)
  );
  AND2_X1 _42154_ (
    .A1(_22152_),
    .A2(_07750_),
    .ZN(_07751_)
  );
  INV_X1 _42155_ (
    .A(_07751_),
    .ZN(_07752_)
  );
  AND2_X1 _42156_ (
    .A1(_07744_),
    .A2(_07752_),
    .ZN(_07753_)
  );
  AND2_X1 _42157_ (
    .A1(_21682_),
    .A2(_00007_[2]),
    .ZN(_07754_)
  );
  INV_X1 _42158_ (
    .A(_07754_),
    .ZN(_07755_)
  );
  AND2_X1 _42159_ (
    .A1(_21966_),
    .A2(_22077_),
    .ZN(_07756_)
  );
  INV_X1 _42160_ (
    .A(_07756_),
    .ZN(_07757_)
  );
  AND2_X1 _42161_ (
    .A1(_07755_),
    .A2(_07757_),
    .ZN(_07758_)
  );
  AND2_X1 _42162_ (
    .A1(_22152_),
    .A2(_07758_),
    .ZN(_07759_)
  );
  INV_X1 _42163_ (
    .A(_07759_),
    .ZN(_07760_)
  );
  AND2_X1 _42164_ (
    .A1(_21525_),
    .A2(_22077_),
    .ZN(_07761_)
  );
  INV_X1 _42165_ (
    .A(_07761_),
    .ZN(_07762_)
  );
  AND2_X1 _42166_ (
    .A1(_21745_),
    .A2(_00007_[2]),
    .ZN(_07763_)
  );
  INV_X1 _42167_ (
    .A(_07763_),
    .ZN(_07764_)
  );
  AND2_X1 _42168_ (
    .A1(_00007_[0]),
    .A2(_07764_),
    .ZN(_07765_)
  );
  AND2_X1 _42169_ (
    .A1(_07762_),
    .A2(_07765_),
    .ZN(_07766_)
  );
  INV_X1 _42170_ (
    .A(_07766_),
    .ZN(_07767_)
  );
  AND2_X1 _42171_ (
    .A1(_07760_),
    .A2(_07767_),
    .ZN(_07768_)
  );
  AND2_X1 _42172_ (
    .A1(_22152_),
    .A2(_07691_),
    .ZN(_07769_)
  );
  AND2_X1 _42173_ (
    .A1(_07689_),
    .A2(_07769_),
    .ZN(_07770_)
  );
  INV_X1 _42174_ (
    .A(_07770_),
    .ZN(_07771_)
  );
  AND2_X1 _42175_ (
    .A1(_00007_[0]),
    .A2(_07693_),
    .ZN(_07772_)
  );
  AND2_X1 _42176_ (
    .A1(_07695_),
    .A2(_07772_),
    .ZN(_07773_)
  );
  INV_X1 _42177_ (
    .A(_07773_),
    .ZN(_07774_)
  );
  AND2_X1 _42178_ (
    .A1(_07771_),
    .A2(_07774_),
    .ZN(_07775_)
  );
  AND2_X1 _42179_ (
    .A1(_00007_[1]),
    .A2(_07775_),
    .ZN(_07776_)
  );
  INV_X1 _42180_ (
    .A(_07776_),
    .ZN(_07777_)
  );
  AND2_X1 _42181_ (
    .A1(_00007_[0]),
    .A2(_07736_),
    .ZN(_07778_)
  );
  AND2_X1 _42182_ (
    .A1(_07734_),
    .A2(_07778_),
    .ZN(_07779_)
  );
  INV_X1 _42183_ (
    .A(_07779_),
    .ZN(_07780_)
  );
  AND2_X1 _42184_ (
    .A1(_22152_),
    .A2(_07732_),
    .ZN(_07781_)
  );
  INV_X1 _42185_ (
    .A(_07781_),
    .ZN(_07782_)
  );
  AND2_X1 _42186_ (
    .A1(_07780_),
    .A2(_07782_),
    .ZN(_07783_)
  );
  AND2_X1 _42187_ (
    .A1(_22078_),
    .A2(_07783_),
    .ZN(_07784_)
  );
  INV_X1 _42188_ (
    .A(_07784_),
    .ZN(_07785_)
  );
  AND2_X1 _42189_ (
    .A1(_07777_),
    .A2(_07785_),
    .ZN(_07786_)
  );
  AND2_X1 _42190_ (
    .A1(_22109_),
    .A2(_07786_),
    .ZN(_07787_)
  );
  INV_X1 _42191_ (
    .A(_07787_),
    .ZN(_07788_)
  );
  AND2_X1 _42192_ (
    .A1(_21930_),
    .A2(_22077_),
    .ZN(_07789_)
  );
  INV_X1 _42193_ (
    .A(_07789_),
    .ZN(_07790_)
  );
  AND2_X1 _42194_ (
    .A1(_21946_),
    .A2(_00007_[2]),
    .ZN(_07791_)
  );
  INV_X1 _42195_ (
    .A(_07791_),
    .ZN(_07792_)
  );
  AND2_X1 _42196_ (
    .A1(_00007_[0]),
    .A2(_07792_),
    .ZN(_07793_)
  );
  AND2_X1 _42197_ (
    .A1(_07790_),
    .A2(_07793_),
    .ZN(_07794_)
  );
  INV_X1 _42198_ (
    .A(_07794_),
    .ZN(_07795_)
  );
  AND2_X1 _42199_ (
    .A1(_21878_),
    .A2(_22077_),
    .ZN(_07796_)
  );
  INV_X1 _42200_ (
    .A(_07796_),
    .ZN(_07797_)
  );
  AND2_X1 _42201_ (
    .A1(_21858_),
    .A2(_00007_[2]),
    .ZN(_07798_)
  );
  INV_X1 _42202_ (
    .A(_07798_),
    .ZN(_07799_)
  );
  AND2_X1 _42203_ (
    .A1(_07797_),
    .A2(_07799_),
    .ZN(_07800_)
  );
  AND2_X1 _42204_ (
    .A1(_22152_),
    .A2(_07800_),
    .ZN(_07801_)
  );
  INV_X1 _42205_ (
    .A(_07801_),
    .ZN(_07802_)
  );
  AND2_X1 _42206_ (
    .A1(_07795_),
    .A2(_07802_),
    .ZN(_07803_)
  );
  AND2_X1 _42207_ (
    .A1(_00007_[1]),
    .A2(_07803_),
    .ZN(_07804_)
  );
  INV_X1 _42208_ (
    .A(_07804_),
    .ZN(_07805_)
  );
  AND2_X1 _42209_ (
    .A1(_21842_),
    .A2(_22077_),
    .ZN(_07806_)
  );
  INV_X1 _42210_ (
    .A(_07806_),
    .ZN(_07807_)
  );
  AND2_X1 _42211_ (
    .A1(_21898_),
    .A2(_00007_[2]),
    .ZN(_07808_)
  );
  INV_X1 _42212_ (
    .A(_07808_),
    .ZN(_07809_)
  );
  AND2_X1 _42213_ (
    .A1(_00007_[0]),
    .A2(_07809_),
    .ZN(_07810_)
  );
  AND2_X1 _42214_ (
    .A1(_07807_),
    .A2(_07810_),
    .ZN(_07811_)
  );
  INV_X1 _42215_ (
    .A(_07811_),
    .ZN(_07812_)
  );
  AND2_X1 _42216_ (
    .A1(_21576_),
    .A2(_22077_),
    .ZN(_07813_)
  );
  INV_X1 _42217_ (
    .A(_07813_),
    .ZN(_07814_)
  );
  AND2_X1 _42218_ (
    .A1(_21914_),
    .A2(_00007_[2]),
    .ZN(_07815_)
  );
  INV_X1 _42219_ (
    .A(_07815_),
    .ZN(_07816_)
  );
  AND2_X1 _42220_ (
    .A1(_07814_),
    .A2(_07816_),
    .ZN(_07817_)
  );
  AND2_X1 _42221_ (
    .A1(_22152_),
    .A2(_07817_),
    .ZN(_07818_)
  );
  INV_X1 _42222_ (
    .A(_07818_),
    .ZN(_07819_)
  );
  AND2_X1 _42223_ (
    .A1(_07812_),
    .A2(_07819_),
    .ZN(_07820_)
  );
  AND2_X1 _42224_ (
    .A1(_22078_),
    .A2(_07820_),
    .ZN(_07821_)
  );
  INV_X1 _42225_ (
    .A(_07821_),
    .ZN(_07822_)
  );
  AND2_X1 _42226_ (
    .A1(_00007_[3]),
    .A2(_07822_),
    .ZN(_07823_)
  );
  AND2_X1 _42227_ (
    .A1(_07805_),
    .A2(_07823_),
    .ZN(_07824_)
  );
  INV_X1 _42228_ (
    .A(_07824_),
    .ZN(_07825_)
  );
  AND2_X1 _42229_ (
    .A1(_00007_[4]),
    .A2(_07825_),
    .ZN(_07826_)
  );
  AND2_X1 _42230_ (
    .A1(_07788_),
    .A2(_07826_),
    .ZN(_07827_)
  );
  INV_X1 _42231_ (
    .A(_07827_),
    .ZN(_07828_)
  );
  AND2_X1 _42232_ (
    .A1(_00007_[1]),
    .A2(_07727_),
    .ZN(_07829_)
  );
  INV_X1 _42233_ (
    .A(_07829_),
    .ZN(_07830_)
  );
  AND2_X1 _42234_ (
    .A1(_22078_),
    .A2(_07768_),
    .ZN(_07831_)
  );
  INV_X1 _42235_ (
    .A(_07831_),
    .ZN(_07832_)
  );
  AND2_X1 _42236_ (
    .A1(_22109_),
    .A2(_07832_),
    .ZN(_07833_)
  );
  AND2_X1 _42237_ (
    .A1(_07830_),
    .A2(_07833_),
    .ZN(_07834_)
  );
  INV_X1 _42238_ (
    .A(_07834_),
    .ZN(_07835_)
  );
  AND2_X1 _42239_ (
    .A1(_00007_[1]),
    .A2(_07712_),
    .ZN(_07836_)
  );
  INV_X1 _42240_ (
    .A(_07836_),
    .ZN(_07837_)
  );
  AND2_X1 _42241_ (
    .A1(_22078_),
    .A2(_07753_),
    .ZN(_07838_)
  );
  INV_X1 _42242_ (
    .A(_07838_),
    .ZN(_07839_)
  );
  AND2_X1 _42243_ (
    .A1(_00007_[3]),
    .A2(_07839_),
    .ZN(_07840_)
  );
  AND2_X1 _42244_ (
    .A1(_07837_),
    .A2(_07840_),
    .ZN(_07841_)
  );
  INV_X1 _42245_ (
    .A(_07841_),
    .ZN(_07842_)
  );
  AND2_X1 _42246_ (
    .A1(_07835_),
    .A2(_07842_),
    .ZN(_07843_)
  );
  AND2_X1 _42247_ (
    .A1(_22144_),
    .A2(_07843_),
    .ZN(_07844_)
  );
  INV_X1 _42248_ (
    .A(_07844_),
    .ZN(_07845_)
  );
  AND2_X1 _42249_ (
    .A1(_07828_),
    .A2(_07845_),
    .ZN(_07846_)
  );
  AND2_X1 _42250_ (
    .A1(_05842_),
    .A2(_07846_),
    .ZN(_07847_)
  );
  INV_X1 _42251_ (
    .A(_07847_),
    .ZN(_07848_)
  );
  AND2_X1 _42252_ (
    .A1(_21216_),
    .A2(_04963_),
    .ZN(_07849_)
  );
  INV_X1 _42253_ (
    .A(_07849_),
    .ZN(_07850_)
  );
  AND2_X1 _42254_ (
    .A1(_04962_),
    .A2(_07848_),
    .ZN(_07851_)
  );
  AND2_X1 _42255_ (
    .A1(_07687_),
    .A2(_07851_),
    .ZN(_07852_)
  );
  INV_X1 _42256_ (
    .A(_07852_),
    .ZN(_07853_)
  );
  AND2_X1 _42257_ (
    .A1(_07850_),
    .A2(_07853_),
    .ZN(_00297_)
  );
  AND2_X1 _42258_ (
    .A1(\cpuregs[29] [17]),
    .A2(_00007_[2]),
    .ZN(_07854_)
  );
  INV_X1 _42259_ (
    .A(_07854_),
    .ZN(_07855_)
  );
  AND2_X1 _42260_ (
    .A1(\cpuregs[25] [17]),
    .A2(_22077_),
    .ZN(_07856_)
  );
  INV_X1 _42261_ (
    .A(_07856_),
    .ZN(_07857_)
  );
  AND2_X1 _42262_ (
    .A1(_00007_[0]),
    .A2(_07857_),
    .ZN(_07858_)
  );
  AND2_X1 _42263_ (
    .A1(_07855_),
    .A2(_07858_),
    .ZN(_07859_)
  );
  INV_X1 _42264_ (
    .A(_07859_),
    .ZN(_07860_)
  );
  AND2_X1 _42265_ (
    .A1(\cpuregs[24] [17]),
    .A2(_22077_),
    .ZN(_07861_)
  );
  INV_X1 _42266_ (
    .A(_07861_),
    .ZN(_07862_)
  );
  AND2_X1 _42267_ (
    .A1(\cpuregs[28] [17]),
    .A2(_00007_[2]),
    .ZN(_07863_)
  );
  INV_X1 _42268_ (
    .A(_07863_),
    .ZN(_07864_)
  );
  AND2_X1 _42269_ (
    .A1(_22152_),
    .A2(_07864_),
    .ZN(_07865_)
  );
  AND2_X1 _42270_ (
    .A1(_07862_),
    .A2(_07865_),
    .ZN(_07866_)
  );
  INV_X1 _42271_ (
    .A(_07866_),
    .ZN(_07867_)
  );
  AND2_X1 _42272_ (
    .A1(_22078_),
    .A2(_07867_),
    .ZN(_07868_)
  );
  AND2_X1 _42273_ (
    .A1(_07860_),
    .A2(_07868_),
    .ZN(_07869_)
  );
  INV_X1 _42274_ (
    .A(_07869_),
    .ZN(_07870_)
  );
  AND2_X1 _42275_ (
    .A1(\cpuregs[31] [17]),
    .A2(_00007_[2]),
    .ZN(_07871_)
  );
  INV_X1 _42276_ (
    .A(_07871_),
    .ZN(_07872_)
  );
  AND2_X1 _42277_ (
    .A1(\cpuregs[27] [17]),
    .A2(_22077_),
    .ZN(_07873_)
  );
  INV_X1 _42278_ (
    .A(_07873_),
    .ZN(_07874_)
  );
  AND2_X1 _42279_ (
    .A1(_00007_[0]),
    .A2(_07874_),
    .ZN(_07875_)
  );
  AND2_X1 _42280_ (
    .A1(_07872_),
    .A2(_07875_),
    .ZN(_07876_)
  );
  INV_X1 _42281_ (
    .A(_07876_),
    .ZN(_07877_)
  );
  AND2_X1 _42282_ (
    .A1(\cpuregs[26] [17]),
    .A2(_22077_),
    .ZN(_07878_)
  );
  INV_X1 _42283_ (
    .A(_07878_),
    .ZN(_07879_)
  );
  AND2_X1 _42284_ (
    .A1(\cpuregs[30] [17]),
    .A2(_00007_[2]),
    .ZN(_07880_)
  );
  INV_X1 _42285_ (
    .A(_07880_),
    .ZN(_07881_)
  );
  AND2_X1 _42286_ (
    .A1(_22152_),
    .A2(_07881_),
    .ZN(_07882_)
  );
  AND2_X1 _42287_ (
    .A1(_07879_),
    .A2(_07882_),
    .ZN(_07883_)
  );
  INV_X1 _42288_ (
    .A(_07883_),
    .ZN(_07884_)
  );
  AND2_X1 _42289_ (
    .A1(_00007_[1]),
    .A2(_07884_),
    .ZN(_07885_)
  );
  AND2_X1 _42290_ (
    .A1(_07877_),
    .A2(_07885_),
    .ZN(_07886_)
  );
  INV_X1 _42291_ (
    .A(_07886_),
    .ZN(_07887_)
  );
  AND2_X1 _42292_ (
    .A1(_07870_),
    .A2(_07887_),
    .ZN(_07888_)
  );
  INV_X1 _42293_ (
    .A(_07888_),
    .ZN(_07889_)
  );
  AND2_X1 _42294_ (
    .A1(_21586_),
    .A2(_22077_),
    .ZN(_07890_)
  );
  INV_X1 _42295_ (
    .A(_07890_),
    .ZN(_07891_)
  );
  AND2_X1 _42296_ (
    .A1(_21404_),
    .A2(_00007_[2]),
    .ZN(_07892_)
  );
  INV_X1 _42297_ (
    .A(_07892_),
    .ZN(_07893_)
  );
  AND2_X1 _42298_ (
    .A1(_00007_[0]),
    .A2(_07893_),
    .ZN(_07894_)
  );
  AND2_X1 _42299_ (
    .A1(_07891_),
    .A2(_07894_),
    .ZN(_07895_)
  );
  INV_X1 _42300_ (
    .A(_07895_),
    .ZN(_07896_)
  );
  AND2_X1 _42301_ (
    .A1(\cpuregs[14] [17]),
    .A2(_00007_[2]),
    .ZN(_07897_)
  );
  INV_X1 _42302_ (
    .A(_07897_),
    .ZN(_07898_)
  );
  AND2_X1 _42303_ (
    .A1(\cpuregs[10] [17]),
    .A2(_22077_),
    .ZN(_07899_)
  );
  INV_X1 _42304_ (
    .A(_07899_),
    .ZN(_07900_)
  );
  AND2_X1 _42305_ (
    .A1(_07898_),
    .A2(_07900_),
    .ZN(_07901_)
  );
  INV_X1 _42306_ (
    .A(_07901_),
    .ZN(_07902_)
  );
  AND2_X1 _42307_ (
    .A1(_22152_),
    .A2(_07902_),
    .ZN(_07903_)
  );
  INV_X1 _42308_ (
    .A(_07903_),
    .ZN(_07904_)
  );
  AND2_X1 _42309_ (
    .A1(_07896_),
    .A2(_07904_),
    .ZN(_07905_)
  );
  AND2_X1 _42310_ (
    .A1(_21721_),
    .A2(_22077_),
    .ZN(_07906_)
  );
  INV_X1 _42311_ (
    .A(_07906_),
    .ZN(_07907_)
  );
  AND2_X1 _42312_ (
    .A1(_21643_),
    .A2(_00007_[2]),
    .ZN(_07908_)
  );
  INV_X1 _42313_ (
    .A(_07908_),
    .ZN(_07909_)
  );
  AND2_X1 _42314_ (
    .A1(_00007_[0]),
    .A2(_07909_),
    .ZN(_07910_)
  );
  AND2_X1 _42315_ (
    .A1(_07907_),
    .A2(_07910_),
    .ZN(_07911_)
  );
  INV_X1 _42316_ (
    .A(_07911_),
    .ZN(_07912_)
  );
  AND2_X1 _42317_ (
    .A1(\cpuregs[12] [17]),
    .A2(_00007_[2]),
    .ZN(_07913_)
  );
  INV_X1 _42318_ (
    .A(_07913_),
    .ZN(_07914_)
  );
  AND2_X1 _42319_ (
    .A1(\cpuregs[8] [17]),
    .A2(_22077_),
    .ZN(_07915_)
  );
  INV_X1 _42320_ (
    .A(_07915_),
    .ZN(_07916_)
  );
  AND2_X1 _42321_ (
    .A1(_07914_),
    .A2(_07916_),
    .ZN(_07917_)
  );
  INV_X1 _42322_ (
    .A(_07917_),
    .ZN(_07918_)
  );
  AND2_X1 _42323_ (
    .A1(_22152_),
    .A2(_07918_),
    .ZN(_07919_)
  );
  INV_X1 _42324_ (
    .A(_07919_),
    .ZN(_07920_)
  );
  AND2_X1 _42325_ (
    .A1(_07912_),
    .A2(_07920_),
    .ZN(_07921_)
  );
  AND2_X1 _42326_ (
    .A1(_21449_),
    .A2(_22077_),
    .ZN(_07922_)
  );
  INV_X1 _42327_ (
    .A(_07922_),
    .ZN(_07923_)
  );
  AND2_X1 _42328_ (
    .A1(_21660_),
    .A2(_00007_[2]),
    .ZN(_07924_)
  );
  INV_X1 _42329_ (
    .A(_07924_),
    .ZN(_07925_)
  );
  AND2_X1 _42330_ (
    .A1(_07923_),
    .A2(_07925_),
    .ZN(_07926_)
  );
  AND2_X1 _42331_ (
    .A1(_21471_),
    .A2(_22077_),
    .ZN(_07927_)
  );
  INV_X1 _42332_ (
    .A(_07927_),
    .ZN(_07928_)
  );
  AND2_X1 _42333_ (
    .A1(_21770_),
    .A2(_00007_[2]),
    .ZN(_07929_)
  );
  INV_X1 _42334_ (
    .A(_07929_),
    .ZN(_07930_)
  );
  AND2_X1 _42335_ (
    .A1(_00007_[0]),
    .A2(_07930_),
    .ZN(_07931_)
  );
  AND2_X1 _42336_ (
    .A1(_07928_),
    .A2(_07931_),
    .ZN(_07932_)
  );
  INV_X1 _42337_ (
    .A(_07932_),
    .ZN(_07933_)
  );
  AND2_X1 _42338_ (
    .A1(_22152_),
    .A2(_07926_),
    .ZN(_07934_)
  );
  INV_X1 _42339_ (
    .A(_07934_),
    .ZN(_07935_)
  );
  AND2_X1 _42340_ (
    .A1(_07933_),
    .A2(_07935_),
    .ZN(_07936_)
  );
  AND2_X1 _42341_ (
    .A1(_21604_),
    .A2(_22077_),
    .ZN(_07937_)
  );
  INV_X1 _42342_ (
    .A(_07937_),
    .ZN(_07938_)
  );
  AND2_X1 _42343_ (
    .A1(_21424_),
    .A2(_00007_[2]),
    .ZN(_07939_)
  );
  INV_X1 _42344_ (
    .A(_07939_),
    .ZN(_07940_)
  );
  AND2_X1 _42345_ (
    .A1(_21383_),
    .A2(_00007_[2]),
    .ZN(_07941_)
  );
  INV_X1 _42346_ (
    .A(_07941_),
    .ZN(_07942_)
  );
  AND2_X1 _42347_ (
    .A1(_21629_),
    .A2(_22077_),
    .ZN(_07943_)
  );
  INV_X1 _42348_ (
    .A(_07943_),
    .ZN(_07944_)
  );
  AND2_X1 _42349_ (
    .A1(_22152_),
    .A2(_07940_),
    .ZN(_07945_)
  );
  AND2_X1 _42350_ (
    .A1(_07938_),
    .A2(_07945_),
    .ZN(_07946_)
  );
  INV_X1 _42351_ (
    .A(_07946_),
    .ZN(_07947_)
  );
  AND2_X1 _42352_ (
    .A1(_00007_[0]),
    .A2(_07942_),
    .ZN(_07948_)
  );
  AND2_X1 _42353_ (
    .A1(_07944_),
    .A2(_07948_),
    .ZN(_07949_)
  );
  INV_X1 _42354_ (
    .A(_07949_),
    .ZN(_07950_)
  );
  AND2_X1 _42355_ (
    .A1(_07947_),
    .A2(_07950_),
    .ZN(_07951_)
  );
  AND2_X1 _42356_ (
    .A1(_21554_),
    .A2(_22077_),
    .ZN(_07952_)
  );
  INV_X1 _42357_ (
    .A(_07952_),
    .ZN(_07953_)
  );
  AND2_X1 _42358_ (
    .A1(_21820_),
    .A2(_00007_[2]),
    .ZN(_07954_)
  );
  INV_X1 _42359_ (
    .A(_07954_),
    .ZN(_07955_)
  );
  AND2_X1 _42360_ (
    .A1(_22152_),
    .A2(_07955_),
    .ZN(_07956_)
  );
  AND2_X1 _42361_ (
    .A1(_07953_),
    .A2(_07956_),
    .ZN(_07957_)
  );
  INV_X1 _42362_ (
    .A(_07957_),
    .ZN(_07958_)
  );
  AND2_X1 _42363_ (
    .A1(_21501_),
    .A2(_22077_),
    .ZN(_07959_)
  );
  INV_X1 _42364_ (
    .A(_07959_),
    .ZN(_07960_)
  );
  AND2_X1 _42365_ (
    .A1(_21793_),
    .A2(_00007_[2]),
    .ZN(_07961_)
  );
  INV_X1 _42366_ (
    .A(_07961_),
    .ZN(_07962_)
  );
  AND2_X1 _42367_ (
    .A1(_00007_[0]),
    .A2(_07960_),
    .ZN(_07963_)
  );
  AND2_X1 _42368_ (
    .A1(_07962_),
    .A2(_07963_),
    .ZN(_07964_)
  );
  INV_X1 _42369_ (
    .A(_07964_),
    .ZN(_07965_)
  );
  AND2_X1 _42370_ (
    .A1(_07958_),
    .A2(_07965_),
    .ZN(_07966_)
  );
  AND2_X1 _42371_ (
    .A1(_21526_),
    .A2(_22077_),
    .ZN(_07967_)
  );
  INV_X1 _42372_ (
    .A(_07967_),
    .ZN(_07968_)
  );
  AND2_X1 _42373_ (
    .A1(_21746_),
    .A2(_00007_[2]),
    .ZN(_07969_)
  );
  INV_X1 _42374_ (
    .A(_07969_),
    .ZN(_07970_)
  );
  AND2_X1 _42375_ (
    .A1(_00007_[0]),
    .A2(_07970_),
    .ZN(_07971_)
  );
  AND2_X1 _42376_ (
    .A1(_07968_),
    .A2(_07971_),
    .ZN(_07972_)
  );
  INV_X1 _42377_ (
    .A(_07972_),
    .ZN(_07973_)
  );
  AND2_X1 _42378_ (
    .A1(\cpuregs[4] [17]),
    .A2(_00007_[2]),
    .ZN(_07974_)
  );
  INV_X1 _42379_ (
    .A(_07974_),
    .ZN(_07975_)
  );
  AND2_X1 _42380_ (
    .A1(\cpuregs[0] [17]),
    .A2(_22077_),
    .ZN(_07976_)
  );
  INV_X1 _42381_ (
    .A(_07976_),
    .ZN(_07977_)
  );
  AND2_X1 _42382_ (
    .A1(_07975_),
    .A2(_07977_),
    .ZN(_07978_)
  );
  INV_X1 _42383_ (
    .A(_07978_),
    .ZN(_07979_)
  );
  AND2_X1 _42384_ (
    .A1(_22152_),
    .A2(_07979_),
    .ZN(_07980_)
  );
  INV_X1 _42385_ (
    .A(_07980_),
    .ZN(_07981_)
  );
  AND2_X1 _42386_ (
    .A1(_07973_),
    .A2(_07981_),
    .ZN(_07982_)
  );
  AND2_X1 _42387_ (
    .A1(_00007_[1]),
    .A2(_07966_),
    .ZN(_07983_)
  );
  INV_X1 _42388_ (
    .A(_07983_),
    .ZN(_07984_)
  );
  AND2_X1 _42389_ (
    .A1(_22078_),
    .A2(_07982_),
    .ZN(_07985_)
  );
  INV_X1 _42390_ (
    .A(_07985_),
    .ZN(_07986_)
  );
  AND2_X1 _42391_ (
    .A1(_07984_),
    .A2(_07986_),
    .ZN(_07987_)
  );
  AND2_X1 _42392_ (
    .A1(_00007_[1]),
    .A2(_07951_),
    .ZN(_07988_)
  );
  INV_X1 _42393_ (
    .A(_07988_),
    .ZN(_07989_)
  );
  AND2_X1 _42394_ (
    .A1(_22078_),
    .A2(_07936_),
    .ZN(_07990_)
  );
  INV_X1 _42395_ (
    .A(_07990_),
    .ZN(_07991_)
  );
  AND2_X1 _42396_ (
    .A1(_22109_),
    .A2(_07991_),
    .ZN(_07992_)
  );
  AND2_X1 _42397_ (
    .A1(_07989_),
    .A2(_07992_),
    .ZN(_07993_)
  );
  INV_X1 _42398_ (
    .A(_07993_),
    .ZN(_07994_)
  );
  AND2_X1 _42399_ (
    .A1(_00007_[3]),
    .A2(_07889_),
    .ZN(_07995_)
  );
  INV_X1 _42400_ (
    .A(_07995_),
    .ZN(_07996_)
  );
  AND2_X1 _42401_ (
    .A1(_00007_[4]),
    .A2(_07996_),
    .ZN(_07997_)
  );
  AND2_X1 _42402_ (
    .A1(_07994_),
    .A2(_07997_),
    .ZN(_07998_)
  );
  INV_X1 _42403_ (
    .A(_07998_),
    .ZN(_07999_)
  );
  AND2_X1 _42404_ (
    .A1(_22109_),
    .A2(_07987_),
    .ZN(_08000_)
  );
  INV_X1 _42405_ (
    .A(_08000_),
    .ZN(_08001_)
  );
  AND2_X1 _42406_ (
    .A1(_00007_[1]),
    .A2(_07905_),
    .ZN(_08002_)
  );
  INV_X1 _42407_ (
    .A(_08002_),
    .ZN(_08003_)
  );
  AND2_X1 _42408_ (
    .A1(_22078_),
    .A2(_07921_),
    .ZN(_08004_)
  );
  INV_X1 _42409_ (
    .A(_08004_),
    .ZN(_08005_)
  );
  AND2_X1 _42410_ (
    .A1(_00007_[3]),
    .A2(_08005_),
    .ZN(_08006_)
  );
  AND2_X1 _42411_ (
    .A1(_08003_),
    .A2(_08006_),
    .ZN(_08007_)
  );
  INV_X1 _42412_ (
    .A(_08007_),
    .ZN(_08008_)
  );
  AND2_X1 _42413_ (
    .A1(_08001_),
    .A2(_08008_),
    .ZN(_08009_)
  );
  AND2_X1 _42414_ (
    .A1(_22144_),
    .A2(_08009_),
    .ZN(_08010_)
  );
  INV_X1 _42415_ (
    .A(_08010_),
    .ZN(_08011_)
  );
  AND2_X1 _42416_ (
    .A1(_07999_),
    .A2(_08011_),
    .ZN(_08012_)
  );
  AND2_X1 _42417_ (
    .A1(_05842_),
    .A2(_08012_),
    .ZN(_08013_)
  );
  INV_X1 _42418_ (
    .A(_08013_),
    .ZN(_08014_)
  );
  AND2_X1 _42419_ (
    .A1(decoded_imm[17]),
    .A2(_04966_),
    .ZN(_08015_)
  );
  INV_X1 _42420_ (
    .A(_08015_),
    .ZN(_08016_)
  );
  AND2_X1 _42421_ (
    .A1(_21217_),
    .A2(_04963_),
    .ZN(_08017_)
  );
  INV_X1 _42422_ (
    .A(_08017_),
    .ZN(_08018_)
  );
  AND2_X1 _42423_ (
    .A1(_04962_),
    .A2(_08016_),
    .ZN(_08019_)
  );
  AND2_X1 _42424_ (
    .A1(_08014_),
    .A2(_08019_),
    .ZN(_08020_)
  );
  INV_X1 _42425_ (
    .A(_08020_),
    .ZN(_08021_)
  );
  AND2_X1 _42426_ (
    .A1(_08018_),
    .A2(_08021_),
    .ZN(_00298_)
  );
  AND2_X1 _42427_ (
    .A1(decoded_imm[18]),
    .A2(_04966_),
    .ZN(_08022_)
  );
  INV_X1 _42428_ (
    .A(_08022_),
    .ZN(_08023_)
  );
  AND2_X1 _42429_ (
    .A1(\cpuregs[19] [18]),
    .A2(_22077_),
    .ZN(_08024_)
  );
  INV_X1 _42430_ (
    .A(_08024_),
    .ZN(_08025_)
  );
  AND2_X1 _42431_ (
    .A1(\cpuregs[23] [18]),
    .A2(_00007_[2]),
    .ZN(_08026_)
  );
  INV_X1 _42432_ (
    .A(_08026_),
    .ZN(_08027_)
  );
  AND2_X1 _42433_ (
    .A1(_08025_),
    .A2(_08027_),
    .ZN(_08028_)
  );
  INV_X1 _42434_ (
    .A(_08028_),
    .ZN(_08029_)
  );
  AND2_X1 _42435_ (
    .A1(_00007_[0]),
    .A2(_08029_),
    .ZN(_08030_)
  );
  INV_X1 _42436_ (
    .A(_08030_),
    .ZN(_08031_)
  );
  AND2_X1 _42437_ (
    .A1(\cpuregs[22] [18]),
    .A2(_00007_[2]),
    .ZN(_08032_)
  );
  INV_X1 _42438_ (
    .A(_08032_),
    .ZN(_08033_)
  );
  AND2_X1 _42439_ (
    .A1(\cpuregs[18] [18]),
    .A2(_22077_),
    .ZN(_08034_)
  );
  INV_X1 _42440_ (
    .A(_08034_),
    .ZN(_08035_)
  );
  AND2_X1 _42441_ (
    .A1(_08033_),
    .A2(_08035_),
    .ZN(_08036_)
  );
  INV_X1 _42442_ (
    .A(_08036_),
    .ZN(_08037_)
  );
  AND2_X1 _42443_ (
    .A1(_22152_),
    .A2(_08037_),
    .ZN(_08038_)
  );
  INV_X1 _42444_ (
    .A(_08038_),
    .ZN(_08039_)
  );
  AND2_X1 _42445_ (
    .A1(_21502_),
    .A2(_22077_),
    .ZN(_08040_)
  );
  INV_X1 _42446_ (
    .A(_08040_),
    .ZN(_08041_)
  );
  AND2_X1 _42447_ (
    .A1(_21794_),
    .A2(_00007_[2]),
    .ZN(_08042_)
  );
  INV_X1 _42448_ (
    .A(_08042_),
    .ZN(_08043_)
  );
  AND2_X1 _42449_ (
    .A1(_00007_[0]),
    .A2(_08043_),
    .ZN(_08044_)
  );
  AND2_X1 _42450_ (
    .A1(_08041_),
    .A2(_08044_),
    .ZN(_08045_)
  );
  INV_X1 _42451_ (
    .A(_08045_),
    .ZN(_08046_)
  );
  AND2_X1 _42452_ (
    .A1(_21821_),
    .A2(_00007_[2]),
    .ZN(_08047_)
  );
  INV_X1 _42453_ (
    .A(_08047_),
    .ZN(_08048_)
  );
  AND2_X1 _42454_ (
    .A1(_21555_),
    .A2(_22077_),
    .ZN(_08049_)
  );
  INV_X1 _42455_ (
    .A(_08049_),
    .ZN(_08050_)
  );
  AND2_X1 _42456_ (
    .A1(_22152_),
    .A2(_08050_),
    .ZN(_08051_)
  );
  AND2_X1 _42457_ (
    .A1(_08048_),
    .A2(_08051_),
    .ZN(_08052_)
  );
  INV_X1 _42458_ (
    .A(_08052_),
    .ZN(_08053_)
  );
  AND2_X1 _42459_ (
    .A1(\cpuregs[17] [18]),
    .A2(_22077_),
    .ZN(_08054_)
  );
  INV_X1 _42460_ (
    .A(_08054_),
    .ZN(_08055_)
  );
  AND2_X1 _42461_ (
    .A1(\cpuregs[21] [18]),
    .A2(_00007_[2]),
    .ZN(_08056_)
  );
  INV_X1 _42462_ (
    .A(_08056_),
    .ZN(_08057_)
  );
  AND2_X1 _42463_ (
    .A1(_08055_),
    .A2(_08057_),
    .ZN(_08058_)
  );
  INV_X1 _42464_ (
    .A(_08058_),
    .ZN(_08059_)
  );
  AND2_X1 _42465_ (
    .A1(_00007_[0]),
    .A2(_08059_),
    .ZN(_08060_)
  );
  INV_X1 _42466_ (
    .A(_08060_),
    .ZN(_08061_)
  );
  AND2_X1 _42467_ (
    .A1(\cpuregs[16] [18]),
    .A2(_22077_),
    .ZN(_08062_)
  );
  INV_X1 _42468_ (
    .A(_08062_),
    .ZN(_08063_)
  );
  AND2_X1 _42469_ (
    .A1(\cpuregs[20] [18]),
    .A2(_00007_[2]),
    .ZN(_08064_)
  );
  INV_X1 _42470_ (
    .A(_08064_),
    .ZN(_08065_)
  );
  AND2_X1 _42471_ (
    .A1(_08063_),
    .A2(_08065_),
    .ZN(_08066_)
  );
  INV_X1 _42472_ (
    .A(_08066_),
    .ZN(_08067_)
  );
  AND2_X1 _42473_ (
    .A1(_22152_),
    .A2(_08067_),
    .ZN(_08068_)
  );
  INV_X1 _42474_ (
    .A(_08068_),
    .ZN(_08069_)
  );
  AND2_X1 _42475_ (
    .A1(_08061_),
    .A2(_08069_),
    .ZN(_08070_)
  );
  AND2_X1 _42476_ (
    .A1(_21527_),
    .A2(_22077_),
    .ZN(_08071_)
  );
  INV_X1 _42477_ (
    .A(_08071_),
    .ZN(_08072_)
  );
  AND2_X1 _42478_ (
    .A1(_21747_),
    .A2(_00007_[2]),
    .ZN(_08073_)
  );
  INV_X1 _42479_ (
    .A(_08073_),
    .ZN(_08074_)
  );
  AND2_X1 _42480_ (
    .A1(_00007_[0]),
    .A2(_08074_),
    .ZN(_08075_)
  );
  AND2_X1 _42481_ (
    .A1(_08072_),
    .A2(_08075_),
    .ZN(_08076_)
  );
  INV_X1 _42482_ (
    .A(_08076_),
    .ZN(_08077_)
  );
  AND2_X1 _42483_ (
    .A1(_21968_),
    .A2(_22077_),
    .ZN(_08078_)
  );
  INV_X1 _42484_ (
    .A(_08078_),
    .ZN(_08079_)
  );
  AND2_X1 _42485_ (
    .A1(_21684_),
    .A2(_00007_[2]),
    .ZN(_08080_)
  );
  INV_X1 _42486_ (
    .A(_08080_),
    .ZN(_08081_)
  );
  AND2_X1 _42487_ (
    .A1(_08079_),
    .A2(_08081_),
    .ZN(_08082_)
  );
  AND2_X1 _42488_ (
    .A1(_22152_),
    .A2(_08082_),
    .ZN(_08083_)
  );
  INV_X1 _42489_ (
    .A(_08083_),
    .ZN(_08084_)
  );
  AND2_X1 _42490_ (
    .A1(_08077_),
    .A2(_08084_),
    .ZN(_08085_)
  );
  AND2_X1 _42491_ (
    .A1(_22078_),
    .A2(_08085_),
    .ZN(_08086_)
  );
  INV_X1 _42492_ (
    .A(_08086_),
    .ZN(_08087_)
  );
  AND2_X1 _42493_ (
    .A1(_00007_[1]),
    .A2(_08053_),
    .ZN(_08088_)
  );
  AND2_X1 _42494_ (
    .A1(_08046_),
    .A2(_08088_),
    .ZN(_08089_)
  );
  INV_X1 _42495_ (
    .A(_08089_),
    .ZN(_08090_)
  );
  AND2_X1 _42496_ (
    .A1(_08087_),
    .A2(_08090_),
    .ZN(_08091_)
  );
  AND2_X1 _42497_ (
    .A1(_22144_),
    .A2(_08091_),
    .ZN(_08092_)
  );
  INV_X1 _42498_ (
    .A(_08092_),
    .ZN(_08093_)
  );
  AND2_X1 _42499_ (
    .A1(_00007_[1]),
    .A2(_08039_),
    .ZN(_08094_)
  );
  AND2_X1 _42500_ (
    .A1(_08031_),
    .A2(_08094_),
    .ZN(_08095_)
  );
  INV_X1 _42501_ (
    .A(_08095_),
    .ZN(_08096_)
  );
  AND2_X1 _42502_ (
    .A1(_22078_),
    .A2(_08070_),
    .ZN(_08097_)
  );
  INV_X1 _42503_ (
    .A(_08097_),
    .ZN(_08098_)
  );
  AND2_X1 _42504_ (
    .A1(_08096_),
    .A2(_08098_),
    .ZN(_08099_)
  );
  AND2_X1 _42505_ (
    .A1(_00007_[4]),
    .A2(_08099_),
    .ZN(_08100_)
  );
  INV_X1 _42506_ (
    .A(_08100_),
    .ZN(_08101_)
  );
  AND2_X1 _42507_ (
    .A1(_08093_),
    .A2(_08101_),
    .ZN(_08102_)
  );
  AND2_X1 _42508_ (
    .A1(\cpuregs[26] [18]),
    .A2(_22077_),
    .ZN(_08103_)
  );
  INV_X1 _42509_ (
    .A(_08103_),
    .ZN(_08104_)
  );
  AND2_X1 _42510_ (
    .A1(\cpuregs[30] [18]),
    .A2(_00007_[2]),
    .ZN(_08105_)
  );
  INV_X1 _42511_ (
    .A(_08105_),
    .ZN(_08106_)
  );
  AND2_X1 _42512_ (
    .A1(_00007_[1]),
    .A2(_08106_),
    .ZN(_08107_)
  );
  AND2_X1 _42513_ (
    .A1(_08104_),
    .A2(_08107_),
    .ZN(_08108_)
  );
  INV_X1 _42514_ (
    .A(_08108_),
    .ZN(_08109_)
  );
  AND2_X1 _42515_ (
    .A1(\cpuregs[28] [18]),
    .A2(_00007_[2]),
    .ZN(_08110_)
  );
  INV_X1 _42516_ (
    .A(_08110_),
    .ZN(_08111_)
  );
  AND2_X1 _42517_ (
    .A1(\cpuregs[24] [18]),
    .A2(_22077_),
    .ZN(_08112_)
  );
  INV_X1 _42518_ (
    .A(_08112_),
    .ZN(_08113_)
  );
  AND2_X1 _42519_ (
    .A1(_22078_),
    .A2(_08113_),
    .ZN(_08114_)
  );
  AND2_X1 _42520_ (
    .A1(_08111_),
    .A2(_08114_),
    .ZN(_08115_)
  );
  INV_X1 _42521_ (
    .A(_08115_),
    .ZN(_08116_)
  );
  AND2_X1 _42522_ (
    .A1(_22152_),
    .A2(_08116_),
    .ZN(_08117_)
  );
  AND2_X1 _42523_ (
    .A1(_08109_),
    .A2(_08117_),
    .ZN(_08118_)
  );
  INV_X1 _42524_ (
    .A(_08118_),
    .ZN(_08119_)
  );
  AND2_X1 _42525_ (
    .A1(\cpuregs[27] [18]),
    .A2(_22077_),
    .ZN(_08120_)
  );
  INV_X1 _42526_ (
    .A(_08120_),
    .ZN(_08121_)
  );
  AND2_X1 _42527_ (
    .A1(\cpuregs[31] [18]),
    .A2(_00007_[2]),
    .ZN(_08122_)
  );
  INV_X1 _42528_ (
    .A(_08122_),
    .ZN(_08123_)
  );
  AND2_X1 _42529_ (
    .A1(_00007_[1]),
    .A2(_08123_),
    .ZN(_08124_)
  );
  AND2_X1 _42530_ (
    .A1(_08121_),
    .A2(_08124_),
    .ZN(_08125_)
  );
  INV_X1 _42531_ (
    .A(_08125_),
    .ZN(_08126_)
  );
  AND2_X1 _42532_ (
    .A1(\cpuregs[29] [18]),
    .A2(_00007_[2]),
    .ZN(_08127_)
  );
  INV_X1 _42533_ (
    .A(_08127_),
    .ZN(_08128_)
  );
  AND2_X1 _42534_ (
    .A1(\cpuregs[25] [18]),
    .A2(_22077_),
    .ZN(_08129_)
  );
  INV_X1 _42535_ (
    .A(_08129_),
    .ZN(_08130_)
  );
  AND2_X1 _42536_ (
    .A1(_22078_),
    .A2(_08130_),
    .ZN(_08131_)
  );
  AND2_X1 _42537_ (
    .A1(_08128_),
    .A2(_08131_),
    .ZN(_08132_)
  );
  INV_X1 _42538_ (
    .A(_08132_),
    .ZN(_08133_)
  );
  AND2_X1 _42539_ (
    .A1(_00007_[0]),
    .A2(_08133_),
    .ZN(_08134_)
  );
  AND2_X1 _42540_ (
    .A1(_08126_),
    .A2(_08134_),
    .ZN(_08135_)
  );
  INV_X1 _42541_ (
    .A(_08135_),
    .ZN(_08136_)
  );
  AND2_X1 _42542_ (
    .A1(_08119_),
    .A2(_08136_),
    .ZN(_08137_)
  );
  INV_X1 _42543_ (
    .A(_08137_),
    .ZN(_08138_)
  );
  AND2_X1 _42544_ (
    .A1(_00007_[4]),
    .A2(_08138_),
    .ZN(_08139_)
  );
  INV_X1 _42545_ (
    .A(_08139_),
    .ZN(_08140_)
  );
  AND2_X1 _42546_ (
    .A1(\cpuregs[12] [18]),
    .A2(_22078_),
    .ZN(_08141_)
  );
  INV_X1 _42547_ (
    .A(_08141_),
    .ZN(_08142_)
  );
  AND2_X1 _42548_ (
    .A1(\cpuregs[14] [18]),
    .A2(_00007_[1]),
    .ZN(_08143_)
  );
  INV_X1 _42549_ (
    .A(_08143_),
    .ZN(_08144_)
  );
  AND2_X1 _42550_ (
    .A1(_00007_[2]),
    .A2(_08144_),
    .ZN(_08145_)
  );
  AND2_X1 _42551_ (
    .A1(_08142_),
    .A2(_08145_),
    .ZN(_08146_)
  );
  INV_X1 _42552_ (
    .A(_08146_),
    .ZN(_08147_)
  );
  AND2_X1 _42553_ (
    .A1(\cpuregs[8] [18]),
    .A2(_22078_),
    .ZN(_08148_)
  );
  INV_X1 _42554_ (
    .A(_08148_),
    .ZN(_08149_)
  );
  AND2_X1 _42555_ (
    .A1(\cpuregs[10] [18]),
    .A2(_00007_[1]),
    .ZN(_08150_)
  );
  INV_X1 _42556_ (
    .A(_08150_),
    .ZN(_08151_)
  );
  AND2_X1 _42557_ (
    .A1(_22077_),
    .A2(_08151_),
    .ZN(_08152_)
  );
  AND2_X1 _42558_ (
    .A1(_08149_),
    .A2(_08152_),
    .ZN(_08153_)
  );
  INV_X1 _42559_ (
    .A(_08153_),
    .ZN(_08154_)
  );
  AND2_X1 _42560_ (
    .A1(_22152_),
    .A2(_08154_),
    .ZN(_08155_)
  );
  AND2_X1 _42561_ (
    .A1(_08147_),
    .A2(_08155_),
    .ZN(_08156_)
  );
  INV_X1 _42562_ (
    .A(_08156_),
    .ZN(_08157_)
  );
  AND2_X1 _42563_ (
    .A1(\cpuregs[13] [18]),
    .A2(_22078_),
    .ZN(_08158_)
  );
  INV_X1 _42564_ (
    .A(_08158_),
    .ZN(_08159_)
  );
  AND2_X1 _42565_ (
    .A1(\cpuregs[15] [18]),
    .A2(_00007_[1]),
    .ZN(_08160_)
  );
  INV_X1 _42566_ (
    .A(_08160_),
    .ZN(_08161_)
  );
  AND2_X1 _42567_ (
    .A1(_00007_[2]),
    .A2(_08161_),
    .ZN(_08162_)
  );
  AND2_X1 _42568_ (
    .A1(_08159_),
    .A2(_08162_),
    .ZN(_08163_)
  );
  INV_X1 _42569_ (
    .A(_08163_),
    .ZN(_08164_)
  );
  AND2_X1 _42570_ (
    .A1(\cpuregs[9] [18]),
    .A2(_22078_),
    .ZN(_08165_)
  );
  INV_X1 _42571_ (
    .A(_08165_),
    .ZN(_08166_)
  );
  AND2_X1 _42572_ (
    .A1(\cpuregs[11] [18]),
    .A2(_00007_[1]),
    .ZN(_08167_)
  );
  INV_X1 _42573_ (
    .A(_08167_),
    .ZN(_08168_)
  );
  AND2_X1 _42574_ (
    .A1(_22077_),
    .A2(_08168_),
    .ZN(_08169_)
  );
  AND2_X1 _42575_ (
    .A1(_08166_),
    .A2(_08169_),
    .ZN(_08170_)
  );
  INV_X1 _42576_ (
    .A(_08170_),
    .ZN(_08171_)
  );
  AND2_X1 _42577_ (
    .A1(_00007_[0]),
    .A2(_08171_),
    .ZN(_08172_)
  );
  AND2_X1 _42578_ (
    .A1(_08164_),
    .A2(_08172_),
    .ZN(_08173_)
  );
  INV_X1 _42579_ (
    .A(_08173_),
    .ZN(_08174_)
  );
  AND2_X1 _42580_ (
    .A1(_08157_),
    .A2(_08174_),
    .ZN(_08175_)
  );
  INV_X1 _42581_ (
    .A(_08175_),
    .ZN(_08176_)
  );
  AND2_X1 _42582_ (
    .A1(_22144_),
    .A2(_08176_),
    .ZN(_08177_)
  );
  INV_X1 _42583_ (
    .A(_08177_),
    .ZN(_08178_)
  );
  AND2_X1 _42584_ (
    .A1(_00007_[3]),
    .A2(_08178_),
    .ZN(_08179_)
  );
  AND2_X1 _42585_ (
    .A1(_08140_),
    .A2(_08179_),
    .ZN(_08180_)
  );
  INV_X1 _42586_ (
    .A(_08180_),
    .ZN(_08181_)
  );
  AND2_X1 _42587_ (
    .A1(_22109_),
    .A2(_08102_),
    .ZN(_08182_)
  );
  INV_X1 _42588_ (
    .A(_08182_),
    .ZN(_08183_)
  );
  AND2_X1 _42589_ (
    .A1(_08181_),
    .A2(_08183_),
    .ZN(_08184_)
  );
  AND2_X1 _42590_ (
    .A1(_05842_),
    .A2(_08184_),
    .ZN(_08185_)
  );
  INV_X1 _42591_ (
    .A(_08185_),
    .ZN(_08186_)
  );
  AND2_X1 _42592_ (
    .A1(_21218_),
    .A2(_04963_),
    .ZN(_08187_)
  );
  INV_X1 _42593_ (
    .A(_08187_),
    .ZN(_08188_)
  );
  AND2_X1 _42594_ (
    .A1(_04962_),
    .A2(_08186_),
    .ZN(_08189_)
  );
  AND2_X1 _42595_ (
    .A1(_08023_),
    .A2(_08189_),
    .ZN(_08190_)
  );
  INV_X1 _42596_ (
    .A(_08190_),
    .ZN(_08191_)
  );
  AND2_X1 _42597_ (
    .A1(_08188_),
    .A2(_08191_),
    .ZN(_00299_)
  );
  AND2_X1 _42598_ (
    .A1(_21605_),
    .A2(_22077_),
    .ZN(_08192_)
  );
  INV_X1 _42599_ (
    .A(_08192_),
    .ZN(_08193_)
  );
  AND2_X1 _42600_ (
    .A1(_21425_),
    .A2(_00007_[2]),
    .ZN(_08194_)
  );
  INV_X1 _42601_ (
    .A(_08194_),
    .ZN(_08195_)
  );
  AND2_X1 _42602_ (
    .A1(_21384_),
    .A2(_00007_[2]),
    .ZN(_08196_)
  );
  INV_X1 _42603_ (
    .A(_08196_),
    .ZN(_08197_)
  );
  AND2_X1 _42604_ (
    .A1(_21630_),
    .A2(_22077_),
    .ZN(_08198_)
  );
  INV_X1 _42605_ (
    .A(_08198_),
    .ZN(_08199_)
  );
  AND2_X1 _42606_ (
    .A1(\cpuregs[11] [19]),
    .A2(_22077_),
    .ZN(_08200_)
  );
  INV_X1 _42607_ (
    .A(_08200_),
    .ZN(_08201_)
  );
  AND2_X1 _42608_ (
    .A1(\cpuregs[15] [19]),
    .A2(_00007_[2]),
    .ZN(_08202_)
  );
  INV_X1 _42609_ (
    .A(_08202_),
    .ZN(_08203_)
  );
  AND2_X1 _42610_ (
    .A1(_08201_),
    .A2(_08203_),
    .ZN(_08204_)
  );
  INV_X1 _42611_ (
    .A(_08204_),
    .ZN(_08205_)
  );
  AND2_X1 _42612_ (
    .A1(_00007_[0]),
    .A2(_08205_),
    .ZN(_08206_)
  );
  INV_X1 _42613_ (
    .A(_08206_),
    .ZN(_08207_)
  );
  AND2_X1 _42614_ (
    .A1(\cpuregs[14] [19]),
    .A2(_00007_[2]),
    .ZN(_08208_)
  );
  INV_X1 _42615_ (
    .A(_08208_),
    .ZN(_08209_)
  );
  AND2_X1 _42616_ (
    .A1(\cpuregs[10] [19]),
    .A2(_22077_),
    .ZN(_08210_)
  );
  INV_X1 _42617_ (
    .A(_08210_),
    .ZN(_08211_)
  );
  AND2_X1 _42618_ (
    .A1(_08209_),
    .A2(_08211_),
    .ZN(_08212_)
  );
  INV_X1 _42619_ (
    .A(_08212_),
    .ZN(_08213_)
  );
  AND2_X1 _42620_ (
    .A1(_22152_),
    .A2(_08213_),
    .ZN(_08214_)
  );
  INV_X1 _42621_ (
    .A(_08214_),
    .ZN(_08215_)
  );
  AND2_X1 _42622_ (
    .A1(_08207_),
    .A2(_08215_),
    .ZN(_08216_)
  );
  AND2_X1 _42623_ (
    .A1(_21556_),
    .A2(_22077_),
    .ZN(_08217_)
  );
  INV_X1 _42624_ (
    .A(_08217_),
    .ZN(_08218_)
  );
  AND2_X1 _42625_ (
    .A1(_21822_),
    .A2(_00007_[2]),
    .ZN(_08219_)
  );
  INV_X1 _42626_ (
    .A(_08219_),
    .ZN(_08220_)
  );
  AND2_X1 _42627_ (
    .A1(_22152_),
    .A2(_08220_),
    .ZN(_08221_)
  );
  AND2_X1 _42628_ (
    .A1(_08218_),
    .A2(_08221_),
    .ZN(_08222_)
  );
  INV_X1 _42629_ (
    .A(_08222_),
    .ZN(_08223_)
  );
  AND2_X1 _42630_ (
    .A1(_21795_),
    .A2(_00007_[2]),
    .ZN(_08224_)
  );
  INV_X1 _42631_ (
    .A(_08224_),
    .ZN(_08225_)
  );
  AND2_X1 _42632_ (
    .A1(_21503_),
    .A2(_22077_),
    .ZN(_08226_)
  );
  INV_X1 _42633_ (
    .A(_08226_),
    .ZN(_08227_)
  );
  AND2_X1 _42634_ (
    .A1(_00007_[0]),
    .A2(_08227_),
    .ZN(_08228_)
  );
  AND2_X1 _42635_ (
    .A1(_08225_),
    .A2(_08228_),
    .ZN(_08229_)
  );
  INV_X1 _42636_ (
    .A(_08229_),
    .ZN(_08230_)
  );
  AND2_X1 _42637_ (
    .A1(_08223_),
    .A2(_08230_),
    .ZN(_08231_)
  );
  AND2_X1 _42638_ (
    .A1(_21450_),
    .A2(_22077_),
    .ZN(_08232_)
  );
  INV_X1 _42639_ (
    .A(_08232_),
    .ZN(_08233_)
  );
  AND2_X1 _42640_ (
    .A1(_21661_),
    .A2(_00007_[2]),
    .ZN(_08234_)
  );
  INV_X1 _42641_ (
    .A(_08234_),
    .ZN(_08235_)
  );
  AND2_X1 _42642_ (
    .A1(_08233_),
    .A2(_08235_),
    .ZN(_08236_)
  );
  AND2_X1 _42643_ (
    .A1(_21472_),
    .A2(_22077_),
    .ZN(_08237_)
  );
  INV_X1 _42644_ (
    .A(_08237_),
    .ZN(_08238_)
  );
  AND2_X1 _42645_ (
    .A1(_21771_),
    .A2(_00007_[2]),
    .ZN(_08239_)
  );
  INV_X1 _42646_ (
    .A(_08239_),
    .ZN(_08240_)
  );
  AND2_X1 _42647_ (
    .A1(\cpuregs[9] [19]),
    .A2(_22077_),
    .ZN(_08241_)
  );
  INV_X1 _42648_ (
    .A(_08241_),
    .ZN(_08242_)
  );
  AND2_X1 _42649_ (
    .A1(\cpuregs[13] [19]),
    .A2(_00007_[2]),
    .ZN(_08243_)
  );
  INV_X1 _42650_ (
    .A(_08243_),
    .ZN(_08244_)
  );
  AND2_X1 _42651_ (
    .A1(_08242_),
    .A2(_08244_),
    .ZN(_08245_)
  );
  INV_X1 _42652_ (
    .A(_08245_),
    .ZN(_08246_)
  );
  AND2_X1 _42653_ (
    .A1(_00007_[0]),
    .A2(_08246_),
    .ZN(_08247_)
  );
  INV_X1 _42654_ (
    .A(_08247_),
    .ZN(_08248_)
  );
  AND2_X1 _42655_ (
    .A1(\cpuregs[12] [19]),
    .A2(_00007_[2]),
    .ZN(_08249_)
  );
  INV_X1 _42656_ (
    .A(_08249_),
    .ZN(_08250_)
  );
  AND2_X1 _42657_ (
    .A1(\cpuregs[8] [19]),
    .A2(_22077_),
    .ZN(_08251_)
  );
  INV_X1 _42658_ (
    .A(_08251_),
    .ZN(_08252_)
  );
  AND2_X1 _42659_ (
    .A1(_08250_),
    .A2(_08252_),
    .ZN(_08253_)
  );
  INV_X1 _42660_ (
    .A(_08253_),
    .ZN(_08254_)
  );
  AND2_X1 _42661_ (
    .A1(_22152_),
    .A2(_08254_),
    .ZN(_08255_)
  );
  INV_X1 _42662_ (
    .A(_08255_),
    .ZN(_08256_)
  );
  AND2_X1 _42663_ (
    .A1(_08248_),
    .A2(_08256_),
    .ZN(_08257_)
  );
  AND2_X1 _42664_ (
    .A1(_21685_),
    .A2(_00007_[2]),
    .ZN(_08258_)
  );
  INV_X1 _42665_ (
    .A(_08258_),
    .ZN(_08259_)
  );
  AND2_X1 _42666_ (
    .A1(_21969_),
    .A2(_22077_),
    .ZN(_08260_)
  );
  INV_X1 _42667_ (
    .A(_08260_),
    .ZN(_08261_)
  );
  AND2_X1 _42668_ (
    .A1(_08259_),
    .A2(_08261_),
    .ZN(_08262_)
  );
  AND2_X1 _42669_ (
    .A1(_22152_),
    .A2(_08262_),
    .ZN(_08263_)
  );
  INV_X1 _42670_ (
    .A(_08263_),
    .ZN(_08264_)
  );
  AND2_X1 _42671_ (
    .A1(_21528_),
    .A2(_22077_),
    .ZN(_08265_)
  );
  INV_X1 _42672_ (
    .A(_08265_),
    .ZN(_08266_)
  );
  AND2_X1 _42673_ (
    .A1(_21748_),
    .A2(_00007_[2]),
    .ZN(_08267_)
  );
  INV_X1 _42674_ (
    .A(_08267_),
    .ZN(_08268_)
  );
  AND2_X1 _42675_ (
    .A1(_00007_[0]),
    .A2(_08268_),
    .ZN(_08269_)
  );
  AND2_X1 _42676_ (
    .A1(_08266_),
    .A2(_08269_),
    .ZN(_08270_)
  );
  INV_X1 _42677_ (
    .A(_08270_),
    .ZN(_08271_)
  );
  AND2_X1 _42678_ (
    .A1(_08264_),
    .A2(_08271_),
    .ZN(_08272_)
  );
  AND2_X1 _42679_ (
    .A1(_22152_),
    .A2(_08195_),
    .ZN(_08273_)
  );
  AND2_X1 _42680_ (
    .A1(_08193_),
    .A2(_08273_),
    .ZN(_08274_)
  );
  INV_X1 _42681_ (
    .A(_08274_),
    .ZN(_08275_)
  );
  AND2_X1 _42682_ (
    .A1(_00007_[0]),
    .A2(_08197_),
    .ZN(_08276_)
  );
  AND2_X1 _42683_ (
    .A1(_08199_),
    .A2(_08276_),
    .ZN(_08277_)
  );
  INV_X1 _42684_ (
    .A(_08277_),
    .ZN(_08278_)
  );
  AND2_X1 _42685_ (
    .A1(_08275_),
    .A2(_08278_),
    .ZN(_08279_)
  );
  AND2_X1 _42686_ (
    .A1(_00007_[1]),
    .A2(_08279_),
    .ZN(_08280_)
  );
  INV_X1 _42687_ (
    .A(_08280_),
    .ZN(_08281_)
  );
  AND2_X1 _42688_ (
    .A1(_00007_[0]),
    .A2(_08240_),
    .ZN(_08282_)
  );
  AND2_X1 _42689_ (
    .A1(_08238_),
    .A2(_08282_),
    .ZN(_08283_)
  );
  INV_X1 _42690_ (
    .A(_08283_),
    .ZN(_08284_)
  );
  AND2_X1 _42691_ (
    .A1(_22152_),
    .A2(_08236_),
    .ZN(_08285_)
  );
  INV_X1 _42692_ (
    .A(_08285_),
    .ZN(_08286_)
  );
  AND2_X1 _42693_ (
    .A1(_08284_),
    .A2(_08286_),
    .ZN(_08287_)
  );
  AND2_X1 _42694_ (
    .A1(_22078_),
    .A2(_08287_),
    .ZN(_08288_)
  );
  INV_X1 _42695_ (
    .A(_08288_),
    .ZN(_08289_)
  );
  AND2_X1 _42696_ (
    .A1(_22109_),
    .A2(_08289_),
    .ZN(_08290_)
  );
  AND2_X1 _42697_ (
    .A1(_08281_),
    .A2(_08290_),
    .ZN(_08291_)
  );
  INV_X1 _42698_ (
    .A(_08291_),
    .ZN(_08292_)
  );
  AND2_X1 _42699_ (
    .A1(_21931_),
    .A2(_22077_),
    .ZN(_08293_)
  );
  INV_X1 _42700_ (
    .A(_08293_),
    .ZN(_08294_)
  );
  AND2_X1 _42701_ (
    .A1(_21947_),
    .A2(_00007_[2]),
    .ZN(_08295_)
  );
  INV_X1 _42702_ (
    .A(_08295_),
    .ZN(_08296_)
  );
  AND2_X1 _42703_ (
    .A1(_00007_[0]),
    .A2(_08296_),
    .ZN(_08297_)
  );
  AND2_X1 _42704_ (
    .A1(_08294_),
    .A2(_08297_),
    .ZN(_08298_)
  );
  INV_X1 _42705_ (
    .A(_08298_),
    .ZN(_08299_)
  );
  AND2_X1 _42706_ (
    .A1(_21880_),
    .A2(_22077_),
    .ZN(_08300_)
  );
  INV_X1 _42707_ (
    .A(_08300_),
    .ZN(_08301_)
  );
  AND2_X1 _42708_ (
    .A1(_21859_),
    .A2(_00007_[2]),
    .ZN(_08302_)
  );
  INV_X1 _42709_ (
    .A(_08302_),
    .ZN(_08303_)
  );
  AND2_X1 _42710_ (
    .A1(_08301_),
    .A2(_08303_),
    .ZN(_08304_)
  );
  AND2_X1 _42711_ (
    .A1(_22152_),
    .A2(_08304_),
    .ZN(_08305_)
  );
  INV_X1 _42712_ (
    .A(_08305_),
    .ZN(_08306_)
  );
  AND2_X1 _42713_ (
    .A1(_08299_),
    .A2(_08306_),
    .ZN(_08307_)
  );
  AND2_X1 _42714_ (
    .A1(_00007_[1]),
    .A2(_08307_),
    .ZN(_08308_)
  );
  INV_X1 _42715_ (
    .A(_08308_),
    .ZN(_08309_)
  );
  AND2_X1 _42716_ (
    .A1(_21843_),
    .A2(_22077_),
    .ZN(_08310_)
  );
  INV_X1 _42717_ (
    .A(_08310_),
    .ZN(_08311_)
  );
  AND2_X1 _42718_ (
    .A1(_21899_),
    .A2(_00007_[2]),
    .ZN(_08312_)
  );
  INV_X1 _42719_ (
    .A(_08312_),
    .ZN(_08313_)
  );
  AND2_X1 _42720_ (
    .A1(_00007_[0]),
    .A2(_08313_),
    .ZN(_08314_)
  );
  AND2_X1 _42721_ (
    .A1(_08311_),
    .A2(_08314_),
    .ZN(_08315_)
  );
  INV_X1 _42722_ (
    .A(_08315_),
    .ZN(_08316_)
  );
  AND2_X1 _42723_ (
    .A1(_21577_),
    .A2(_22077_),
    .ZN(_08317_)
  );
  INV_X1 _42724_ (
    .A(_08317_),
    .ZN(_08318_)
  );
  AND2_X1 _42725_ (
    .A1(_21915_),
    .A2(_00007_[2]),
    .ZN(_08319_)
  );
  INV_X1 _42726_ (
    .A(_08319_),
    .ZN(_08320_)
  );
  AND2_X1 _42727_ (
    .A1(_08318_),
    .A2(_08320_),
    .ZN(_08321_)
  );
  AND2_X1 _42728_ (
    .A1(_22152_),
    .A2(_08321_),
    .ZN(_08322_)
  );
  INV_X1 _42729_ (
    .A(_08322_),
    .ZN(_08323_)
  );
  AND2_X1 _42730_ (
    .A1(_08316_),
    .A2(_08323_),
    .ZN(_08324_)
  );
  AND2_X1 _42731_ (
    .A1(_22078_),
    .A2(_08324_),
    .ZN(_08325_)
  );
  INV_X1 _42732_ (
    .A(_08325_),
    .ZN(_08326_)
  );
  AND2_X1 _42733_ (
    .A1(_00007_[3]),
    .A2(_08326_),
    .ZN(_08327_)
  );
  AND2_X1 _42734_ (
    .A1(_08309_),
    .A2(_08327_),
    .ZN(_08328_)
  );
  INV_X1 _42735_ (
    .A(_08328_),
    .ZN(_08329_)
  );
  AND2_X1 _42736_ (
    .A1(_00007_[4]),
    .A2(_08329_),
    .ZN(_08330_)
  );
  AND2_X1 _42737_ (
    .A1(_08292_),
    .A2(_08330_),
    .ZN(_08331_)
  );
  INV_X1 _42738_ (
    .A(_08331_),
    .ZN(_08332_)
  );
  AND2_X1 _42739_ (
    .A1(_00007_[1]),
    .A2(_08231_),
    .ZN(_08333_)
  );
  INV_X1 _42740_ (
    .A(_08333_),
    .ZN(_08334_)
  );
  AND2_X1 _42741_ (
    .A1(_22078_),
    .A2(_08272_),
    .ZN(_08335_)
  );
  INV_X1 _42742_ (
    .A(_08335_),
    .ZN(_08336_)
  );
  AND2_X1 _42743_ (
    .A1(_22109_),
    .A2(_08336_),
    .ZN(_08337_)
  );
  AND2_X1 _42744_ (
    .A1(_08334_),
    .A2(_08337_),
    .ZN(_08338_)
  );
  INV_X1 _42745_ (
    .A(_08338_),
    .ZN(_08339_)
  );
  AND2_X1 _42746_ (
    .A1(_00007_[1]),
    .A2(_08216_),
    .ZN(_08340_)
  );
  INV_X1 _42747_ (
    .A(_08340_),
    .ZN(_08341_)
  );
  AND2_X1 _42748_ (
    .A1(_22078_),
    .A2(_08257_),
    .ZN(_08342_)
  );
  INV_X1 _42749_ (
    .A(_08342_),
    .ZN(_08343_)
  );
  AND2_X1 _42750_ (
    .A1(_00007_[3]),
    .A2(_08343_),
    .ZN(_08344_)
  );
  AND2_X1 _42751_ (
    .A1(_08341_),
    .A2(_08344_),
    .ZN(_08345_)
  );
  INV_X1 _42752_ (
    .A(_08345_),
    .ZN(_08346_)
  );
  AND2_X1 _42753_ (
    .A1(_08339_),
    .A2(_08346_),
    .ZN(_08347_)
  );
  AND2_X1 _42754_ (
    .A1(_22144_),
    .A2(_08347_),
    .ZN(_08348_)
  );
  INV_X1 _42755_ (
    .A(_08348_),
    .ZN(_08349_)
  );
  AND2_X1 _42756_ (
    .A1(_08332_),
    .A2(_08349_),
    .ZN(_08350_)
  );
  AND2_X1 _42757_ (
    .A1(_05842_),
    .A2(_08350_),
    .ZN(_08351_)
  );
  INV_X1 _42758_ (
    .A(_08351_),
    .ZN(_08352_)
  );
  AND2_X1 _42759_ (
    .A1(decoded_imm[19]),
    .A2(_04966_),
    .ZN(_08353_)
  );
  INV_X1 _42760_ (
    .A(_08353_),
    .ZN(_08354_)
  );
  AND2_X1 _42761_ (
    .A1(_21219_),
    .A2(_04963_),
    .ZN(_08355_)
  );
  INV_X1 _42762_ (
    .A(_08355_),
    .ZN(_08356_)
  );
  AND2_X1 _42763_ (
    .A1(_04962_),
    .A2(_08354_),
    .ZN(_08357_)
  );
  AND2_X1 _42764_ (
    .A1(_08352_),
    .A2(_08357_),
    .ZN(_08358_)
  );
  INV_X1 _42765_ (
    .A(_08358_),
    .ZN(_08359_)
  );
  AND2_X1 _42766_ (
    .A1(_08356_),
    .A2(_08359_),
    .ZN(_00300_)
  );
  AND2_X1 _42767_ (
    .A1(decoded_imm[20]),
    .A2(_04966_),
    .ZN(_08360_)
  );
  INV_X1 _42768_ (
    .A(_08360_),
    .ZN(_08361_)
  );
  AND2_X1 _42769_ (
    .A1(\cpuregs[29] [20]),
    .A2(_00007_[2]),
    .ZN(_08362_)
  );
  INV_X1 _42770_ (
    .A(_08362_),
    .ZN(_08363_)
  );
  AND2_X1 _42771_ (
    .A1(\cpuregs[25] [20]),
    .A2(_22077_),
    .ZN(_08364_)
  );
  INV_X1 _42772_ (
    .A(_08364_),
    .ZN(_08365_)
  );
  AND2_X1 _42773_ (
    .A1(_00007_[0]),
    .A2(_08365_),
    .ZN(_08366_)
  );
  AND2_X1 _42774_ (
    .A1(_08363_),
    .A2(_08366_),
    .ZN(_08367_)
  );
  INV_X1 _42775_ (
    .A(_08367_),
    .ZN(_08368_)
  );
  AND2_X1 _42776_ (
    .A1(\cpuregs[24] [20]),
    .A2(_22077_),
    .ZN(_08369_)
  );
  INV_X1 _42777_ (
    .A(_08369_),
    .ZN(_08370_)
  );
  AND2_X1 _42778_ (
    .A1(\cpuregs[28] [20]),
    .A2(_00007_[2]),
    .ZN(_08371_)
  );
  INV_X1 _42779_ (
    .A(_08371_),
    .ZN(_08372_)
  );
  AND2_X1 _42780_ (
    .A1(_22152_),
    .A2(_08372_),
    .ZN(_08373_)
  );
  AND2_X1 _42781_ (
    .A1(_08370_),
    .A2(_08373_),
    .ZN(_08374_)
  );
  INV_X1 _42782_ (
    .A(_08374_),
    .ZN(_08375_)
  );
  AND2_X1 _42783_ (
    .A1(_22078_),
    .A2(_08375_),
    .ZN(_08376_)
  );
  AND2_X1 _42784_ (
    .A1(_08368_),
    .A2(_08376_),
    .ZN(_08377_)
  );
  INV_X1 _42785_ (
    .A(_08377_),
    .ZN(_08378_)
  );
  AND2_X1 _42786_ (
    .A1(\cpuregs[31] [20]),
    .A2(_00007_[2]),
    .ZN(_08379_)
  );
  INV_X1 _42787_ (
    .A(_08379_),
    .ZN(_08380_)
  );
  AND2_X1 _42788_ (
    .A1(\cpuregs[27] [20]),
    .A2(_22077_),
    .ZN(_08381_)
  );
  INV_X1 _42789_ (
    .A(_08381_),
    .ZN(_08382_)
  );
  AND2_X1 _42790_ (
    .A1(_00007_[0]),
    .A2(_08382_),
    .ZN(_08383_)
  );
  AND2_X1 _42791_ (
    .A1(_08380_),
    .A2(_08383_),
    .ZN(_08384_)
  );
  INV_X1 _42792_ (
    .A(_08384_),
    .ZN(_08385_)
  );
  AND2_X1 _42793_ (
    .A1(\cpuregs[26] [20]),
    .A2(_22077_),
    .ZN(_08386_)
  );
  INV_X1 _42794_ (
    .A(_08386_),
    .ZN(_08387_)
  );
  AND2_X1 _42795_ (
    .A1(\cpuregs[30] [20]),
    .A2(_00007_[2]),
    .ZN(_08388_)
  );
  INV_X1 _42796_ (
    .A(_08388_),
    .ZN(_08389_)
  );
  AND2_X1 _42797_ (
    .A1(_22152_),
    .A2(_08389_),
    .ZN(_08390_)
  );
  AND2_X1 _42798_ (
    .A1(_08387_),
    .A2(_08390_),
    .ZN(_08391_)
  );
  INV_X1 _42799_ (
    .A(_08391_),
    .ZN(_08392_)
  );
  AND2_X1 _42800_ (
    .A1(_00007_[1]),
    .A2(_08392_),
    .ZN(_08393_)
  );
  AND2_X1 _42801_ (
    .A1(_08385_),
    .A2(_08393_),
    .ZN(_08394_)
  );
  INV_X1 _42802_ (
    .A(_08394_),
    .ZN(_08395_)
  );
  AND2_X1 _42803_ (
    .A1(_08378_),
    .A2(_08395_),
    .ZN(_08396_)
  );
  INV_X1 _42804_ (
    .A(_08396_),
    .ZN(_08397_)
  );
  AND2_X1 _42805_ (
    .A1(\cpuregs[11] [20]),
    .A2(_22077_),
    .ZN(_08398_)
  );
  INV_X1 _42806_ (
    .A(_08398_),
    .ZN(_08399_)
  );
  AND2_X1 _42807_ (
    .A1(\cpuregs[15] [20]),
    .A2(_00007_[2]),
    .ZN(_08400_)
  );
  INV_X1 _42808_ (
    .A(_08400_),
    .ZN(_08401_)
  );
  AND2_X1 _42809_ (
    .A1(_08399_),
    .A2(_08401_),
    .ZN(_08402_)
  );
  INV_X1 _42810_ (
    .A(_08402_),
    .ZN(_08403_)
  );
  AND2_X1 _42811_ (
    .A1(_00007_[0]),
    .A2(_08403_),
    .ZN(_08404_)
  );
  INV_X1 _42812_ (
    .A(_08404_),
    .ZN(_08405_)
  );
  AND2_X1 _42813_ (
    .A1(\cpuregs[14] [20]),
    .A2(_00007_[2]),
    .ZN(_08406_)
  );
  INV_X1 _42814_ (
    .A(_08406_),
    .ZN(_08407_)
  );
  AND2_X1 _42815_ (
    .A1(\cpuregs[10] [20]),
    .A2(_22077_),
    .ZN(_08408_)
  );
  INV_X1 _42816_ (
    .A(_08408_),
    .ZN(_08409_)
  );
  AND2_X1 _42817_ (
    .A1(_08407_),
    .A2(_08409_),
    .ZN(_08410_)
  );
  INV_X1 _42818_ (
    .A(_08410_),
    .ZN(_08411_)
  );
  AND2_X1 _42819_ (
    .A1(_22152_),
    .A2(_08411_),
    .ZN(_08412_)
  );
  INV_X1 _42820_ (
    .A(_08412_),
    .ZN(_08413_)
  );
  AND2_X1 _42821_ (
    .A1(_08405_),
    .A2(_08413_),
    .ZN(_08414_)
  );
  AND2_X1 _42822_ (
    .A1(\cpuregs[9] [20]),
    .A2(_22077_),
    .ZN(_08415_)
  );
  INV_X1 _42823_ (
    .A(_08415_),
    .ZN(_08416_)
  );
  AND2_X1 _42824_ (
    .A1(\cpuregs[13] [20]),
    .A2(_00007_[2]),
    .ZN(_08417_)
  );
  INV_X1 _42825_ (
    .A(_08417_),
    .ZN(_08418_)
  );
  AND2_X1 _42826_ (
    .A1(_08416_),
    .A2(_08418_),
    .ZN(_08419_)
  );
  INV_X1 _42827_ (
    .A(_08419_),
    .ZN(_08420_)
  );
  AND2_X1 _42828_ (
    .A1(_00007_[0]),
    .A2(_08420_),
    .ZN(_08421_)
  );
  INV_X1 _42829_ (
    .A(_08421_),
    .ZN(_08422_)
  );
  AND2_X1 _42830_ (
    .A1(\cpuregs[12] [20]),
    .A2(_00007_[2]),
    .ZN(_08423_)
  );
  INV_X1 _42831_ (
    .A(_08423_),
    .ZN(_08424_)
  );
  AND2_X1 _42832_ (
    .A1(\cpuregs[8] [20]),
    .A2(_22077_),
    .ZN(_08425_)
  );
  INV_X1 _42833_ (
    .A(_08425_),
    .ZN(_08426_)
  );
  AND2_X1 _42834_ (
    .A1(_08424_),
    .A2(_08426_),
    .ZN(_08427_)
  );
  INV_X1 _42835_ (
    .A(_08427_),
    .ZN(_08428_)
  );
  AND2_X1 _42836_ (
    .A1(_22152_),
    .A2(_08428_),
    .ZN(_08429_)
  );
  INV_X1 _42837_ (
    .A(_08429_),
    .ZN(_08430_)
  );
  AND2_X1 _42838_ (
    .A1(_08422_),
    .A2(_08430_),
    .ZN(_08431_)
  );
  AND2_X1 _42839_ (
    .A1(_21451_),
    .A2(_22077_),
    .ZN(_08432_)
  );
  INV_X1 _42840_ (
    .A(_08432_),
    .ZN(_08433_)
  );
  AND2_X1 _42841_ (
    .A1(_21662_),
    .A2(_00007_[2]),
    .ZN(_08434_)
  );
  INV_X1 _42842_ (
    .A(_08434_),
    .ZN(_08435_)
  );
  AND2_X1 _42843_ (
    .A1(_08433_),
    .A2(_08435_),
    .ZN(_08436_)
  );
  AND2_X1 _42844_ (
    .A1(_21473_),
    .A2(_22077_),
    .ZN(_08437_)
  );
  INV_X1 _42845_ (
    .A(_08437_),
    .ZN(_08438_)
  );
  AND2_X1 _42846_ (
    .A1(_21772_),
    .A2(_00007_[2]),
    .ZN(_08439_)
  );
  INV_X1 _42847_ (
    .A(_08439_),
    .ZN(_08440_)
  );
  AND2_X1 _42848_ (
    .A1(_00007_[0]),
    .A2(_08440_),
    .ZN(_08441_)
  );
  AND2_X1 _42849_ (
    .A1(_08438_),
    .A2(_08441_),
    .ZN(_08442_)
  );
  INV_X1 _42850_ (
    .A(_08442_),
    .ZN(_08443_)
  );
  AND2_X1 _42851_ (
    .A1(_22152_),
    .A2(_08436_),
    .ZN(_08444_)
  );
  INV_X1 _42852_ (
    .A(_08444_),
    .ZN(_08445_)
  );
  AND2_X1 _42853_ (
    .A1(_08443_),
    .A2(_08445_),
    .ZN(_08446_)
  );
  AND2_X1 _42854_ (
    .A1(_21606_),
    .A2(_22077_),
    .ZN(_08447_)
  );
  INV_X1 _42855_ (
    .A(_08447_),
    .ZN(_08448_)
  );
  AND2_X1 _42856_ (
    .A1(_21426_),
    .A2(_00007_[2]),
    .ZN(_08449_)
  );
  INV_X1 _42857_ (
    .A(_08449_),
    .ZN(_08450_)
  );
  AND2_X1 _42858_ (
    .A1(_21385_),
    .A2(_00007_[2]),
    .ZN(_08451_)
  );
  INV_X1 _42859_ (
    .A(_08451_),
    .ZN(_08452_)
  );
  AND2_X1 _42860_ (
    .A1(_21631_),
    .A2(_22077_),
    .ZN(_08453_)
  );
  INV_X1 _42861_ (
    .A(_08453_),
    .ZN(_08454_)
  );
  AND2_X1 _42862_ (
    .A1(_22152_),
    .A2(_08450_),
    .ZN(_08455_)
  );
  AND2_X1 _42863_ (
    .A1(_08448_),
    .A2(_08455_),
    .ZN(_08456_)
  );
  INV_X1 _42864_ (
    .A(_08456_),
    .ZN(_08457_)
  );
  AND2_X1 _42865_ (
    .A1(_00007_[0]),
    .A2(_08452_),
    .ZN(_08458_)
  );
  AND2_X1 _42866_ (
    .A1(_08454_),
    .A2(_08458_),
    .ZN(_08459_)
  );
  INV_X1 _42867_ (
    .A(_08459_),
    .ZN(_08460_)
  );
  AND2_X1 _42868_ (
    .A1(_08457_),
    .A2(_08460_),
    .ZN(_08461_)
  );
  AND2_X1 _42869_ (
    .A1(_00007_[1]),
    .A2(_08461_),
    .ZN(_08462_)
  );
  INV_X1 _42870_ (
    .A(_08462_),
    .ZN(_08463_)
  );
  AND2_X1 _42871_ (
    .A1(_22078_),
    .A2(_08446_),
    .ZN(_08464_)
  );
  INV_X1 _42872_ (
    .A(_08464_),
    .ZN(_08465_)
  );
  AND2_X1 _42873_ (
    .A1(_08463_),
    .A2(_08465_),
    .ZN(_08466_)
  );
  AND2_X1 _42874_ (
    .A1(\cpuregs[2] [20]),
    .A2(_22077_),
    .ZN(_08467_)
  );
  INV_X1 _42875_ (
    .A(_08467_),
    .ZN(_08468_)
  );
  AND2_X1 _42876_ (
    .A1(\cpuregs[6] [20]),
    .A2(_00007_[2]),
    .ZN(_08469_)
  );
  INV_X1 _42877_ (
    .A(_08469_),
    .ZN(_08470_)
  );
  AND2_X1 _42878_ (
    .A1(_08468_),
    .A2(_08470_),
    .ZN(_08471_)
  );
  INV_X1 _42879_ (
    .A(_08471_),
    .ZN(_08472_)
  );
  AND2_X1 _42880_ (
    .A1(_22152_),
    .A2(_08472_),
    .ZN(_08473_)
  );
  INV_X1 _42881_ (
    .A(_08473_),
    .ZN(_08474_)
  );
  AND2_X1 _42882_ (
    .A1(\cpuregs[7] [20]),
    .A2(_00007_[2]),
    .ZN(_08475_)
  );
  INV_X1 _42883_ (
    .A(_08475_),
    .ZN(_08476_)
  );
  AND2_X1 _42884_ (
    .A1(\cpuregs[3] [20]),
    .A2(_22077_),
    .ZN(_08477_)
  );
  INV_X1 _42885_ (
    .A(_08477_),
    .ZN(_08478_)
  );
  AND2_X1 _42886_ (
    .A1(_08476_),
    .A2(_08478_),
    .ZN(_08479_)
  );
  INV_X1 _42887_ (
    .A(_08479_),
    .ZN(_08480_)
  );
  AND2_X1 _42888_ (
    .A1(_00007_[0]),
    .A2(_08480_),
    .ZN(_08481_)
  );
  INV_X1 _42889_ (
    .A(_08481_),
    .ZN(_08482_)
  );
  AND2_X1 _42890_ (
    .A1(_08474_),
    .A2(_08482_),
    .ZN(_08483_)
  );
  AND2_X1 _42891_ (
    .A1(\cpuregs[1] [20]),
    .A2(_22077_),
    .ZN(_08484_)
  );
  INV_X1 _42892_ (
    .A(_08484_),
    .ZN(_08485_)
  );
  AND2_X1 _42893_ (
    .A1(\cpuregs[5] [20]),
    .A2(_00007_[2]),
    .ZN(_08486_)
  );
  INV_X1 _42894_ (
    .A(_08486_),
    .ZN(_08487_)
  );
  AND2_X1 _42895_ (
    .A1(_08485_),
    .A2(_08487_),
    .ZN(_08488_)
  );
  INV_X1 _42896_ (
    .A(_08488_),
    .ZN(_08489_)
  );
  AND2_X1 _42897_ (
    .A1(_00007_[0]),
    .A2(_08489_),
    .ZN(_08490_)
  );
  INV_X1 _42898_ (
    .A(_08490_),
    .ZN(_08491_)
  );
  AND2_X1 _42899_ (
    .A1(\cpuregs[4] [20]),
    .A2(_00007_[2]),
    .ZN(_08492_)
  );
  INV_X1 _42900_ (
    .A(_08492_),
    .ZN(_08493_)
  );
  AND2_X1 _42901_ (
    .A1(\cpuregs[0] [20]),
    .A2(_22077_),
    .ZN(_08494_)
  );
  INV_X1 _42902_ (
    .A(_08494_),
    .ZN(_08495_)
  );
  AND2_X1 _42903_ (
    .A1(_08493_),
    .A2(_08495_),
    .ZN(_08496_)
  );
  INV_X1 _42904_ (
    .A(_08496_),
    .ZN(_08497_)
  );
  AND2_X1 _42905_ (
    .A1(_22152_),
    .A2(_08497_),
    .ZN(_08498_)
  );
  INV_X1 _42906_ (
    .A(_08498_),
    .ZN(_08499_)
  );
  AND2_X1 _42907_ (
    .A1(_08491_),
    .A2(_08499_),
    .ZN(_08500_)
  );
  AND2_X1 _42908_ (
    .A1(_00007_[1]),
    .A2(_08483_),
    .ZN(_08501_)
  );
  INV_X1 _42909_ (
    .A(_08501_),
    .ZN(_08502_)
  );
  AND2_X1 _42910_ (
    .A1(_22078_),
    .A2(_08500_),
    .ZN(_08503_)
  );
  INV_X1 _42911_ (
    .A(_08503_),
    .ZN(_08504_)
  );
  AND2_X1 _42912_ (
    .A1(_08502_),
    .A2(_08504_),
    .ZN(_08505_)
  );
  AND2_X1 _42913_ (
    .A1(_22109_),
    .A2(_08466_),
    .ZN(_08506_)
  );
  INV_X1 _42914_ (
    .A(_08506_),
    .ZN(_08507_)
  );
  AND2_X1 _42915_ (
    .A1(_00007_[3]),
    .A2(_08397_),
    .ZN(_08508_)
  );
  INV_X1 _42916_ (
    .A(_08508_),
    .ZN(_08509_)
  );
  AND2_X1 _42917_ (
    .A1(_00007_[4]),
    .A2(_08509_),
    .ZN(_08510_)
  );
  AND2_X1 _42918_ (
    .A1(_08507_),
    .A2(_08510_),
    .ZN(_08511_)
  );
  INV_X1 _42919_ (
    .A(_08511_),
    .ZN(_08512_)
  );
  AND2_X1 _42920_ (
    .A1(_00007_[1]),
    .A2(_08414_),
    .ZN(_08513_)
  );
  INV_X1 _42921_ (
    .A(_08513_),
    .ZN(_08514_)
  );
  AND2_X1 _42922_ (
    .A1(_22078_),
    .A2(_08431_),
    .ZN(_08515_)
  );
  INV_X1 _42923_ (
    .A(_08515_),
    .ZN(_08516_)
  );
  AND2_X1 _42924_ (
    .A1(_00007_[3]),
    .A2(_08516_),
    .ZN(_08517_)
  );
  AND2_X1 _42925_ (
    .A1(_08514_),
    .A2(_08517_),
    .ZN(_08518_)
  );
  INV_X1 _42926_ (
    .A(_08518_),
    .ZN(_08519_)
  );
  AND2_X1 _42927_ (
    .A1(_22109_),
    .A2(_08505_),
    .ZN(_08520_)
  );
  INV_X1 _42928_ (
    .A(_08520_),
    .ZN(_08521_)
  );
  AND2_X1 _42929_ (
    .A1(_08519_),
    .A2(_08521_),
    .ZN(_08522_)
  );
  AND2_X1 _42930_ (
    .A1(_22144_),
    .A2(_08522_),
    .ZN(_08523_)
  );
  INV_X1 _42931_ (
    .A(_08523_),
    .ZN(_08524_)
  );
  AND2_X1 _42932_ (
    .A1(_08512_),
    .A2(_08524_),
    .ZN(_08525_)
  );
  AND2_X1 _42933_ (
    .A1(_05842_),
    .A2(_08525_),
    .ZN(_08526_)
  );
  INV_X1 _42934_ (
    .A(_08526_),
    .ZN(_08527_)
  );
  AND2_X1 _42935_ (
    .A1(_21220_),
    .A2(_04963_),
    .ZN(_08528_)
  );
  INV_X1 _42936_ (
    .A(_08528_),
    .ZN(_08529_)
  );
  AND2_X1 _42937_ (
    .A1(_04962_),
    .A2(_08527_),
    .ZN(_08530_)
  );
  AND2_X1 _42938_ (
    .A1(_08361_),
    .A2(_08530_),
    .ZN(_08531_)
  );
  INV_X1 _42939_ (
    .A(_08531_),
    .ZN(_08532_)
  );
  AND2_X1 _42940_ (
    .A1(_08529_),
    .A2(_08532_),
    .ZN(_00301_)
  );
  AND2_X1 _42941_ (
    .A1(decoded_imm[21]),
    .A2(_04966_),
    .ZN(_08533_)
  );
  INV_X1 _42942_ (
    .A(_08533_),
    .ZN(_08534_)
  );
  AND2_X1 _42943_ (
    .A1(\cpuregs[19] [21]),
    .A2(_22077_),
    .ZN(_08535_)
  );
  INV_X1 _42944_ (
    .A(_08535_),
    .ZN(_08536_)
  );
  AND2_X1 _42945_ (
    .A1(\cpuregs[23] [21]),
    .A2(_00007_[2]),
    .ZN(_08537_)
  );
  INV_X1 _42946_ (
    .A(_08537_),
    .ZN(_08538_)
  );
  AND2_X1 _42947_ (
    .A1(_08536_),
    .A2(_08538_),
    .ZN(_08539_)
  );
  INV_X1 _42948_ (
    .A(_08539_),
    .ZN(_08540_)
  );
  AND2_X1 _42949_ (
    .A1(_00007_[0]),
    .A2(_08540_),
    .ZN(_08541_)
  );
  INV_X1 _42950_ (
    .A(_08541_),
    .ZN(_08542_)
  );
  AND2_X1 _42951_ (
    .A1(\cpuregs[22] [21]),
    .A2(_00007_[2]),
    .ZN(_08543_)
  );
  INV_X1 _42952_ (
    .A(_08543_),
    .ZN(_08544_)
  );
  AND2_X1 _42953_ (
    .A1(\cpuregs[18] [21]),
    .A2(_22077_),
    .ZN(_08545_)
  );
  INV_X1 _42954_ (
    .A(_08545_),
    .ZN(_08546_)
  );
  AND2_X1 _42955_ (
    .A1(_08544_),
    .A2(_08546_),
    .ZN(_08547_)
  );
  INV_X1 _42956_ (
    .A(_08547_),
    .ZN(_08548_)
  );
  AND2_X1 _42957_ (
    .A1(_22152_),
    .A2(_08548_),
    .ZN(_08549_)
  );
  INV_X1 _42958_ (
    .A(_08549_),
    .ZN(_08550_)
  );
  AND2_X1 _42959_ (
    .A1(_21504_),
    .A2(_22077_),
    .ZN(_08551_)
  );
  INV_X1 _42960_ (
    .A(_08551_),
    .ZN(_08552_)
  );
  AND2_X1 _42961_ (
    .A1(_21796_),
    .A2(_00007_[2]),
    .ZN(_08553_)
  );
  INV_X1 _42962_ (
    .A(_08553_),
    .ZN(_08554_)
  );
  AND2_X1 _42963_ (
    .A1(_00007_[0]),
    .A2(_08554_),
    .ZN(_08555_)
  );
  AND2_X1 _42964_ (
    .A1(_08552_),
    .A2(_08555_),
    .ZN(_08556_)
  );
  INV_X1 _42965_ (
    .A(_08556_),
    .ZN(_08557_)
  );
  AND2_X1 _42966_ (
    .A1(_21823_),
    .A2(_00007_[2]),
    .ZN(_08558_)
  );
  INV_X1 _42967_ (
    .A(_08558_),
    .ZN(_08559_)
  );
  AND2_X1 _42968_ (
    .A1(_21557_),
    .A2(_22077_),
    .ZN(_08560_)
  );
  INV_X1 _42969_ (
    .A(_08560_),
    .ZN(_08561_)
  );
  AND2_X1 _42970_ (
    .A1(_22152_),
    .A2(_08561_),
    .ZN(_08562_)
  );
  AND2_X1 _42971_ (
    .A1(_08559_),
    .A2(_08562_),
    .ZN(_08563_)
  );
  INV_X1 _42972_ (
    .A(_08563_),
    .ZN(_08564_)
  );
  AND2_X1 _42973_ (
    .A1(\cpuregs[17] [21]),
    .A2(_22077_),
    .ZN(_08565_)
  );
  INV_X1 _42974_ (
    .A(_08565_),
    .ZN(_08566_)
  );
  AND2_X1 _42975_ (
    .A1(\cpuregs[21] [21]),
    .A2(_00007_[2]),
    .ZN(_08567_)
  );
  INV_X1 _42976_ (
    .A(_08567_),
    .ZN(_08568_)
  );
  AND2_X1 _42977_ (
    .A1(_08566_),
    .A2(_08568_),
    .ZN(_08569_)
  );
  INV_X1 _42978_ (
    .A(_08569_),
    .ZN(_08570_)
  );
  AND2_X1 _42979_ (
    .A1(_00007_[0]),
    .A2(_08570_),
    .ZN(_08571_)
  );
  INV_X1 _42980_ (
    .A(_08571_),
    .ZN(_08572_)
  );
  AND2_X1 _42981_ (
    .A1(\cpuregs[16] [21]),
    .A2(_22077_),
    .ZN(_08573_)
  );
  INV_X1 _42982_ (
    .A(_08573_),
    .ZN(_08574_)
  );
  AND2_X1 _42983_ (
    .A1(\cpuregs[20] [21]),
    .A2(_00007_[2]),
    .ZN(_08575_)
  );
  INV_X1 _42984_ (
    .A(_08575_),
    .ZN(_08576_)
  );
  AND2_X1 _42985_ (
    .A1(_08574_),
    .A2(_08576_),
    .ZN(_08577_)
  );
  INV_X1 _42986_ (
    .A(_08577_),
    .ZN(_08578_)
  );
  AND2_X1 _42987_ (
    .A1(_22152_),
    .A2(_08578_),
    .ZN(_08579_)
  );
  INV_X1 _42988_ (
    .A(_08579_),
    .ZN(_08580_)
  );
  AND2_X1 _42989_ (
    .A1(_08572_),
    .A2(_08580_),
    .ZN(_08581_)
  );
  AND2_X1 _42990_ (
    .A1(_21529_),
    .A2(_22077_),
    .ZN(_08582_)
  );
  INV_X1 _42991_ (
    .A(_08582_),
    .ZN(_08583_)
  );
  AND2_X1 _42992_ (
    .A1(_21749_),
    .A2(_00007_[2]),
    .ZN(_08584_)
  );
  INV_X1 _42993_ (
    .A(_08584_),
    .ZN(_08585_)
  );
  AND2_X1 _42994_ (
    .A1(_00007_[0]),
    .A2(_08585_),
    .ZN(_08586_)
  );
  AND2_X1 _42995_ (
    .A1(_08583_),
    .A2(_08586_),
    .ZN(_08587_)
  );
  INV_X1 _42996_ (
    .A(_08587_),
    .ZN(_08588_)
  );
  AND2_X1 _42997_ (
    .A1(_21970_),
    .A2(_22077_),
    .ZN(_08589_)
  );
  INV_X1 _42998_ (
    .A(_08589_),
    .ZN(_08590_)
  );
  AND2_X1 _42999_ (
    .A1(_21686_),
    .A2(_00007_[2]),
    .ZN(_08591_)
  );
  INV_X1 _43000_ (
    .A(_08591_),
    .ZN(_08592_)
  );
  AND2_X1 _43001_ (
    .A1(_08590_),
    .A2(_08592_),
    .ZN(_08593_)
  );
  AND2_X1 _43002_ (
    .A1(_22152_),
    .A2(_08593_),
    .ZN(_08594_)
  );
  INV_X1 _43003_ (
    .A(_08594_),
    .ZN(_08595_)
  );
  AND2_X1 _43004_ (
    .A1(_08588_),
    .A2(_08595_),
    .ZN(_08596_)
  );
  AND2_X1 _43005_ (
    .A1(_22078_),
    .A2(_08596_),
    .ZN(_08597_)
  );
  INV_X1 _43006_ (
    .A(_08597_),
    .ZN(_08598_)
  );
  AND2_X1 _43007_ (
    .A1(_00007_[1]),
    .A2(_08564_),
    .ZN(_08599_)
  );
  AND2_X1 _43008_ (
    .A1(_08557_),
    .A2(_08599_),
    .ZN(_08600_)
  );
  INV_X1 _43009_ (
    .A(_08600_),
    .ZN(_08601_)
  );
  AND2_X1 _43010_ (
    .A1(_08598_),
    .A2(_08601_),
    .ZN(_08602_)
  );
  AND2_X1 _43011_ (
    .A1(_22144_),
    .A2(_08602_),
    .ZN(_08603_)
  );
  INV_X1 _43012_ (
    .A(_08603_),
    .ZN(_08604_)
  );
  AND2_X1 _43013_ (
    .A1(_00007_[1]),
    .A2(_08550_),
    .ZN(_08605_)
  );
  AND2_X1 _43014_ (
    .A1(_08542_),
    .A2(_08605_),
    .ZN(_08606_)
  );
  INV_X1 _43015_ (
    .A(_08606_),
    .ZN(_08607_)
  );
  AND2_X1 _43016_ (
    .A1(_22078_),
    .A2(_08581_),
    .ZN(_08608_)
  );
  INV_X1 _43017_ (
    .A(_08608_),
    .ZN(_08609_)
  );
  AND2_X1 _43018_ (
    .A1(_08607_),
    .A2(_08609_),
    .ZN(_08610_)
  );
  AND2_X1 _43019_ (
    .A1(_00007_[4]),
    .A2(_08610_),
    .ZN(_08611_)
  );
  INV_X1 _43020_ (
    .A(_08611_),
    .ZN(_08612_)
  );
  AND2_X1 _43021_ (
    .A1(_08604_),
    .A2(_08612_),
    .ZN(_08613_)
  );
  AND2_X1 _43022_ (
    .A1(\cpuregs[26] [21]),
    .A2(_22077_),
    .ZN(_08614_)
  );
  INV_X1 _43023_ (
    .A(_08614_),
    .ZN(_08615_)
  );
  AND2_X1 _43024_ (
    .A1(\cpuregs[30] [21]),
    .A2(_00007_[2]),
    .ZN(_08616_)
  );
  INV_X1 _43025_ (
    .A(_08616_),
    .ZN(_08617_)
  );
  AND2_X1 _43026_ (
    .A1(_00007_[1]),
    .A2(_08617_),
    .ZN(_08618_)
  );
  AND2_X1 _43027_ (
    .A1(_08615_),
    .A2(_08618_),
    .ZN(_08619_)
  );
  INV_X1 _43028_ (
    .A(_08619_),
    .ZN(_08620_)
  );
  AND2_X1 _43029_ (
    .A1(\cpuregs[28] [21]),
    .A2(_00007_[2]),
    .ZN(_08621_)
  );
  INV_X1 _43030_ (
    .A(_08621_),
    .ZN(_08622_)
  );
  AND2_X1 _43031_ (
    .A1(\cpuregs[24] [21]),
    .A2(_22077_),
    .ZN(_08623_)
  );
  INV_X1 _43032_ (
    .A(_08623_),
    .ZN(_08624_)
  );
  AND2_X1 _43033_ (
    .A1(_22078_),
    .A2(_08624_),
    .ZN(_08625_)
  );
  AND2_X1 _43034_ (
    .A1(_08622_),
    .A2(_08625_),
    .ZN(_08626_)
  );
  INV_X1 _43035_ (
    .A(_08626_),
    .ZN(_08627_)
  );
  AND2_X1 _43036_ (
    .A1(_22152_),
    .A2(_08627_),
    .ZN(_08628_)
  );
  AND2_X1 _43037_ (
    .A1(_08620_),
    .A2(_08628_),
    .ZN(_08629_)
  );
  INV_X1 _43038_ (
    .A(_08629_),
    .ZN(_08630_)
  );
  AND2_X1 _43039_ (
    .A1(\cpuregs[27] [21]),
    .A2(_22077_),
    .ZN(_08631_)
  );
  INV_X1 _43040_ (
    .A(_08631_),
    .ZN(_08632_)
  );
  AND2_X1 _43041_ (
    .A1(\cpuregs[31] [21]),
    .A2(_00007_[2]),
    .ZN(_08633_)
  );
  INV_X1 _43042_ (
    .A(_08633_),
    .ZN(_08634_)
  );
  AND2_X1 _43043_ (
    .A1(_00007_[1]),
    .A2(_08634_),
    .ZN(_08635_)
  );
  AND2_X1 _43044_ (
    .A1(_08632_),
    .A2(_08635_),
    .ZN(_08636_)
  );
  INV_X1 _43045_ (
    .A(_08636_),
    .ZN(_08637_)
  );
  AND2_X1 _43046_ (
    .A1(\cpuregs[29] [21]),
    .A2(_00007_[2]),
    .ZN(_08638_)
  );
  INV_X1 _43047_ (
    .A(_08638_),
    .ZN(_08639_)
  );
  AND2_X1 _43048_ (
    .A1(\cpuregs[25] [21]),
    .A2(_22077_),
    .ZN(_08640_)
  );
  INV_X1 _43049_ (
    .A(_08640_),
    .ZN(_08641_)
  );
  AND2_X1 _43050_ (
    .A1(_22078_),
    .A2(_08641_),
    .ZN(_08642_)
  );
  AND2_X1 _43051_ (
    .A1(_08639_),
    .A2(_08642_),
    .ZN(_08643_)
  );
  INV_X1 _43052_ (
    .A(_08643_),
    .ZN(_08644_)
  );
  AND2_X1 _43053_ (
    .A1(_00007_[0]),
    .A2(_08644_),
    .ZN(_08645_)
  );
  AND2_X1 _43054_ (
    .A1(_08637_),
    .A2(_08645_),
    .ZN(_08646_)
  );
  INV_X1 _43055_ (
    .A(_08646_),
    .ZN(_08647_)
  );
  AND2_X1 _43056_ (
    .A1(_08630_),
    .A2(_08647_),
    .ZN(_08648_)
  );
  INV_X1 _43057_ (
    .A(_08648_),
    .ZN(_08649_)
  );
  AND2_X1 _43058_ (
    .A1(_00007_[4]),
    .A2(_08649_),
    .ZN(_08650_)
  );
  INV_X1 _43059_ (
    .A(_08650_),
    .ZN(_08651_)
  );
  AND2_X1 _43060_ (
    .A1(\cpuregs[12] [21]),
    .A2(_22078_),
    .ZN(_08652_)
  );
  INV_X1 _43061_ (
    .A(_08652_),
    .ZN(_08653_)
  );
  AND2_X1 _43062_ (
    .A1(\cpuregs[14] [21]),
    .A2(_00007_[1]),
    .ZN(_08654_)
  );
  INV_X1 _43063_ (
    .A(_08654_),
    .ZN(_08655_)
  );
  AND2_X1 _43064_ (
    .A1(_00007_[2]),
    .A2(_08655_),
    .ZN(_08656_)
  );
  AND2_X1 _43065_ (
    .A1(_08653_),
    .A2(_08656_),
    .ZN(_08657_)
  );
  INV_X1 _43066_ (
    .A(_08657_),
    .ZN(_08658_)
  );
  AND2_X1 _43067_ (
    .A1(\cpuregs[8] [21]),
    .A2(_22078_),
    .ZN(_08659_)
  );
  INV_X1 _43068_ (
    .A(_08659_),
    .ZN(_08660_)
  );
  AND2_X1 _43069_ (
    .A1(\cpuregs[10] [21]),
    .A2(_00007_[1]),
    .ZN(_08661_)
  );
  INV_X1 _43070_ (
    .A(_08661_),
    .ZN(_08662_)
  );
  AND2_X1 _43071_ (
    .A1(_22077_),
    .A2(_08662_),
    .ZN(_08663_)
  );
  AND2_X1 _43072_ (
    .A1(_08660_),
    .A2(_08663_),
    .ZN(_08664_)
  );
  INV_X1 _43073_ (
    .A(_08664_),
    .ZN(_08665_)
  );
  AND2_X1 _43074_ (
    .A1(_22152_),
    .A2(_08665_),
    .ZN(_08666_)
  );
  AND2_X1 _43075_ (
    .A1(_08658_),
    .A2(_08666_),
    .ZN(_08667_)
  );
  INV_X1 _43076_ (
    .A(_08667_),
    .ZN(_08668_)
  );
  AND2_X1 _43077_ (
    .A1(\cpuregs[13] [21]),
    .A2(_22078_),
    .ZN(_08669_)
  );
  INV_X1 _43078_ (
    .A(_08669_),
    .ZN(_08670_)
  );
  AND2_X1 _43079_ (
    .A1(\cpuregs[15] [21]),
    .A2(_00007_[1]),
    .ZN(_08671_)
  );
  INV_X1 _43080_ (
    .A(_08671_),
    .ZN(_08672_)
  );
  AND2_X1 _43081_ (
    .A1(_00007_[2]),
    .A2(_08672_),
    .ZN(_08673_)
  );
  AND2_X1 _43082_ (
    .A1(_08670_),
    .A2(_08673_),
    .ZN(_08674_)
  );
  INV_X1 _43083_ (
    .A(_08674_),
    .ZN(_08675_)
  );
  AND2_X1 _43084_ (
    .A1(\cpuregs[9] [21]),
    .A2(_22078_),
    .ZN(_08676_)
  );
  INV_X1 _43085_ (
    .A(_08676_),
    .ZN(_08677_)
  );
  AND2_X1 _43086_ (
    .A1(\cpuregs[11] [21]),
    .A2(_00007_[1]),
    .ZN(_08678_)
  );
  INV_X1 _43087_ (
    .A(_08678_),
    .ZN(_08679_)
  );
  AND2_X1 _43088_ (
    .A1(_22077_),
    .A2(_08679_),
    .ZN(_08680_)
  );
  AND2_X1 _43089_ (
    .A1(_08677_),
    .A2(_08680_),
    .ZN(_08681_)
  );
  INV_X1 _43090_ (
    .A(_08681_),
    .ZN(_08682_)
  );
  AND2_X1 _43091_ (
    .A1(_00007_[0]),
    .A2(_08682_),
    .ZN(_08683_)
  );
  AND2_X1 _43092_ (
    .A1(_08675_),
    .A2(_08683_),
    .ZN(_08684_)
  );
  INV_X1 _43093_ (
    .A(_08684_),
    .ZN(_08685_)
  );
  AND2_X1 _43094_ (
    .A1(_08668_),
    .A2(_08685_),
    .ZN(_08686_)
  );
  INV_X1 _43095_ (
    .A(_08686_),
    .ZN(_08687_)
  );
  AND2_X1 _43096_ (
    .A1(_22144_),
    .A2(_08687_),
    .ZN(_08688_)
  );
  INV_X1 _43097_ (
    .A(_08688_),
    .ZN(_08689_)
  );
  AND2_X1 _43098_ (
    .A1(_00007_[3]),
    .A2(_08689_),
    .ZN(_08690_)
  );
  AND2_X1 _43099_ (
    .A1(_08651_),
    .A2(_08690_),
    .ZN(_08691_)
  );
  INV_X1 _43100_ (
    .A(_08691_),
    .ZN(_08692_)
  );
  AND2_X1 _43101_ (
    .A1(_22109_),
    .A2(_08613_),
    .ZN(_08693_)
  );
  INV_X1 _43102_ (
    .A(_08693_),
    .ZN(_08694_)
  );
  AND2_X1 _43103_ (
    .A1(_08692_),
    .A2(_08694_),
    .ZN(_08695_)
  );
  AND2_X1 _43104_ (
    .A1(_05842_),
    .A2(_08695_),
    .ZN(_08696_)
  );
  INV_X1 _43105_ (
    .A(_08696_),
    .ZN(_08697_)
  );
  AND2_X1 _43106_ (
    .A1(_21221_),
    .A2(_04963_),
    .ZN(_08698_)
  );
  INV_X1 _43107_ (
    .A(_08698_),
    .ZN(_08699_)
  );
  AND2_X1 _43108_ (
    .A1(_04962_),
    .A2(_08697_),
    .ZN(_08700_)
  );
  AND2_X1 _43109_ (
    .A1(_08534_),
    .A2(_08700_),
    .ZN(_08701_)
  );
  INV_X1 _43110_ (
    .A(_08701_),
    .ZN(_08702_)
  );
  AND2_X1 _43111_ (
    .A1(_08699_),
    .A2(_08702_),
    .ZN(_00302_)
  );
  AND2_X1 _43112_ (
    .A1(\cpuregs[29] [22]),
    .A2(_00007_[2]),
    .ZN(_08703_)
  );
  INV_X1 _43113_ (
    .A(_08703_),
    .ZN(_08704_)
  );
  AND2_X1 _43114_ (
    .A1(\cpuregs[25] [22]),
    .A2(_22077_),
    .ZN(_08705_)
  );
  INV_X1 _43115_ (
    .A(_08705_),
    .ZN(_08706_)
  );
  AND2_X1 _43116_ (
    .A1(_00007_[0]),
    .A2(_08706_),
    .ZN(_08707_)
  );
  AND2_X1 _43117_ (
    .A1(_08704_),
    .A2(_08707_),
    .ZN(_08708_)
  );
  INV_X1 _43118_ (
    .A(_08708_),
    .ZN(_08709_)
  );
  AND2_X1 _43119_ (
    .A1(\cpuregs[24] [22]),
    .A2(_22077_),
    .ZN(_08710_)
  );
  INV_X1 _43120_ (
    .A(_08710_),
    .ZN(_08711_)
  );
  AND2_X1 _43121_ (
    .A1(\cpuregs[28] [22]),
    .A2(_00007_[2]),
    .ZN(_08712_)
  );
  INV_X1 _43122_ (
    .A(_08712_),
    .ZN(_08713_)
  );
  AND2_X1 _43123_ (
    .A1(_22152_),
    .A2(_08713_),
    .ZN(_08714_)
  );
  AND2_X1 _43124_ (
    .A1(_08711_),
    .A2(_08714_),
    .ZN(_08715_)
  );
  INV_X1 _43125_ (
    .A(_08715_),
    .ZN(_08716_)
  );
  AND2_X1 _43126_ (
    .A1(_22078_),
    .A2(_08716_),
    .ZN(_08717_)
  );
  AND2_X1 _43127_ (
    .A1(_08709_),
    .A2(_08717_),
    .ZN(_08718_)
  );
  INV_X1 _43128_ (
    .A(_08718_),
    .ZN(_08719_)
  );
  AND2_X1 _43129_ (
    .A1(\cpuregs[31] [22]),
    .A2(_00007_[2]),
    .ZN(_08720_)
  );
  INV_X1 _43130_ (
    .A(_08720_),
    .ZN(_08721_)
  );
  AND2_X1 _43131_ (
    .A1(\cpuregs[27] [22]),
    .A2(_22077_),
    .ZN(_08722_)
  );
  INV_X1 _43132_ (
    .A(_08722_),
    .ZN(_08723_)
  );
  AND2_X1 _43133_ (
    .A1(_00007_[0]),
    .A2(_08723_),
    .ZN(_08724_)
  );
  AND2_X1 _43134_ (
    .A1(_08721_),
    .A2(_08724_),
    .ZN(_08725_)
  );
  INV_X1 _43135_ (
    .A(_08725_),
    .ZN(_08726_)
  );
  AND2_X1 _43136_ (
    .A1(\cpuregs[26] [22]),
    .A2(_22077_),
    .ZN(_08727_)
  );
  INV_X1 _43137_ (
    .A(_08727_),
    .ZN(_08728_)
  );
  AND2_X1 _43138_ (
    .A1(\cpuregs[30] [22]),
    .A2(_00007_[2]),
    .ZN(_08729_)
  );
  INV_X1 _43139_ (
    .A(_08729_),
    .ZN(_08730_)
  );
  AND2_X1 _43140_ (
    .A1(_22152_),
    .A2(_08730_),
    .ZN(_08731_)
  );
  AND2_X1 _43141_ (
    .A1(_08728_),
    .A2(_08731_),
    .ZN(_08732_)
  );
  INV_X1 _43142_ (
    .A(_08732_),
    .ZN(_08733_)
  );
  AND2_X1 _43143_ (
    .A1(_00007_[1]),
    .A2(_08733_),
    .ZN(_08734_)
  );
  AND2_X1 _43144_ (
    .A1(_08726_),
    .A2(_08734_),
    .ZN(_08735_)
  );
  INV_X1 _43145_ (
    .A(_08735_),
    .ZN(_08736_)
  );
  AND2_X1 _43146_ (
    .A1(_08719_),
    .A2(_08736_),
    .ZN(_08737_)
  );
  INV_X1 _43147_ (
    .A(_08737_),
    .ZN(_08738_)
  );
  AND2_X1 _43148_ (
    .A1(\cpuregs[11] [22]),
    .A2(_22077_),
    .ZN(_08739_)
  );
  INV_X1 _43149_ (
    .A(_08739_),
    .ZN(_08740_)
  );
  AND2_X1 _43150_ (
    .A1(\cpuregs[15] [22]),
    .A2(_00007_[2]),
    .ZN(_08741_)
  );
  INV_X1 _43151_ (
    .A(_08741_),
    .ZN(_08742_)
  );
  AND2_X1 _43152_ (
    .A1(_08740_),
    .A2(_08742_),
    .ZN(_08743_)
  );
  INV_X1 _43153_ (
    .A(_08743_),
    .ZN(_08744_)
  );
  AND2_X1 _43154_ (
    .A1(_00007_[0]),
    .A2(_08744_),
    .ZN(_08745_)
  );
  INV_X1 _43155_ (
    .A(_08745_),
    .ZN(_08746_)
  );
  AND2_X1 _43156_ (
    .A1(\cpuregs[14] [22]),
    .A2(_00007_[2]),
    .ZN(_08747_)
  );
  INV_X1 _43157_ (
    .A(_08747_),
    .ZN(_08748_)
  );
  AND2_X1 _43158_ (
    .A1(\cpuregs[10] [22]),
    .A2(_22077_),
    .ZN(_08749_)
  );
  INV_X1 _43159_ (
    .A(_08749_),
    .ZN(_08750_)
  );
  AND2_X1 _43160_ (
    .A1(_08748_),
    .A2(_08750_),
    .ZN(_08751_)
  );
  INV_X1 _43161_ (
    .A(_08751_),
    .ZN(_08752_)
  );
  AND2_X1 _43162_ (
    .A1(_22152_),
    .A2(_08752_),
    .ZN(_08753_)
  );
  INV_X1 _43163_ (
    .A(_08753_),
    .ZN(_08754_)
  );
  AND2_X1 _43164_ (
    .A1(_08746_),
    .A2(_08754_),
    .ZN(_08755_)
  );
  AND2_X1 _43165_ (
    .A1(\cpuregs[9] [22]),
    .A2(_22077_),
    .ZN(_08756_)
  );
  INV_X1 _43166_ (
    .A(_08756_),
    .ZN(_08757_)
  );
  AND2_X1 _43167_ (
    .A1(\cpuregs[13] [22]),
    .A2(_00007_[2]),
    .ZN(_08758_)
  );
  INV_X1 _43168_ (
    .A(_08758_),
    .ZN(_08759_)
  );
  AND2_X1 _43169_ (
    .A1(_08757_),
    .A2(_08759_),
    .ZN(_08760_)
  );
  INV_X1 _43170_ (
    .A(_08760_),
    .ZN(_08761_)
  );
  AND2_X1 _43171_ (
    .A1(_00007_[0]),
    .A2(_08761_),
    .ZN(_08762_)
  );
  INV_X1 _43172_ (
    .A(_08762_),
    .ZN(_08763_)
  );
  AND2_X1 _43173_ (
    .A1(\cpuregs[12] [22]),
    .A2(_00007_[2]),
    .ZN(_08764_)
  );
  INV_X1 _43174_ (
    .A(_08764_),
    .ZN(_08765_)
  );
  AND2_X1 _43175_ (
    .A1(\cpuregs[8] [22]),
    .A2(_22077_),
    .ZN(_08766_)
  );
  INV_X1 _43176_ (
    .A(_08766_),
    .ZN(_08767_)
  );
  AND2_X1 _43177_ (
    .A1(_08765_),
    .A2(_08767_),
    .ZN(_08768_)
  );
  INV_X1 _43178_ (
    .A(_08768_),
    .ZN(_08769_)
  );
  AND2_X1 _43179_ (
    .A1(_22152_),
    .A2(_08769_),
    .ZN(_08770_)
  );
  INV_X1 _43180_ (
    .A(_08770_),
    .ZN(_08771_)
  );
  AND2_X1 _43181_ (
    .A1(_08763_),
    .A2(_08771_),
    .ZN(_08772_)
  );
  AND2_X1 _43182_ (
    .A1(_21452_),
    .A2(_22077_),
    .ZN(_08773_)
  );
  INV_X1 _43183_ (
    .A(_08773_),
    .ZN(_08774_)
  );
  AND2_X1 _43184_ (
    .A1(_21663_),
    .A2(_00007_[2]),
    .ZN(_08775_)
  );
  INV_X1 _43185_ (
    .A(_08775_),
    .ZN(_08776_)
  );
  AND2_X1 _43186_ (
    .A1(_08774_),
    .A2(_08776_),
    .ZN(_08777_)
  );
  AND2_X1 _43187_ (
    .A1(_21474_),
    .A2(_22077_),
    .ZN(_08778_)
  );
  INV_X1 _43188_ (
    .A(_08778_),
    .ZN(_08779_)
  );
  AND2_X1 _43189_ (
    .A1(_21773_),
    .A2(_00007_[2]),
    .ZN(_08780_)
  );
  INV_X1 _43190_ (
    .A(_08780_),
    .ZN(_08781_)
  );
  AND2_X1 _43191_ (
    .A1(_00007_[0]),
    .A2(_08781_),
    .ZN(_08782_)
  );
  AND2_X1 _43192_ (
    .A1(_08779_),
    .A2(_08782_),
    .ZN(_08783_)
  );
  INV_X1 _43193_ (
    .A(_08783_),
    .ZN(_08784_)
  );
  AND2_X1 _43194_ (
    .A1(_22152_),
    .A2(_08777_),
    .ZN(_08785_)
  );
  INV_X1 _43195_ (
    .A(_08785_),
    .ZN(_08786_)
  );
  AND2_X1 _43196_ (
    .A1(_08784_),
    .A2(_08786_),
    .ZN(_08787_)
  );
  AND2_X1 _43197_ (
    .A1(_21607_),
    .A2(_22077_),
    .ZN(_08788_)
  );
  INV_X1 _43198_ (
    .A(_08788_),
    .ZN(_08789_)
  );
  AND2_X1 _43199_ (
    .A1(_21427_),
    .A2(_00007_[2]),
    .ZN(_08790_)
  );
  INV_X1 _43200_ (
    .A(_08790_),
    .ZN(_08791_)
  );
  AND2_X1 _43201_ (
    .A1(_21386_),
    .A2(_00007_[2]),
    .ZN(_08792_)
  );
  INV_X1 _43202_ (
    .A(_08792_),
    .ZN(_08793_)
  );
  AND2_X1 _43203_ (
    .A1(_21632_),
    .A2(_22077_),
    .ZN(_08794_)
  );
  INV_X1 _43204_ (
    .A(_08794_),
    .ZN(_08795_)
  );
  AND2_X1 _43205_ (
    .A1(_22152_),
    .A2(_08791_),
    .ZN(_08796_)
  );
  AND2_X1 _43206_ (
    .A1(_08789_),
    .A2(_08796_),
    .ZN(_08797_)
  );
  INV_X1 _43207_ (
    .A(_08797_),
    .ZN(_08798_)
  );
  AND2_X1 _43208_ (
    .A1(_00007_[0]),
    .A2(_08793_),
    .ZN(_08799_)
  );
  AND2_X1 _43209_ (
    .A1(_08795_),
    .A2(_08799_),
    .ZN(_08800_)
  );
  INV_X1 _43210_ (
    .A(_08800_),
    .ZN(_08801_)
  );
  AND2_X1 _43211_ (
    .A1(_08798_),
    .A2(_08801_),
    .ZN(_08802_)
  );
  AND2_X1 _43212_ (
    .A1(_21558_),
    .A2(_22077_),
    .ZN(_08803_)
  );
  INV_X1 _43213_ (
    .A(_08803_),
    .ZN(_08804_)
  );
  AND2_X1 _43214_ (
    .A1(_21824_),
    .A2(_00007_[2]),
    .ZN(_08805_)
  );
  INV_X1 _43215_ (
    .A(_08805_),
    .ZN(_08806_)
  );
  AND2_X1 _43216_ (
    .A1(_22152_),
    .A2(_08806_),
    .ZN(_08807_)
  );
  AND2_X1 _43217_ (
    .A1(_08804_),
    .A2(_08807_),
    .ZN(_08808_)
  );
  INV_X1 _43218_ (
    .A(_08808_),
    .ZN(_08809_)
  );
  AND2_X1 _43219_ (
    .A1(\cpuregs[7] [22]),
    .A2(_00007_[2]),
    .ZN(_08810_)
  );
  INV_X1 _43220_ (
    .A(_08810_),
    .ZN(_08811_)
  );
  AND2_X1 _43221_ (
    .A1(\cpuregs[3] [22]),
    .A2(_22077_),
    .ZN(_08812_)
  );
  INV_X1 _43222_ (
    .A(_08812_),
    .ZN(_08813_)
  );
  AND2_X1 _43223_ (
    .A1(_08811_),
    .A2(_08813_),
    .ZN(_08814_)
  );
  INV_X1 _43224_ (
    .A(_08814_),
    .ZN(_08815_)
  );
  AND2_X1 _43225_ (
    .A1(_00007_[0]),
    .A2(_08815_),
    .ZN(_08816_)
  );
  INV_X1 _43226_ (
    .A(_08816_),
    .ZN(_08817_)
  );
  AND2_X1 _43227_ (
    .A1(_08809_),
    .A2(_08817_),
    .ZN(_08818_)
  );
  AND2_X1 _43228_ (
    .A1(\cpuregs[1] [22]),
    .A2(_22077_),
    .ZN(_08819_)
  );
  INV_X1 _43229_ (
    .A(_08819_),
    .ZN(_08820_)
  );
  AND2_X1 _43230_ (
    .A1(\cpuregs[5] [22]),
    .A2(_00007_[2]),
    .ZN(_08821_)
  );
  INV_X1 _43231_ (
    .A(_08821_),
    .ZN(_08822_)
  );
  AND2_X1 _43232_ (
    .A1(_08820_),
    .A2(_08822_),
    .ZN(_08823_)
  );
  INV_X1 _43233_ (
    .A(_08823_),
    .ZN(_08824_)
  );
  AND2_X1 _43234_ (
    .A1(_00007_[0]),
    .A2(_08824_),
    .ZN(_08825_)
  );
  INV_X1 _43235_ (
    .A(_08825_),
    .ZN(_08826_)
  );
  AND2_X1 _43236_ (
    .A1(\cpuregs[4] [22]),
    .A2(_00007_[2]),
    .ZN(_08827_)
  );
  INV_X1 _43237_ (
    .A(_08827_),
    .ZN(_08828_)
  );
  AND2_X1 _43238_ (
    .A1(\cpuregs[0] [22]),
    .A2(_22077_),
    .ZN(_08829_)
  );
  INV_X1 _43239_ (
    .A(_08829_),
    .ZN(_08830_)
  );
  AND2_X1 _43240_ (
    .A1(_08828_),
    .A2(_08830_),
    .ZN(_08831_)
  );
  INV_X1 _43241_ (
    .A(_08831_),
    .ZN(_08832_)
  );
  AND2_X1 _43242_ (
    .A1(_22152_),
    .A2(_08832_),
    .ZN(_08833_)
  );
  INV_X1 _43243_ (
    .A(_08833_),
    .ZN(_08834_)
  );
  AND2_X1 _43244_ (
    .A1(_08826_),
    .A2(_08834_),
    .ZN(_08835_)
  );
  AND2_X1 _43245_ (
    .A1(_00007_[1]),
    .A2(_08818_),
    .ZN(_08836_)
  );
  INV_X1 _43246_ (
    .A(_08836_),
    .ZN(_08837_)
  );
  AND2_X1 _43247_ (
    .A1(_22078_),
    .A2(_08835_),
    .ZN(_08838_)
  );
  INV_X1 _43248_ (
    .A(_08838_),
    .ZN(_08839_)
  );
  AND2_X1 _43249_ (
    .A1(_08837_),
    .A2(_08839_),
    .ZN(_08840_)
  );
  AND2_X1 _43250_ (
    .A1(_00007_[1]),
    .A2(_08802_),
    .ZN(_08841_)
  );
  INV_X1 _43251_ (
    .A(_08841_),
    .ZN(_08842_)
  );
  AND2_X1 _43252_ (
    .A1(_22078_),
    .A2(_08787_),
    .ZN(_08843_)
  );
  INV_X1 _43253_ (
    .A(_08843_),
    .ZN(_08844_)
  );
  AND2_X1 _43254_ (
    .A1(_22109_),
    .A2(_08844_),
    .ZN(_08845_)
  );
  AND2_X1 _43255_ (
    .A1(_08842_),
    .A2(_08845_),
    .ZN(_08846_)
  );
  INV_X1 _43256_ (
    .A(_08846_),
    .ZN(_08847_)
  );
  AND2_X1 _43257_ (
    .A1(_00007_[3]),
    .A2(_08738_),
    .ZN(_08848_)
  );
  INV_X1 _43258_ (
    .A(_08848_),
    .ZN(_08849_)
  );
  AND2_X1 _43259_ (
    .A1(_00007_[4]),
    .A2(_08849_),
    .ZN(_08850_)
  );
  AND2_X1 _43260_ (
    .A1(_08847_),
    .A2(_08850_),
    .ZN(_08851_)
  );
  INV_X1 _43261_ (
    .A(_08851_),
    .ZN(_08852_)
  );
  AND2_X1 _43262_ (
    .A1(_22109_),
    .A2(_08840_),
    .ZN(_08853_)
  );
  INV_X1 _43263_ (
    .A(_08853_),
    .ZN(_08854_)
  );
  AND2_X1 _43264_ (
    .A1(_00007_[1]),
    .A2(_08755_),
    .ZN(_08855_)
  );
  INV_X1 _43265_ (
    .A(_08855_),
    .ZN(_08856_)
  );
  AND2_X1 _43266_ (
    .A1(_22078_),
    .A2(_08772_),
    .ZN(_08857_)
  );
  INV_X1 _43267_ (
    .A(_08857_),
    .ZN(_08858_)
  );
  AND2_X1 _43268_ (
    .A1(_00007_[3]),
    .A2(_08858_),
    .ZN(_08859_)
  );
  AND2_X1 _43269_ (
    .A1(_08856_),
    .A2(_08859_),
    .ZN(_08860_)
  );
  INV_X1 _43270_ (
    .A(_08860_),
    .ZN(_08861_)
  );
  AND2_X1 _43271_ (
    .A1(_08854_),
    .A2(_08861_),
    .ZN(_08862_)
  );
  AND2_X1 _43272_ (
    .A1(_22144_),
    .A2(_08862_),
    .ZN(_08863_)
  );
  INV_X1 _43273_ (
    .A(_08863_),
    .ZN(_08864_)
  );
  AND2_X1 _43274_ (
    .A1(_08852_),
    .A2(_08864_),
    .ZN(_08865_)
  );
  AND2_X1 _43275_ (
    .A1(_05842_),
    .A2(_08865_),
    .ZN(_08866_)
  );
  INV_X1 _43276_ (
    .A(_08866_),
    .ZN(_08867_)
  );
  AND2_X1 _43277_ (
    .A1(decoded_imm[22]),
    .A2(_04966_),
    .ZN(_08868_)
  );
  INV_X1 _43278_ (
    .A(_08868_),
    .ZN(_08869_)
  );
  AND2_X1 _43279_ (
    .A1(_21222_),
    .A2(_04963_),
    .ZN(_08870_)
  );
  INV_X1 _43280_ (
    .A(_08870_),
    .ZN(_08871_)
  );
  AND2_X1 _43281_ (
    .A1(_04962_),
    .A2(_08869_),
    .ZN(_08872_)
  );
  AND2_X1 _43282_ (
    .A1(_08867_),
    .A2(_08872_),
    .ZN(_08873_)
  );
  INV_X1 _43283_ (
    .A(_08873_),
    .ZN(_08874_)
  );
  AND2_X1 _43284_ (
    .A1(_08871_),
    .A2(_08874_),
    .ZN(_00303_)
  );
  AND2_X1 _43285_ (
    .A1(decoded_imm[23]),
    .A2(_04966_),
    .ZN(_08875_)
  );
  INV_X1 _43286_ (
    .A(_08875_),
    .ZN(_08876_)
  );
  AND2_X1 _43287_ (
    .A1(_21633_),
    .A2(_22077_),
    .ZN(_08877_)
  );
  INV_X1 _43288_ (
    .A(_08877_),
    .ZN(_08878_)
  );
  AND2_X1 _43289_ (
    .A1(_21387_),
    .A2(_00007_[2]),
    .ZN(_08879_)
  );
  INV_X1 _43290_ (
    .A(_08879_),
    .ZN(_08880_)
  );
  AND2_X1 _43291_ (
    .A1(_00007_[0]),
    .A2(_08878_),
    .ZN(_08881_)
  );
  AND2_X1 _43292_ (
    .A1(_08880_),
    .A2(_08881_),
    .ZN(_08882_)
  );
  INV_X1 _43293_ (
    .A(_08882_),
    .ZN(_08883_)
  );
  AND2_X1 _43294_ (
    .A1(_21608_),
    .A2(_22077_),
    .ZN(_08884_)
  );
  INV_X1 _43295_ (
    .A(_08884_),
    .ZN(_08885_)
  );
  AND2_X1 _43296_ (
    .A1(_21428_),
    .A2(_00007_[2]),
    .ZN(_08886_)
  );
  INV_X1 _43297_ (
    .A(_08886_),
    .ZN(_08887_)
  );
  AND2_X1 _43298_ (
    .A1(_22152_),
    .A2(_08887_),
    .ZN(_08888_)
  );
  AND2_X1 _43299_ (
    .A1(_08885_),
    .A2(_08888_),
    .ZN(_08889_)
  );
  INV_X1 _43300_ (
    .A(_08889_),
    .ZN(_08890_)
  );
  AND2_X1 _43301_ (
    .A1(_21505_),
    .A2(_22077_),
    .ZN(_08891_)
  );
  INV_X1 _43302_ (
    .A(_08891_),
    .ZN(_08892_)
  );
  AND2_X1 _43303_ (
    .A1(_21797_),
    .A2(_00007_[2]),
    .ZN(_08893_)
  );
  INV_X1 _43304_ (
    .A(_08893_),
    .ZN(_08894_)
  );
  AND2_X1 _43305_ (
    .A1(_00007_[0]),
    .A2(_08894_),
    .ZN(_08895_)
  );
  AND2_X1 _43306_ (
    .A1(_08892_),
    .A2(_08895_),
    .ZN(_08896_)
  );
  INV_X1 _43307_ (
    .A(_08896_),
    .ZN(_08897_)
  );
  AND2_X1 _43308_ (
    .A1(_21825_),
    .A2(_00007_[2]),
    .ZN(_08898_)
  );
  INV_X1 _43309_ (
    .A(_08898_),
    .ZN(_08899_)
  );
  AND2_X1 _43310_ (
    .A1(_21559_),
    .A2(_22077_),
    .ZN(_08900_)
  );
  INV_X1 _43311_ (
    .A(_08900_),
    .ZN(_08901_)
  );
  AND2_X1 _43312_ (
    .A1(_22152_),
    .A2(_08901_),
    .ZN(_08902_)
  );
  AND2_X1 _43313_ (
    .A1(_08899_),
    .A2(_08902_),
    .ZN(_08903_)
  );
  INV_X1 _43314_ (
    .A(_08903_),
    .ZN(_08904_)
  );
  AND2_X1 _43315_ (
    .A1(\cpuregs[17] [23]),
    .A2(_22077_),
    .ZN(_08905_)
  );
  INV_X1 _43316_ (
    .A(_08905_),
    .ZN(_08906_)
  );
  AND2_X1 _43317_ (
    .A1(\cpuregs[21] [23]),
    .A2(_00007_[2]),
    .ZN(_08907_)
  );
  INV_X1 _43318_ (
    .A(_08907_),
    .ZN(_08908_)
  );
  AND2_X1 _43319_ (
    .A1(_08906_),
    .A2(_08908_),
    .ZN(_08909_)
  );
  INV_X1 _43320_ (
    .A(_08909_),
    .ZN(_08910_)
  );
  AND2_X1 _43321_ (
    .A1(_00007_[0]),
    .A2(_08910_),
    .ZN(_08911_)
  );
  INV_X1 _43322_ (
    .A(_08911_),
    .ZN(_08912_)
  );
  AND2_X1 _43323_ (
    .A1(\cpuregs[16] [23]),
    .A2(_22077_),
    .ZN(_08913_)
  );
  INV_X1 _43324_ (
    .A(_08913_),
    .ZN(_08914_)
  );
  AND2_X1 _43325_ (
    .A1(\cpuregs[20] [23]),
    .A2(_00007_[2]),
    .ZN(_08915_)
  );
  INV_X1 _43326_ (
    .A(_08915_),
    .ZN(_08916_)
  );
  AND2_X1 _43327_ (
    .A1(_08914_),
    .A2(_08916_),
    .ZN(_08917_)
  );
  INV_X1 _43328_ (
    .A(_08917_),
    .ZN(_08918_)
  );
  AND2_X1 _43329_ (
    .A1(_22152_),
    .A2(_08918_),
    .ZN(_08919_)
  );
  INV_X1 _43330_ (
    .A(_08919_),
    .ZN(_08920_)
  );
  AND2_X1 _43331_ (
    .A1(_08912_),
    .A2(_08920_),
    .ZN(_08921_)
  );
  AND2_X1 _43332_ (
    .A1(_21530_),
    .A2(_22077_),
    .ZN(_08922_)
  );
  INV_X1 _43333_ (
    .A(_08922_),
    .ZN(_08923_)
  );
  AND2_X1 _43334_ (
    .A1(_21750_),
    .A2(_00007_[2]),
    .ZN(_08924_)
  );
  INV_X1 _43335_ (
    .A(_08924_),
    .ZN(_08925_)
  );
  AND2_X1 _43336_ (
    .A1(_00007_[0]),
    .A2(_08925_),
    .ZN(_08926_)
  );
  AND2_X1 _43337_ (
    .A1(_08923_),
    .A2(_08926_),
    .ZN(_08927_)
  );
  INV_X1 _43338_ (
    .A(_08927_),
    .ZN(_08928_)
  );
  AND2_X1 _43339_ (
    .A1(_21971_),
    .A2(_22077_),
    .ZN(_08929_)
  );
  INV_X1 _43340_ (
    .A(_08929_),
    .ZN(_08930_)
  );
  AND2_X1 _43341_ (
    .A1(_21687_),
    .A2(_00007_[2]),
    .ZN(_08931_)
  );
  INV_X1 _43342_ (
    .A(_08931_),
    .ZN(_08932_)
  );
  AND2_X1 _43343_ (
    .A1(_08930_),
    .A2(_08932_),
    .ZN(_08933_)
  );
  AND2_X1 _43344_ (
    .A1(_22152_),
    .A2(_08933_),
    .ZN(_08934_)
  );
  INV_X1 _43345_ (
    .A(_08934_),
    .ZN(_08935_)
  );
  AND2_X1 _43346_ (
    .A1(_08928_),
    .A2(_08935_),
    .ZN(_08936_)
  );
  AND2_X1 _43347_ (
    .A1(_22078_),
    .A2(_08936_),
    .ZN(_08937_)
  );
  INV_X1 _43348_ (
    .A(_08937_),
    .ZN(_08938_)
  );
  AND2_X1 _43349_ (
    .A1(_00007_[1]),
    .A2(_08904_),
    .ZN(_08939_)
  );
  AND2_X1 _43350_ (
    .A1(_08897_),
    .A2(_08939_),
    .ZN(_08940_)
  );
  INV_X1 _43351_ (
    .A(_08940_),
    .ZN(_08941_)
  );
  AND2_X1 _43352_ (
    .A1(_08938_),
    .A2(_08941_),
    .ZN(_08942_)
  );
  AND2_X1 _43353_ (
    .A1(_22144_),
    .A2(_08942_),
    .ZN(_08943_)
  );
  INV_X1 _43354_ (
    .A(_08943_),
    .ZN(_08944_)
  );
  AND2_X1 _43355_ (
    .A1(_00007_[1]),
    .A2(_08890_),
    .ZN(_08945_)
  );
  AND2_X1 _43356_ (
    .A1(_08883_),
    .A2(_08945_),
    .ZN(_08946_)
  );
  INV_X1 _43357_ (
    .A(_08946_),
    .ZN(_08947_)
  );
  AND2_X1 _43358_ (
    .A1(_22078_),
    .A2(_08921_),
    .ZN(_08948_)
  );
  INV_X1 _43359_ (
    .A(_08948_),
    .ZN(_08949_)
  );
  AND2_X1 _43360_ (
    .A1(_08947_),
    .A2(_08949_),
    .ZN(_08950_)
  );
  AND2_X1 _43361_ (
    .A1(_00007_[4]),
    .A2(_08950_),
    .ZN(_08951_)
  );
  INV_X1 _43362_ (
    .A(_08951_),
    .ZN(_08952_)
  );
  AND2_X1 _43363_ (
    .A1(_08944_),
    .A2(_08952_),
    .ZN(_08953_)
  );
  AND2_X1 _43364_ (
    .A1(_21860_),
    .A2(_00007_[2]),
    .ZN(_08954_)
  );
  INV_X1 _43365_ (
    .A(_08954_),
    .ZN(_08955_)
  );
  AND2_X1 _43366_ (
    .A1(_21882_),
    .A2(_22077_),
    .ZN(_08956_)
  );
  INV_X1 _43367_ (
    .A(_08956_),
    .ZN(_08957_)
  );
  AND2_X1 _43368_ (
    .A1(_08955_),
    .A2(_08957_),
    .ZN(_08958_)
  );
  AND2_X1 _43369_ (
    .A1(_22152_),
    .A2(_08958_),
    .ZN(_08959_)
  );
  INV_X1 _43370_ (
    .A(_08959_),
    .ZN(_08960_)
  );
  AND2_X1 _43371_ (
    .A1(_21932_),
    .A2(_22077_),
    .ZN(_08961_)
  );
  INV_X1 _43372_ (
    .A(_08961_),
    .ZN(_08962_)
  );
  AND2_X1 _43373_ (
    .A1(_21948_),
    .A2(_00007_[2]),
    .ZN(_08963_)
  );
  INV_X1 _43374_ (
    .A(_08963_),
    .ZN(_08964_)
  );
  AND2_X1 _43375_ (
    .A1(_00007_[0]),
    .A2(_08964_),
    .ZN(_08965_)
  );
  AND2_X1 _43376_ (
    .A1(_08962_),
    .A2(_08965_),
    .ZN(_08966_)
  );
  INV_X1 _43377_ (
    .A(_08966_),
    .ZN(_08967_)
  );
  AND2_X1 _43378_ (
    .A1(_00007_[1]),
    .A2(_08967_),
    .ZN(_08968_)
  );
  AND2_X1 _43379_ (
    .A1(_08960_),
    .A2(_08968_),
    .ZN(_08969_)
  );
  INV_X1 _43380_ (
    .A(_08969_),
    .ZN(_08970_)
  );
  AND2_X1 _43381_ (
    .A1(_21900_),
    .A2(_00007_[2]),
    .ZN(_08971_)
  );
  INV_X1 _43382_ (
    .A(_08971_),
    .ZN(_08972_)
  );
  AND2_X1 _43383_ (
    .A1(_21844_),
    .A2(_22077_),
    .ZN(_08973_)
  );
  INV_X1 _43384_ (
    .A(_08973_),
    .ZN(_08974_)
  );
  AND2_X1 _43385_ (
    .A1(_00007_[0]),
    .A2(_08974_),
    .ZN(_08975_)
  );
  AND2_X1 _43386_ (
    .A1(_08972_),
    .A2(_08975_),
    .ZN(_08976_)
  );
  INV_X1 _43387_ (
    .A(_08976_),
    .ZN(_08977_)
  );
  AND2_X1 _43388_ (
    .A1(_21578_),
    .A2(_22077_),
    .ZN(_08978_)
  );
  INV_X1 _43389_ (
    .A(_08978_),
    .ZN(_08979_)
  );
  AND2_X1 _43390_ (
    .A1(_21916_),
    .A2(_00007_[2]),
    .ZN(_08980_)
  );
  INV_X1 _43391_ (
    .A(_08980_),
    .ZN(_08981_)
  );
  AND2_X1 _43392_ (
    .A1(_08979_),
    .A2(_08981_),
    .ZN(_08982_)
  );
  AND2_X1 _43393_ (
    .A1(_22152_),
    .A2(_08982_),
    .ZN(_08983_)
  );
  INV_X1 _43394_ (
    .A(_08983_),
    .ZN(_08984_)
  );
  AND2_X1 _43395_ (
    .A1(_08977_),
    .A2(_08984_),
    .ZN(_08985_)
  );
  AND2_X1 _43396_ (
    .A1(_22078_),
    .A2(_08985_),
    .ZN(_08986_)
  );
  INV_X1 _43397_ (
    .A(_08986_),
    .ZN(_08987_)
  );
  AND2_X1 _43398_ (
    .A1(_08970_),
    .A2(_08987_),
    .ZN(_08988_)
  );
  AND2_X1 _43399_ (
    .A1(_00007_[4]),
    .A2(_08988_),
    .ZN(_08989_)
  );
  INV_X1 _43400_ (
    .A(_08989_),
    .ZN(_08990_)
  );
  AND2_X1 _43401_ (
    .A1(_21644_),
    .A2(_00007_[2]),
    .ZN(_08991_)
  );
  INV_X1 _43402_ (
    .A(_08991_),
    .ZN(_08992_)
  );
  AND2_X1 _43403_ (
    .A1(_21722_),
    .A2(_22077_),
    .ZN(_08993_)
  );
  INV_X1 _43404_ (
    .A(_08993_),
    .ZN(_08994_)
  );
  AND2_X1 _43405_ (
    .A1(_00007_[0]),
    .A2(_08994_),
    .ZN(_08995_)
  );
  AND2_X1 _43406_ (
    .A1(_08992_),
    .A2(_08995_),
    .ZN(_08996_)
  );
  INV_X1 _43407_ (
    .A(_08996_),
    .ZN(_08997_)
  );
  AND2_X1 _43408_ (
    .A1(_21729_),
    .A2(_22077_),
    .ZN(_08998_)
  );
  INV_X1 _43409_ (
    .A(_08998_),
    .ZN(_08999_)
  );
  AND2_X1 _43410_ (
    .A1(_21484_),
    .A2(_00007_[2]),
    .ZN(_09000_)
  );
  INV_X1 _43411_ (
    .A(_09000_),
    .ZN(_09001_)
  );
  AND2_X1 _43412_ (
    .A1(_08999_),
    .A2(_09001_),
    .ZN(_09002_)
  );
  AND2_X1 _43413_ (
    .A1(_22152_),
    .A2(_09002_),
    .ZN(_09003_)
  );
  INV_X1 _43414_ (
    .A(_09003_),
    .ZN(_09004_)
  );
  AND2_X1 _43415_ (
    .A1(_08997_),
    .A2(_09004_),
    .ZN(_09005_)
  );
  AND2_X1 _43416_ (
    .A1(_22078_),
    .A2(_09005_),
    .ZN(_09006_)
  );
  INV_X1 _43417_ (
    .A(_09006_),
    .ZN(_09007_)
  );
  AND2_X1 _43418_ (
    .A1(_21398_),
    .A2(_00007_[2]),
    .ZN(_09008_)
  );
  INV_X1 _43419_ (
    .A(_09008_),
    .ZN(_09009_)
  );
  AND2_X1 _43420_ (
    .A1(_21710_),
    .A2(_22077_),
    .ZN(_09010_)
  );
  INV_X1 _43421_ (
    .A(_09010_),
    .ZN(_09011_)
  );
  AND2_X1 _43422_ (
    .A1(_09009_),
    .A2(_09011_),
    .ZN(_09012_)
  );
  AND2_X1 _43423_ (
    .A1(_22152_),
    .A2(_09012_),
    .ZN(_09013_)
  );
  INV_X1 _43424_ (
    .A(_09013_),
    .ZN(_09014_)
  );
  AND2_X1 _43425_ (
    .A1(_21587_),
    .A2(_22077_),
    .ZN(_09015_)
  );
  INV_X1 _43426_ (
    .A(_09015_),
    .ZN(_09016_)
  );
  AND2_X1 _43427_ (
    .A1(_21405_),
    .A2(_00007_[2]),
    .ZN(_09017_)
  );
  INV_X1 _43428_ (
    .A(_09017_),
    .ZN(_09018_)
  );
  AND2_X1 _43429_ (
    .A1(_00007_[0]),
    .A2(_09018_),
    .ZN(_09019_)
  );
  AND2_X1 _43430_ (
    .A1(_09016_),
    .A2(_09019_),
    .ZN(_09020_)
  );
  INV_X1 _43431_ (
    .A(_09020_),
    .ZN(_09021_)
  );
  AND2_X1 _43432_ (
    .A1(_00007_[1]),
    .A2(_09021_),
    .ZN(_09022_)
  );
  AND2_X1 _43433_ (
    .A1(_09014_),
    .A2(_09022_),
    .ZN(_09023_)
  );
  INV_X1 _43434_ (
    .A(_09023_),
    .ZN(_09024_)
  );
  AND2_X1 _43435_ (
    .A1(_09007_),
    .A2(_09024_),
    .ZN(_09025_)
  );
  AND2_X1 _43436_ (
    .A1(_22144_),
    .A2(_09025_),
    .ZN(_09026_)
  );
  INV_X1 _43437_ (
    .A(_09026_),
    .ZN(_09027_)
  );
  AND2_X1 _43438_ (
    .A1(_00007_[3]),
    .A2(_09027_),
    .ZN(_09028_)
  );
  AND2_X1 _43439_ (
    .A1(_08990_),
    .A2(_09028_),
    .ZN(_09029_)
  );
  INV_X1 _43440_ (
    .A(_09029_),
    .ZN(_09030_)
  );
  AND2_X1 _43441_ (
    .A1(_22109_),
    .A2(_08953_),
    .ZN(_09031_)
  );
  INV_X1 _43442_ (
    .A(_09031_),
    .ZN(_09032_)
  );
  AND2_X1 _43443_ (
    .A1(_09030_),
    .A2(_09032_),
    .ZN(_09033_)
  );
  AND2_X1 _43444_ (
    .A1(_05842_),
    .A2(_09033_),
    .ZN(_09034_)
  );
  INV_X1 _43445_ (
    .A(_09034_),
    .ZN(_09035_)
  );
  AND2_X1 _43446_ (
    .A1(_21223_),
    .A2(_04963_),
    .ZN(_09036_)
  );
  INV_X1 _43447_ (
    .A(_09036_),
    .ZN(_09037_)
  );
  AND2_X1 _43448_ (
    .A1(_04962_),
    .A2(_09035_),
    .ZN(_09038_)
  );
  AND2_X1 _43449_ (
    .A1(_08876_),
    .A2(_09038_),
    .ZN(_09039_)
  );
  INV_X1 _43450_ (
    .A(_09039_),
    .ZN(_09040_)
  );
  AND2_X1 _43451_ (
    .A1(_09037_),
    .A2(_09040_),
    .ZN(_00304_)
  );
  AND2_X1 _43452_ (
    .A1(decoded_imm[24]),
    .A2(_04966_),
    .ZN(_09041_)
  );
  INV_X1 _43453_ (
    .A(_09041_),
    .ZN(_09042_)
  );
  AND2_X1 _43454_ (
    .A1(\cpuregs[29] [24]),
    .A2(_00007_[2]),
    .ZN(_09043_)
  );
  INV_X1 _43455_ (
    .A(_09043_),
    .ZN(_09044_)
  );
  AND2_X1 _43456_ (
    .A1(\cpuregs[25] [24]),
    .A2(_22077_),
    .ZN(_09045_)
  );
  INV_X1 _43457_ (
    .A(_09045_),
    .ZN(_09046_)
  );
  AND2_X1 _43458_ (
    .A1(_00007_[0]),
    .A2(_09046_),
    .ZN(_09047_)
  );
  AND2_X1 _43459_ (
    .A1(_09044_),
    .A2(_09047_),
    .ZN(_09048_)
  );
  INV_X1 _43460_ (
    .A(_09048_),
    .ZN(_09049_)
  );
  AND2_X1 _43461_ (
    .A1(\cpuregs[24] [24]),
    .A2(_22077_),
    .ZN(_09050_)
  );
  INV_X1 _43462_ (
    .A(_09050_),
    .ZN(_09051_)
  );
  AND2_X1 _43463_ (
    .A1(\cpuregs[28] [24]),
    .A2(_00007_[2]),
    .ZN(_09052_)
  );
  INV_X1 _43464_ (
    .A(_09052_),
    .ZN(_09053_)
  );
  AND2_X1 _43465_ (
    .A1(_22152_),
    .A2(_09053_),
    .ZN(_09054_)
  );
  AND2_X1 _43466_ (
    .A1(_09051_),
    .A2(_09054_),
    .ZN(_09055_)
  );
  INV_X1 _43467_ (
    .A(_09055_),
    .ZN(_09056_)
  );
  AND2_X1 _43468_ (
    .A1(_22078_),
    .A2(_09056_),
    .ZN(_09057_)
  );
  AND2_X1 _43469_ (
    .A1(_09049_),
    .A2(_09057_),
    .ZN(_09058_)
  );
  INV_X1 _43470_ (
    .A(_09058_),
    .ZN(_09059_)
  );
  AND2_X1 _43471_ (
    .A1(\cpuregs[31] [24]),
    .A2(_00007_[2]),
    .ZN(_09060_)
  );
  INV_X1 _43472_ (
    .A(_09060_),
    .ZN(_09061_)
  );
  AND2_X1 _43473_ (
    .A1(\cpuregs[27] [24]),
    .A2(_22077_),
    .ZN(_09062_)
  );
  INV_X1 _43474_ (
    .A(_09062_),
    .ZN(_09063_)
  );
  AND2_X1 _43475_ (
    .A1(_00007_[0]),
    .A2(_09063_),
    .ZN(_09064_)
  );
  AND2_X1 _43476_ (
    .A1(_09061_),
    .A2(_09064_),
    .ZN(_09065_)
  );
  INV_X1 _43477_ (
    .A(_09065_),
    .ZN(_09066_)
  );
  AND2_X1 _43478_ (
    .A1(\cpuregs[26] [24]),
    .A2(_22077_),
    .ZN(_09067_)
  );
  INV_X1 _43479_ (
    .A(_09067_),
    .ZN(_09068_)
  );
  AND2_X1 _43480_ (
    .A1(\cpuregs[30] [24]),
    .A2(_00007_[2]),
    .ZN(_09069_)
  );
  INV_X1 _43481_ (
    .A(_09069_),
    .ZN(_09070_)
  );
  AND2_X1 _43482_ (
    .A1(_22152_),
    .A2(_09070_),
    .ZN(_09071_)
  );
  AND2_X1 _43483_ (
    .A1(_09068_),
    .A2(_09071_),
    .ZN(_09072_)
  );
  INV_X1 _43484_ (
    .A(_09072_),
    .ZN(_09073_)
  );
  AND2_X1 _43485_ (
    .A1(_00007_[1]),
    .A2(_09073_),
    .ZN(_09074_)
  );
  AND2_X1 _43486_ (
    .A1(_09066_),
    .A2(_09074_),
    .ZN(_09075_)
  );
  INV_X1 _43487_ (
    .A(_09075_),
    .ZN(_09076_)
  );
  AND2_X1 _43488_ (
    .A1(_09059_),
    .A2(_09076_),
    .ZN(_09077_)
  );
  INV_X1 _43489_ (
    .A(_09077_),
    .ZN(_09078_)
  );
  AND2_X1 _43490_ (
    .A1(\cpuregs[11] [24]),
    .A2(_22077_),
    .ZN(_09079_)
  );
  INV_X1 _43491_ (
    .A(_09079_),
    .ZN(_09080_)
  );
  AND2_X1 _43492_ (
    .A1(\cpuregs[15] [24]),
    .A2(_00007_[2]),
    .ZN(_09081_)
  );
  INV_X1 _43493_ (
    .A(_09081_),
    .ZN(_09082_)
  );
  AND2_X1 _43494_ (
    .A1(_09080_),
    .A2(_09082_),
    .ZN(_09083_)
  );
  INV_X1 _43495_ (
    .A(_09083_),
    .ZN(_09084_)
  );
  AND2_X1 _43496_ (
    .A1(_00007_[0]),
    .A2(_09084_),
    .ZN(_09085_)
  );
  INV_X1 _43497_ (
    .A(_09085_),
    .ZN(_09086_)
  );
  AND2_X1 _43498_ (
    .A1(\cpuregs[14] [24]),
    .A2(_00007_[2]),
    .ZN(_09087_)
  );
  INV_X1 _43499_ (
    .A(_09087_),
    .ZN(_09088_)
  );
  AND2_X1 _43500_ (
    .A1(\cpuregs[10] [24]),
    .A2(_22077_),
    .ZN(_09089_)
  );
  INV_X1 _43501_ (
    .A(_09089_),
    .ZN(_09090_)
  );
  AND2_X1 _43502_ (
    .A1(_09088_),
    .A2(_09090_),
    .ZN(_09091_)
  );
  INV_X1 _43503_ (
    .A(_09091_),
    .ZN(_09092_)
  );
  AND2_X1 _43504_ (
    .A1(_22152_),
    .A2(_09092_),
    .ZN(_09093_)
  );
  INV_X1 _43505_ (
    .A(_09093_),
    .ZN(_09094_)
  );
  AND2_X1 _43506_ (
    .A1(_09086_),
    .A2(_09094_),
    .ZN(_09095_)
  );
  AND2_X1 _43507_ (
    .A1(\cpuregs[9] [24]),
    .A2(_22077_),
    .ZN(_09096_)
  );
  INV_X1 _43508_ (
    .A(_09096_),
    .ZN(_09097_)
  );
  AND2_X1 _43509_ (
    .A1(\cpuregs[13] [24]),
    .A2(_00007_[2]),
    .ZN(_09098_)
  );
  INV_X1 _43510_ (
    .A(_09098_),
    .ZN(_09099_)
  );
  AND2_X1 _43511_ (
    .A1(_09097_),
    .A2(_09099_),
    .ZN(_09100_)
  );
  INV_X1 _43512_ (
    .A(_09100_),
    .ZN(_09101_)
  );
  AND2_X1 _43513_ (
    .A1(_00007_[0]),
    .A2(_09101_),
    .ZN(_09102_)
  );
  INV_X1 _43514_ (
    .A(_09102_),
    .ZN(_09103_)
  );
  AND2_X1 _43515_ (
    .A1(\cpuregs[12] [24]),
    .A2(_00007_[2]),
    .ZN(_09104_)
  );
  INV_X1 _43516_ (
    .A(_09104_),
    .ZN(_09105_)
  );
  AND2_X1 _43517_ (
    .A1(\cpuregs[8] [24]),
    .A2(_22077_),
    .ZN(_09106_)
  );
  INV_X1 _43518_ (
    .A(_09106_),
    .ZN(_09107_)
  );
  AND2_X1 _43519_ (
    .A1(_09105_),
    .A2(_09107_),
    .ZN(_09108_)
  );
  INV_X1 _43520_ (
    .A(_09108_),
    .ZN(_09109_)
  );
  AND2_X1 _43521_ (
    .A1(_22152_),
    .A2(_09109_),
    .ZN(_09110_)
  );
  INV_X1 _43522_ (
    .A(_09110_),
    .ZN(_09111_)
  );
  AND2_X1 _43523_ (
    .A1(_09103_),
    .A2(_09111_),
    .ZN(_09112_)
  );
  AND2_X1 _43524_ (
    .A1(_21453_),
    .A2(_22077_),
    .ZN(_09113_)
  );
  INV_X1 _43525_ (
    .A(_09113_),
    .ZN(_09114_)
  );
  AND2_X1 _43526_ (
    .A1(_21664_),
    .A2(_00007_[2]),
    .ZN(_09115_)
  );
  INV_X1 _43527_ (
    .A(_09115_),
    .ZN(_09116_)
  );
  AND2_X1 _43528_ (
    .A1(_09114_),
    .A2(_09116_),
    .ZN(_09117_)
  );
  AND2_X1 _43529_ (
    .A1(_21475_),
    .A2(_22077_),
    .ZN(_09118_)
  );
  INV_X1 _43530_ (
    .A(_09118_),
    .ZN(_09119_)
  );
  AND2_X1 _43531_ (
    .A1(_21774_),
    .A2(_00007_[2]),
    .ZN(_09120_)
  );
  INV_X1 _43532_ (
    .A(_09120_),
    .ZN(_09121_)
  );
  AND2_X1 _43533_ (
    .A1(_00007_[0]),
    .A2(_09121_),
    .ZN(_09122_)
  );
  AND2_X1 _43534_ (
    .A1(_09119_),
    .A2(_09122_),
    .ZN(_09123_)
  );
  INV_X1 _43535_ (
    .A(_09123_),
    .ZN(_09124_)
  );
  AND2_X1 _43536_ (
    .A1(_22152_),
    .A2(_09117_),
    .ZN(_09125_)
  );
  INV_X1 _43537_ (
    .A(_09125_),
    .ZN(_09126_)
  );
  AND2_X1 _43538_ (
    .A1(_09124_),
    .A2(_09126_),
    .ZN(_09127_)
  );
  AND2_X1 _43539_ (
    .A1(_21609_),
    .A2(_22077_),
    .ZN(_09128_)
  );
  INV_X1 _43540_ (
    .A(_09128_),
    .ZN(_09129_)
  );
  AND2_X1 _43541_ (
    .A1(_21429_),
    .A2(_00007_[2]),
    .ZN(_09130_)
  );
  INV_X1 _43542_ (
    .A(_09130_),
    .ZN(_09131_)
  );
  AND2_X1 _43543_ (
    .A1(_21388_),
    .A2(_00007_[2]),
    .ZN(_09132_)
  );
  INV_X1 _43544_ (
    .A(_09132_),
    .ZN(_09133_)
  );
  AND2_X1 _43545_ (
    .A1(_21634_),
    .A2(_22077_),
    .ZN(_09134_)
  );
  INV_X1 _43546_ (
    .A(_09134_),
    .ZN(_09135_)
  );
  AND2_X1 _43547_ (
    .A1(_22152_),
    .A2(_09131_),
    .ZN(_09136_)
  );
  AND2_X1 _43548_ (
    .A1(_09129_),
    .A2(_09136_),
    .ZN(_09137_)
  );
  INV_X1 _43549_ (
    .A(_09137_),
    .ZN(_09138_)
  );
  AND2_X1 _43550_ (
    .A1(_00007_[0]),
    .A2(_09133_),
    .ZN(_09139_)
  );
  AND2_X1 _43551_ (
    .A1(_09135_),
    .A2(_09139_),
    .ZN(_09140_)
  );
  INV_X1 _43552_ (
    .A(_09140_),
    .ZN(_09141_)
  );
  AND2_X1 _43553_ (
    .A1(_09138_),
    .A2(_09141_),
    .ZN(_09142_)
  );
  AND2_X1 _43554_ (
    .A1(_21560_),
    .A2(_22077_),
    .ZN(_09143_)
  );
  INV_X1 _43555_ (
    .A(_09143_),
    .ZN(_09144_)
  );
  AND2_X1 _43556_ (
    .A1(_21826_),
    .A2(_00007_[2]),
    .ZN(_09145_)
  );
  INV_X1 _43557_ (
    .A(_09145_),
    .ZN(_09146_)
  );
  AND2_X1 _43558_ (
    .A1(_22152_),
    .A2(_09146_),
    .ZN(_09147_)
  );
  AND2_X1 _43559_ (
    .A1(_09144_),
    .A2(_09147_),
    .ZN(_09148_)
  );
  INV_X1 _43560_ (
    .A(_09148_),
    .ZN(_09149_)
  );
  AND2_X1 _43561_ (
    .A1(\cpuregs[7] [24]),
    .A2(_00007_[2]),
    .ZN(_09150_)
  );
  INV_X1 _43562_ (
    .A(_09150_),
    .ZN(_09151_)
  );
  AND2_X1 _43563_ (
    .A1(\cpuregs[3] [24]),
    .A2(_22077_),
    .ZN(_09152_)
  );
  INV_X1 _43564_ (
    .A(_09152_),
    .ZN(_09153_)
  );
  AND2_X1 _43565_ (
    .A1(_09151_),
    .A2(_09153_),
    .ZN(_09154_)
  );
  INV_X1 _43566_ (
    .A(_09154_),
    .ZN(_09155_)
  );
  AND2_X1 _43567_ (
    .A1(_00007_[0]),
    .A2(_09155_),
    .ZN(_09156_)
  );
  INV_X1 _43568_ (
    .A(_09156_),
    .ZN(_09157_)
  );
  AND2_X1 _43569_ (
    .A1(_09149_),
    .A2(_09157_),
    .ZN(_09158_)
  );
  AND2_X1 _43570_ (
    .A1(\cpuregs[1] [24]),
    .A2(_22077_),
    .ZN(_09159_)
  );
  INV_X1 _43571_ (
    .A(_09159_),
    .ZN(_09160_)
  );
  AND2_X1 _43572_ (
    .A1(\cpuregs[5] [24]),
    .A2(_00007_[2]),
    .ZN(_09161_)
  );
  INV_X1 _43573_ (
    .A(_09161_),
    .ZN(_09162_)
  );
  AND2_X1 _43574_ (
    .A1(_09160_),
    .A2(_09162_),
    .ZN(_09163_)
  );
  INV_X1 _43575_ (
    .A(_09163_),
    .ZN(_09164_)
  );
  AND2_X1 _43576_ (
    .A1(_00007_[0]),
    .A2(_09164_),
    .ZN(_09165_)
  );
  INV_X1 _43577_ (
    .A(_09165_),
    .ZN(_09166_)
  );
  AND2_X1 _43578_ (
    .A1(\cpuregs[4] [24]),
    .A2(_00007_[2]),
    .ZN(_09167_)
  );
  INV_X1 _43579_ (
    .A(_09167_),
    .ZN(_09168_)
  );
  AND2_X1 _43580_ (
    .A1(\cpuregs[0] [24]),
    .A2(_22077_),
    .ZN(_09169_)
  );
  INV_X1 _43581_ (
    .A(_09169_),
    .ZN(_09170_)
  );
  AND2_X1 _43582_ (
    .A1(_09168_),
    .A2(_09170_),
    .ZN(_09171_)
  );
  INV_X1 _43583_ (
    .A(_09171_),
    .ZN(_09172_)
  );
  AND2_X1 _43584_ (
    .A1(_22152_),
    .A2(_09172_),
    .ZN(_09173_)
  );
  INV_X1 _43585_ (
    .A(_09173_),
    .ZN(_09174_)
  );
  AND2_X1 _43586_ (
    .A1(_09166_),
    .A2(_09174_),
    .ZN(_09175_)
  );
  AND2_X1 _43587_ (
    .A1(_00007_[1]),
    .A2(_09158_),
    .ZN(_09176_)
  );
  INV_X1 _43588_ (
    .A(_09176_),
    .ZN(_09177_)
  );
  AND2_X1 _43589_ (
    .A1(_22078_),
    .A2(_09175_),
    .ZN(_09178_)
  );
  INV_X1 _43590_ (
    .A(_09178_),
    .ZN(_09179_)
  );
  AND2_X1 _43591_ (
    .A1(_09177_),
    .A2(_09179_),
    .ZN(_09180_)
  );
  AND2_X1 _43592_ (
    .A1(_00007_[1]),
    .A2(_09142_),
    .ZN(_09181_)
  );
  INV_X1 _43593_ (
    .A(_09181_),
    .ZN(_09182_)
  );
  AND2_X1 _43594_ (
    .A1(_22078_),
    .A2(_09127_),
    .ZN(_09183_)
  );
  INV_X1 _43595_ (
    .A(_09183_),
    .ZN(_09184_)
  );
  AND2_X1 _43596_ (
    .A1(_22109_),
    .A2(_09184_),
    .ZN(_09185_)
  );
  AND2_X1 _43597_ (
    .A1(_09182_),
    .A2(_09185_),
    .ZN(_09186_)
  );
  INV_X1 _43598_ (
    .A(_09186_),
    .ZN(_09187_)
  );
  AND2_X1 _43599_ (
    .A1(_00007_[3]),
    .A2(_09078_),
    .ZN(_09188_)
  );
  INV_X1 _43600_ (
    .A(_09188_),
    .ZN(_09189_)
  );
  AND2_X1 _43601_ (
    .A1(_00007_[4]),
    .A2(_09189_),
    .ZN(_09190_)
  );
  AND2_X1 _43602_ (
    .A1(_09187_),
    .A2(_09190_),
    .ZN(_09191_)
  );
  INV_X1 _43603_ (
    .A(_09191_),
    .ZN(_09192_)
  );
  AND2_X1 _43604_ (
    .A1(_22109_),
    .A2(_09180_),
    .ZN(_09193_)
  );
  INV_X1 _43605_ (
    .A(_09193_),
    .ZN(_09194_)
  );
  AND2_X1 _43606_ (
    .A1(_00007_[1]),
    .A2(_09095_),
    .ZN(_09195_)
  );
  INV_X1 _43607_ (
    .A(_09195_),
    .ZN(_09196_)
  );
  AND2_X1 _43608_ (
    .A1(_22078_),
    .A2(_09112_),
    .ZN(_09197_)
  );
  INV_X1 _43609_ (
    .A(_09197_),
    .ZN(_09198_)
  );
  AND2_X1 _43610_ (
    .A1(_00007_[3]),
    .A2(_09198_),
    .ZN(_09199_)
  );
  AND2_X1 _43611_ (
    .A1(_09196_),
    .A2(_09199_),
    .ZN(_09200_)
  );
  INV_X1 _43612_ (
    .A(_09200_),
    .ZN(_09201_)
  );
  AND2_X1 _43613_ (
    .A1(_09194_),
    .A2(_09201_),
    .ZN(_09202_)
  );
  AND2_X1 _43614_ (
    .A1(_22144_),
    .A2(_09202_),
    .ZN(_09203_)
  );
  INV_X1 _43615_ (
    .A(_09203_),
    .ZN(_09204_)
  );
  AND2_X1 _43616_ (
    .A1(_09192_),
    .A2(_09204_),
    .ZN(_09205_)
  );
  AND2_X1 _43617_ (
    .A1(_05842_),
    .A2(_09205_),
    .ZN(_09206_)
  );
  INV_X1 _43618_ (
    .A(_09206_),
    .ZN(_09207_)
  );
  AND2_X1 _43619_ (
    .A1(_21224_),
    .A2(_04963_),
    .ZN(_09208_)
  );
  INV_X1 _43620_ (
    .A(_09208_),
    .ZN(_09209_)
  );
  AND2_X1 _43621_ (
    .A1(_04962_),
    .A2(_09207_),
    .ZN(_09210_)
  );
  AND2_X1 _43622_ (
    .A1(_09042_),
    .A2(_09210_),
    .ZN(_09211_)
  );
  INV_X1 _43623_ (
    .A(_09211_),
    .ZN(_09212_)
  );
  AND2_X1 _43624_ (
    .A1(_09209_),
    .A2(_09212_),
    .ZN(_00305_)
  );
  AND2_X1 _43625_ (
    .A1(decoded_imm[25]),
    .A2(_04966_),
    .ZN(_09213_)
  );
  INV_X1 _43626_ (
    .A(_09213_),
    .ZN(_09214_)
  );
  AND2_X1 _43627_ (
    .A1(_21610_),
    .A2(_22077_),
    .ZN(_09215_)
  );
  INV_X1 _43628_ (
    .A(_09215_),
    .ZN(_09216_)
  );
  AND2_X1 _43629_ (
    .A1(_21430_),
    .A2(_00007_[2]),
    .ZN(_09217_)
  );
  INV_X1 _43630_ (
    .A(_09217_),
    .ZN(_09218_)
  );
  AND2_X1 _43631_ (
    .A1(_21389_),
    .A2(_00007_[2]),
    .ZN(_09219_)
  );
  INV_X1 _43632_ (
    .A(_09219_),
    .ZN(_09220_)
  );
  AND2_X1 _43633_ (
    .A1(_21635_),
    .A2(_22077_),
    .ZN(_09221_)
  );
  INV_X1 _43634_ (
    .A(_09221_),
    .ZN(_09222_)
  );
  AND2_X1 _43635_ (
    .A1(\cpuregs[11] [25]),
    .A2(_22077_),
    .ZN(_09223_)
  );
  INV_X1 _43636_ (
    .A(_09223_),
    .ZN(_09224_)
  );
  AND2_X1 _43637_ (
    .A1(\cpuregs[15] [25]),
    .A2(_00007_[2]),
    .ZN(_09225_)
  );
  INV_X1 _43638_ (
    .A(_09225_),
    .ZN(_09226_)
  );
  AND2_X1 _43639_ (
    .A1(_09224_),
    .A2(_09226_),
    .ZN(_09227_)
  );
  INV_X1 _43640_ (
    .A(_09227_),
    .ZN(_09228_)
  );
  AND2_X1 _43641_ (
    .A1(_00007_[0]),
    .A2(_09228_),
    .ZN(_09229_)
  );
  INV_X1 _43642_ (
    .A(_09229_),
    .ZN(_09230_)
  );
  AND2_X1 _43643_ (
    .A1(\cpuregs[14] [25]),
    .A2(_00007_[2]),
    .ZN(_09231_)
  );
  INV_X1 _43644_ (
    .A(_09231_),
    .ZN(_09232_)
  );
  AND2_X1 _43645_ (
    .A1(\cpuregs[10] [25]),
    .A2(_22077_),
    .ZN(_09233_)
  );
  INV_X1 _43646_ (
    .A(_09233_),
    .ZN(_09234_)
  );
  AND2_X1 _43647_ (
    .A1(_09232_),
    .A2(_09234_),
    .ZN(_09235_)
  );
  INV_X1 _43648_ (
    .A(_09235_),
    .ZN(_09236_)
  );
  AND2_X1 _43649_ (
    .A1(_22152_),
    .A2(_09236_),
    .ZN(_09237_)
  );
  INV_X1 _43650_ (
    .A(_09237_),
    .ZN(_09238_)
  );
  AND2_X1 _43651_ (
    .A1(_09230_),
    .A2(_09238_),
    .ZN(_09239_)
  );
  AND2_X1 _43652_ (
    .A1(_21561_),
    .A2(_22077_),
    .ZN(_09240_)
  );
  INV_X1 _43653_ (
    .A(_09240_),
    .ZN(_09241_)
  );
  AND2_X1 _43654_ (
    .A1(_21827_),
    .A2(_00007_[2]),
    .ZN(_09242_)
  );
  INV_X1 _43655_ (
    .A(_09242_),
    .ZN(_09243_)
  );
  AND2_X1 _43656_ (
    .A1(_22152_),
    .A2(_09243_),
    .ZN(_09244_)
  );
  AND2_X1 _43657_ (
    .A1(_09241_),
    .A2(_09244_),
    .ZN(_09245_)
  );
  INV_X1 _43658_ (
    .A(_09245_),
    .ZN(_09246_)
  );
  AND2_X1 _43659_ (
    .A1(_21798_),
    .A2(_00007_[2]),
    .ZN(_09247_)
  );
  INV_X1 _43660_ (
    .A(_09247_),
    .ZN(_09248_)
  );
  AND2_X1 _43661_ (
    .A1(_21506_),
    .A2(_22077_),
    .ZN(_09249_)
  );
  INV_X1 _43662_ (
    .A(_09249_),
    .ZN(_09250_)
  );
  AND2_X1 _43663_ (
    .A1(_00007_[0]),
    .A2(_09250_),
    .ZN(_09251_)
  );
  AND2_X1 _43664_ (
    .A1(_09248_),
    .A2(_09251_),
    .ZN(_09252_)
  );
  INV_X1 _43665_ (
    .A(_09252_),
    .ZN(_09253_)
  );
  AND2_X1 _43666_ (
    .A1(_09246_),
    .A2(_09253_),
    .ZN(_09254_)
  );
  AND2_X1 _43667_ (
    .A1(_21454_),
    .A2(_22077_),
    .ZN(_09255_)
  );
  INV_X1 _43668_ (
    .A(_09255_),
    .ZN(_09256_)
  );
  AND2_X1 _43669_ (
    .A1(_21665_),
    .A2(_00007_[2]),
    .ZN(_09257_)
  );
  INV_X1 _43670_ (
    .A(_09257_),
    .ZN(_09258_)
  );
  AND2_X1 _43671_ (
    .A1(_09256_),
    .A2(_09258_),
    .ZN(_09259_)
  );
  AND2_X1 _43672_ (
    .A1(_21476_),
    .A2(_22077_),
    .ZN(_09260_)
  );
  INV_X1 _43673_ (
    .A(_09260_),
    .ZN(_09261_)
  );
  AND2_X1 _43674_ (
    .A1(_21775_),
    .A2(_00007_[2]),
    .ZN(_09262_)
  );
  INV_X1 _43675_ (
    .A(_09262_),
    .ZN(_09263_)
  );
  AND2_X1 _43676_ (
    .A1(\cpuregs[9] [25]),
    .A2(_22077_),
    .ZN(_09264_)
  );
  INV_X1 _43677_ (
    .A(_09264_),
    .ZN(_09265_)
  );
  AND2_X1 _43678_ (
    .A1(\cpuregs[13] [25]),
    .A2(_00007_[2]),
    .ZN(_09266_)
  );
  INV_X1 _43679_ (
    .A(_09266_),
    .ZN(_09267_)
  );
  AND2_X1 _43680_ (
    .A1(_09265_),
    .A2(_09267_),
    .ZN(_09268_)
  );
  INV_X1 _43681_ (
    .A(_09268_),
    .ZN(_09269_)
  );
  AND2_X1 _43682_ (
    .A1(_00007_[0]),
    .A2(_09269_),
    .ZN(_09270_)
  );
  INV_X1 _43683_ (
    .A(_09270_),
    .ZN(_09271_)
  );
  AND2_X1 _43684_ (
    .A1(\cpuregs[12] [25]),
    .A2(_00007_[2]),
    .ZN(_09272_)
  );
  INV_X1 _43685_ (
    .A(_09272_),
    .ZN(_09273_)
  );
  AND2_X1 _43686_ (
    .A1(\cpuregs[8] [25]),
    .A2(_22077_),
    .ZN(_09274_)
  );
  INV_X1 _43687_ (
    .A(_09274_),
    .ZN(_09275_)
  );
  AND2_X1 _43688_ (
    .A1(_09273_),
    .A2(_09275_),
    .ZN(_09276_)
  );
  INV_X1 _43689_ (
    .A(_09276_),
    .ZN(_09277_)
  );
  AND2_X1 _43690_ (
    .A1(_22152_),
    .A2(_09277_),
    .ZN(_09278_)
  );
  INV_X1 _43691_ (
    .A(_09278_),
    .ZN(_09279_)
  );
  AND2_X1 _43692_ (
    .A1(_09271_),
    .A2(_09279_),
    .ZN(_09280_)
  );
  AND2_X1 _43693_ (
    .A1(_21688_),
    .A2(_00007_[2]),
    .ZN(_09281_)
  );
  INV_X1 _43694_ (
    .A(_09281_),
    .ZN(_09282_)
  );
  AND2_X1 _43695_ (
    .A1(_21972_),
    .A2(_22077_),
    .ZN(_09283_)
  );
  INV_X1 _43696_ (
    .A(_09283_),
    .ZN(_09284_)
  );
  AND2_X1 _43697_ (
    .A1(_09282_),
    .A2(_09284_),
    .ZN(_09285_)
  );
  AND2_X1 _43698_ (
    .A1(_22152_),
    .A2(_09285_),
    .ZN(_09286_)
  );
  INV_X1 _43699_ (
    .A(_09286_),
    .ZN(_09287_)
  );
  AND2_X1 _43700_ (
    .A1(_21531_),
    .A2(_22077_),
    .ZN(_09288_)
  );
  INV_X1 _43701_ (
    .A(_09288_),
    .ZN(_09289_)
  );
  AND2_X1 _43702_ (
    .A1(_21751_),
    .A2(_00007_[2]),
    .ZN(_09290_)
  );
  INV_X1 _43703_ (
    .A(_09290_),
    .ZN(_09291_)
  );
  AND2_X1 _43704_ (
    .A1(_00007_[0]),
    .A2(_09291_),
    .ZN(_09292_)
  );
  AND2_X1 _43705_ (
    .A1(_09289_),
    .A2(_09292_),
    .ZN(_09293_)
  );
  INV_X1 _43706_ (
    .A(_09293_),
    .ZN(_09294_)
  );
  AND2_X1 _43707_ (
    .A1(_09287_),
    .A2(_09294_),
    .ZN(_09295_)
  );
  AND2_X1 _43708_ (
    .A1(_22152_),
    .A2(_09218_),
    .ZN(_09296_)
  );
  AND2_X1 _43709_ (
    .A1(_09216_),
    .A2(_09296_),
    .ZN(_09297_)
  );
  INV_X1 _43710_ (
    .A(_09297_),
    .ZN(_09298_)
  );
  AND2_X1 _43711_ (
    .A1(_00007_[0]),
    .A2(_09220_),
    .ZN(_09299_)
  );
  AND2_X1 _43712_ (
    .A1(_09222_),
    .A2(_09299_),
    .ZN(_09300_)
  );
  INV_X1 _43713_ (
    .A(_09300_),
    .ZN(_09301_)
  );
  AND2_X1 _43714_ (
    .A1(_09298_),
    .A2(_09301_),
    .ZN(_09302_)
  );
  AND2_X1 _43715_ (
    .A1(_00007_[1]),
    .A2(_09302_),
    .ZN(_09303_)
  );
  INV_X1 _43716_ (
    .A(_09303_),
    .ZN(_09304_)
  );
  AND2_X1 _43717_ (
    .A1(_00007_[0]),
    .A2(_09263_),
    .ZN(_09305_)
  );
  AND2_X1 _43718_ (
    .A1(_09261_),
    .A2(_09305_),
    .ZN(_09306_)
  );
  INV_X1 _43719_ (
    .A(_09306_),
    .ZN(_09307_)
  );
  AND2_X1 _43720_ (
    .A1(_22152_),
    .A2(_09259_),
    .ZN(_09308_)
  );
  INV_X1 _43721_ (
    .A(_09308_),
    .ZN(_09309_)
  );
  AND2_X1 _43722_ (
    .A1(_09307_),
    .A2(_09309_),
    .ZN(_09310_)
  );
  AND2_X1 _43723_ (
    .A1(_22078_),
    .A2(_09310_),
    .ZN(_09311_)
  );
  INV_X1 _43724_ (
    .A(_09311_),
    .ZN(_09312_)
  );
  AND2_X1 _43725_ (
    .A1(_22109_),
    .A2(_09312_),
    .ZN(_09313_)
  );
  AND2_X1 _43726_ (
    .A1(_09304_),
    .A2(_09313_),
    .ZN(_09314_)
  );
  INV_X1 _43727_ (
    .A(_09314_),
    .ZN(_09315_)
  );
  AND2_X1 _43728_ (
    .A1(_21933_),
    .A2(_22077_),
    .ZN(_09316_)
  );
  INV_X1 _43729_ (
    .A(_09316_),
    .ZN(_09317_)
  );
  AND2_X1 _43730_ (
    .A1(_21949_),
    .A2(_00007_[2]),
    .ZN(_09318_)
  );
  INV_X1 _43731_ (
    .A(_09318_),
    .ZN(_09319_)
  );
  AND2_X1 _43732_ (
    .A1(_00007_[0]),
    .A2(_09319_),
    .ZN(_09320_)
  );
  AND2_X1 _43733_ (
    .A1(_09317_),
    .A2(_09320_),
    .ZN(_09321_)
  );
  INV_X1 _43734_ (
    .A(_09321_),
    .ZN(_09322_)
  );
  AND2_X1 _43735_ (
    .A1(_21883_),
    .A2(_22077_),
    .ZN(_09323_)
  );
  INV_X1 _43736_ (
    .A(_09323_),
    .ZN(_09324_)
  );
  AND2_X1 _43737_ (
    .A1(_21861_),
    .A2(_00007_[2]),
    .ZN(_09325_)
  );
  INV_X1 _43738_ (
    .A(_09325_),
    .ZN(_09326_)
  );
  AND2_X1 _43739_ (
    .A1(_09324_),
    .A2(_09326_),
    .ZN(_09327_)
  );
  AND2_X1 _43740_ (
    .A1(_22152_),
    .A2(_09327_),
    .ZN(_09328_)
  );
  INV_X1 _43741_ (
    .A(_09328_),
    .ZN(_09329_)
  );
  AND2_X1 _43742_ (
    .A1(_09322_),
    .A2(_09329_),
    .ZN(_09330_)
  );
  AND2_X1 _43743_ (
    .A1(_00007_[1]),
    .A2(_09330_),
    .ZN(_09331_)
  );
  INV_X1 _43744_ (
    .A(_09331_),
    .ZN(_09332_)
  );
  AND2_X1 _43745_ (
    .A1(_21845_),
    .A2(_22077_),
    .ZN(_09333_)
  );
  INV_X1 _43746_ (
    .A(_09333_),
    .ZN(_09334_)
  );
  AND2_X1 _43747_ (
    .A1(_21901_),
    .A2(_00007_[2]),
    .ZN(_09335_)
  );
  INV_X1 _43748_ (
    .A(_09335_),
    .ZN(_09336_)
  );
  AND2_X1 _43749_ (
    .A1(_00007_[0]),
    .A2(_09336_),
    .ZN(_09337_)
  );
  AND2_X1 _43750_ (
    .A1(_09334_),
    .A2(_09337_),
    .ZN(_09338_)
  );
  INV_X1 _43751_ (
    .A(_09338_),
    .ZN(_09339_)
  );
  AND2_X1 _43752_ (
    .A1(_21579_),
    .A2(_22077_),
    .ZN(_09340_)
  );
  INV_X1 _43753_ (
    .A(_09340_),
    .ZN(_09341_)
  );
  AND2_X1 _43754_ (
    .A1(_21917_),
    .A2(_00007_[2]),
    .ZN(_09342_)
  );
  INV_X1 _43755_ (
    .A(_09342_),
    .ZN(_09343_)
  );
  AND2_X1 _43756_ (
    .A1(_09341_),
    .A2(_09343_),
    .ZN(_09344_)
  );
  AND2_X1 _43757_ (
    .A1(_22152_),
    .A2(_09344_),
    .ZN(_09345_)
  );
  INV_X1 _43758_ (
    .A(_09345_),
    .ZN(_09346_)
  );
  AND2_X1 _43759_ (
    .A1(_09339_),
    .A2(_09346_),
    .ZN(_09347_)
  );
  AND2_X1 _43760_ (
    .A1(_22078_),
    .A2(_09347_),
    .ZN(_09348_)
  );
  INV_X1 _43761_ (
    .A(_09348_),
    .ZN(_09349_)
  );
  AND2_X1 _43762_ (
    .A1(_00007_[3]),
    .A2(_09349_),
    .ZN(_09350_)
  );
  AND2_X1 _43763_ (
    .A1(_09332_),
    .A2(_09350_),
    .ZN(_09351_)
  );
  INV_X1 _43764_ (
    .A(_09351_),
    .ZN(_09352_)
  );
  AND2_X1 _43765_ (
    .A1(_00007_[4]),
    .A2(_09352_),
    .ZN(_09353_)
  );
  AND2_X1 _43766_ (
    .A1(_09315_),
    .A2(_09353_),
    .ZN(_09354_)
  );
  INV_X1 _43767_ (
    .A(_09354_),
    .ZN(_09355_)
  );
  AND2_X1 _43768_ (
    .A1(_00007_[1]),
    .A2(_09254_),
    .ZN(_09356_)
  );
  INV_X1 _43769_ (
    .A(_09356_),
    .ZN(_09357_)
  );
  AND2_X1 _43770_ (
    .A1(_22078_),
    .A2(_09295_),
    .ZN(_09358_)
  );
  INV_X1 _43771_ (
    .A(_09358_),
    .ZN(_09359_)
  );
  AND2_X1 _43772_ (
    .A1(_22109_),
    .A2(_09359_),
    .ZN(_09360_)
  );
  AND2_X1 _43773_ (
    .A1(_09357_),
    .A2(_09360_),
    .ZN(_09361_)
  );
  INV_X1 _43774_ (
    .A(_09361_),
    .ZN(_09362_)
  );
  AND2_X1 _43775_ (
    .A1(_00007_[1]),
    .A2(_09239_),
    .ZN(_09363_)
  );
  INV_X1 _43776_ (
    .A(_09363_),
    .ZN(_09364_)
  );
  AND2_X1 _43777_ (
    .A1(_22078_),
    .A2(_09280_),
    .ZN(_09365_)
  );
  INV_X1 _43778_ (
    .A(_09365_),
    .ZN(_09366_)
  );
  AND2_X1 _43779_ (
    .A1(_00007_[3]),
    .A2(_09366_),
    .ZN(_09367_)
  );
  AND2_X1 _43780_ (
    .A1(_09364_),
    .A2(_09367_),
    .ZN(_09368_)
  );
  INV_X1 _43781_ (
    .A(_09368_),
    .ZN(_09369_)
  );
  AND2_X1 _43782_ (
    .A1(_09362_),
    .A2(_09369_),
    .ZN(_09370_)
  );
  AND2_X1 _43783_ (
    .A1(_22144_),
    .A2(_09370_),
    .ZN(_09371_)
  );
  INV_X1 _43784_ (
    .A(_09371_),
    .ZN(_09372_)
  );
  AND2_X1 _43785_ (
    .A1(_09355_),
    .A2(_09372_),
    .ZN(_09373_)
  );
  AND2_X1 _43786_ (
    .A1(_05842_),
    .A2(_09373_),
    .ZN(_09374_)
  );
  INV_X1 _43787_ (
    .A(_09374_),
    .ZN(_09375_)
  );
  AND2_X1 _43788_ (
    .A1(_21225_),
    .A2(_04963_),
    .ZN(_09376_)
  );
  INV_X1 _43789_ (
    .A(_09376_),
    .ZN(_09377_)
  );
  AND2_X1 _43790_ (
    .A1(_04962_),
    .A2(_09375_),
    .ZN(_09378_)
  );
  AND2_X1 _43791_ (
    .A1(_09214_),
    .A2(_09378_),
    .ZN(_09379_)
  );
  INV_X1 _43792_ (
    .A(_09379_),
    .ZN(_09380_)
  );
  AND2_X1 _43793_ (
    .A1(_09377_),
    .A2(_09380_),
    .ZN(_00306_)
  );
  AND2_X1 _43794_ (
    .A1(_21611_),
    .A2(_22077_),
    .ZN(_09381_)
  );
  INV_X1 _43795_ (
    .A(_09381_),
    .ZN(_09382_)
  );
  AND2_X1 _43796_ (
    .A1(_21431_),
    .A2(_00007_[2]),
    .ZN(_09383_)
  );
  INV_X1 _43797_ (
    .A(_09383_),
    .ZN(_09384_)
  );
  AND2_X1 _43798_ (
    .A1(_21390_),
    .A2(_00007_[2]),
    .ZN(_09385_)
  );
  INV_X1 _43799_ (
    .A(_09385_),
    .ZN(_09386_)
  );
  AND2_X1 _43800_ (
    .A1(_21636_),
    .A2(_22077_),
    .ZN(_09387_)
  );
  INV_X1 _43801_ (
    .A(_09387_),
    .ZN(_09388_)
  );
  AND2_X1 _43802_ (
    .A1(\cpuregs[11] [26]),
    .A2(_22077_),
    .ZN(_09389_)
  );
  INV_X1 _43803_ (
    .A(_09389_),
    .ZN(_09390_)
  );
  AND2_X1 _43804_ (
    .A1(\cpuregs[15] [26]),
    .A2(_00007_[2]),
    .ZN(_09391_)
  );
  INV_X1 _43805_ (
    .A(_09391_),
    .ZN(_09392_)
  );
  AND2_X1 _43806_ (
    .A1(_09390_),
    .A2(_09392_),
    .ZN(_09393_)
  );
  INV_X1 _43807_ (
    .A(_09393_),
    .ZN(_09394_)
  );
  AND2_X1 _43808_ (
    .A1(_00007_[0]),
    .A2(_09394_),
    .ZN(_09395_)
  );
  INV_X1 _43809_ (
    .A(_09395_),
    .ZN(_09396_)
  );
  AND2_X1 _43810_ (
    .A1(\cpuregs[14] [26]),
    .A2(_00007_[2]),
    .ZN(_09397_)
  );
  INV_X1 _43811_ (
    .A(_09397_),
    .ZN(_09398_)
  );
  AND2_X1 _43812_ (
    .A1(\cpuregs[10] [26]),
    .A2(_22077_),
    .ZN(_09399_)
  );
  INV_X1 _43813_ (
    .A(_09399_),
    .ZN(_09400_)
  );
  AND2_X1 _43814_ (
    .A1(_09398_),
    .A2(_09400_),
    .ZN(_09401_)
  );
  INV_X1 _43815_ (
    .A(_09401_),
    .ZN(_09402_)
  );
  AND2_X1 _43816_ (
    .A1(_22152_),
    .A2(_09402_),
    .ZN(_09403_)
  );
  INV_X1 _43817_ (
    .A(_09403_),
    .ZN(_09404_)
  );
  AND2_X1 _43818_ (
    .A1(_09396_),
    .A2(_09404_),
    .ZN(_09405_)
  );
  AND2_X1 _43819_ (
    .A1(_21562_),
    .A2(_22077_),
    .ZN(_09406_)
  );
  INV_X1 _43820_ (
    .A(_09406_),
    .ZN(_09407_)
  );
  AND2_X1 _43821_ (
    .A1(_21828_),
    .A2(_00007_[2]),
    .ZN(_09408_)
  );
  INV_X1 _43822_ (
    .A(_09408_),
    .ZN(_09409_)
  );
  AND2_X1 _43823_ (
    .A1(_22152_),
    .A2(_09409_),
    .ZN(_09410_)
  );
  AND2_X1 _43824_ (
    .A1(_09407_),
    .A2(_09410_),
    .ZN(_09411_)
  );
  INV_X1 _43825_ (
    .A(_09411_),
    .ZN(_09412_)
  );
  AND2_X1 _43826_ (
    .A1(_21799_),
    .A2(_00007_[2]),
    .ZN(_09413_)
  );
  INV_X1 _43827_ (
    .A(_09413_),
    .ZN(_09414_)
  );
  AND2_X1 _43828_ (
    .A1(_21507_),
    .A2(_22077_),
    .ZN(_09415_)
  );
  INV_X1 _43829_ (
    .A(_09415_),
    .ZN(_09416_)
  );
  AND2_X1 _43830_ (
    .A1(_00007_[0]),
    .A2(_09416_),
    .ZN(_09417_)
  );
  AND2_X1 _43831_ (
    .A1(_09414_),
    .A2(_09417_),
    .ZN(_09418_)
  );
  INV_X1 _43832_ (
    .A(_09418_),
    .ZN(_09419_)
  );
  AND2_X1 _43833_ (
    .A1(_09412_),
    .A2(_09419_),
    .ZN(_09420_)
  );
  AND2_X1 _43834_ (
    .A1(_21455_),
    .A2(_22077_),
    .ZN(_09421_)
  );
  INV_X1 _43835_ (
    .A(_09421_),
    .ZN(_09422_)
  );
  AND2_X1 _43836_ (
    .A1(_21666_),
    .A2(_00007_[2]),
    .ZN(_09423_)
  );
  INV_X1 _43837_ (
    .A(_09423_),
    .ZN(_09424_)
  );
  AND2_X1 _43838_ (
    .A1(_09422_),
    .A2(_09424_),
    .ZN(_09425_)
  );
  AND2_X1 _43839_ (
    .A1(_21477_),
    .A2(_22077_),
    .ZN(_09426_)
  );
  INV_X1 _43840_ (
    .A(_09426_),
    .ZN(_09427_)
  );
  AND2_X1 _43841_ (
    .A1(_21776_),
    .A2(_00007_[2]),
    .ZN(_09428_)
  );
  INV_X1 _43842_ (
    .A(_09428_),
    .ZN(_09429_)
  );
  AND2_X1 _43843_ (
    .A1(\cpuregs[9] [26]),
    .A2(_22077_),
    .ZN(_09430_)
  );
  INV_X1 _43844_ (
    .A(_09430_),
    .ZN(_09431_)
  );
  AND2_X1 _43845_ (
    .A1(\cpuregs[13] [26]),
    .A2(_00007_[2]),
    .ZN(_09432_)
  );
  INV_X1 _43846_ (
    .A(_09432_),
    .ZN(_09433_)
  );
  AND2_X1 _43847_ (
    .A1(_09431_),
    .A2(_09433_),
    .ZN(_09434_)
  );
  INV_X1 _43848_ (
    .A(_09434_),
    .ZN(_09435_)
  );
  AND2_X1 _43849_ (
    .A1(_00007_[0]),
    .A2(_09435_),
    .ZN(_09436_)
  );
  INV_X1 _43850_ (
    .A(_09436_),
    .ZN(_09437_)
  );
  AND2_X1 _43851_ (
    .A1(\cpuregs[12] [26]),
    .A2(_00007_[2]),
    .ZN(_09438_)
  );
  INV_X1 _43852_ (
    .A(_09438_),
    .ZN(_09439_)
  );
  AND2_X1 _43853_ (
    .A1(\cpuregs[8] [26]),
    .A2(_22077_),
    .ZN(_09440_)
  );
  INV_X1 _43854_ (
    .A(_09440_),
    .ZN(_09441_)
  );
  AND2_X1 _43855_ (
    .A1(_09439_),
    .A2(_09441_),
    .ZN(_09442_)
  );
  INV_X1 _43856_ (
    .A(_09442_),
    .ZN(_09443_)
  );
  AND2_X1 _43857_ (
    .A1(_22152_),
    .A2(_09443_),
    .ZN(_09444_)
  );
  INV_X1 _43858_ (
    .A(_09444_),
    .ZN(_09445_)
  );
  AND2_X1 _43859_ (
    .A1(_09437_),
    .A2(_09445_),
    .ZN(_09446_)
  );
  AND2_X1 _43860_ (
    .A1(_21689_),
    .A2(_00007_[2]),
    .ZN(_09447_)
  );
  INV_X1 _43861_ (
    .A(_09447_),
    .ZN(_09448_)
  );
  AND2_X1 _43862_ (
    .A1(_21973_),
    .A2(_22077_),
    .ZN(_09449_)
  );
  INV_X1 _43863_ (
    .A(_09449_),
    .ZN(_09450_)
  );
  AND2_X1 _43864_ (
    .A1(_09448_),
    .A2(_09450_),
    .ZN(_09451_)
  );
  AND2_X1 _43865_ (
    .A1(_22152_),
    .A2(_09451_),
    .ZN(_09452_)
  );
  INV_X1 _43866_ (
    .A(_09452_),
    .ZN(_09453_)
  );
  AND2_X1 _43867_ (
    .A1(_21532_),
    .A2(_22077_),
    .ZN(_09454_)
  );
  INV_X1 _43868_ (
    .A(_09454_),
    .ZN(_09455_)
  );
  AND2_X1 _43869_ (
    .A1(_21752_),
    .A2(_00007_[2]),
    .ZN(_09456_)
  );
  INV_X1 _43870_ (
    .A(_09456_),
    .ZN(_09457_)
  );
  AND2_X1 _43871_ (
    .A1(_00007_[0]),
    .A2(_09457_),
    .ZN(_09458_)
  );
  AND2_X1 _43872_ (
    .A1(_09455_),
    .A2(_09458_),
    .ZN(_09459_)
  );
  INV_X1 _43873_ (
    .A(_09459_),
    .ZN(_09460_)
  );
  AND2_X1 _43874_ (
    .A1(_09453_),
    .A2(_09460_),
    .ZN(_09461_)
  );
  AND2_X1 _43875_ (
    .A1(_22152_),
    .A2(_09384_),
    .ZN(_09462_)
  );
  AND2_X1 _43876_ (
    .A1(_09382_),
    .A2(_09462_),
    .ZN(_09463_)
  );
  INV_X1 _43877_ (
    .A(_09463_),
    .ZN(_09464_)
  );
  AND2_X1 _43878_ (
    .A1(_00007_[0]),
    .A2(_09386_),
    .ZN(_09465_)
  );
  AND2_X1 _43879_ (
    .A1(_09388_),
    .A2(_09465_),
    .ZN(_09466_)
  );
  INV_X1 _43880_ (
    .A(_09466_),
    .ZN(_09467_)
  );
  AND2_X1 _43881_ (
    .A1(_09464_),
    .A2(_09467_),
    .ZN(_09468_)
  );
  AND2_X1 _43882_ (
    .A1(_00007_[1]),
    .A2(_09468_),
    .ZN(_09469_)
  );
  INV_X1 _43883_ (
    .A(_09469_),
    .ZN(_09470_)
  );
  AND2_X1 _43884_ (
    .A1(_00007_[0]),
    .A2(_09429_),
    .ZN(_09471_)
  );
  AND2_X1 _43885_ (
    .A1(_09427_),
    .A2(_09471_),
    .ZN(_09472_)
  );
  INV_X1 _43886_ (
    .A(_09472_),
    .ZN(_09473_)
  );
  AND2_X1 _43887_ (
    .A1(_22152_),
    .A2(_09425_),
    .ZN(_09474_)
  );
  INV_X1 _43888_ (
    .A(_09474_),
    .ZN(_09475_)
  );
  AND2_X1 _43889_ (
    .A1(_09473_),
    .A2(_09475_),
    .ZN(_09476_)
  );
  AND2_X1 _43890_ (
    .A1(_22078_),
    .A2(_09476_),
    .ZN(_09477_)
  );
  INV_X1 _43891_ (
    .A(_09477_),
    .ZN(_09478_)
  );
  AND2_X1 _43892_ (
    .A1(_22109_),
    .A2(_09478_),
    .ZN(_09479_)
  );
  AND2_X1 _43893_ (
    .A1(_09470_),
    .A2(_09479_),
    .ZN(_09480_)
  );
  INV_X1 _43894_ (
    .A(_09480_),
    .ZN(_09481_)
  );
  AND2_X1 _43895_ (
    .A1(_21934_),
    .A2(_22077_),
    .ZN(_09482_)
  );
  INV_X1 _43896_ (
    .A(_09482_),
    .ZN(_09483_)
  );
  AND2_X1 _43897_ (
    .A1(_21950_),
    .A2(_00007_[2]),
    .ZN(_09484_)
  );
  INV_X1 _43898_ (
    .A(_09484_),
    .ZN(_09485_)
  );
  AND2_X1 _43899_ (
    .A1(_00007_[0]),
    .A2(_09485_),
    .ZN(_09486_)
  );
  AND2_X1 _43900_ (
    .A1(_09483_),
    .A2(_09486_),
    .ZN(_09487_)
  );
  INV_X1 _43901_ (
    .A(_09487_),
    .ZN(_09488_)
  );
  AND2_X1 _43902_ (
    .A1(_21884_),
    .A2(_22077_),
    .ZN(_09489_)
  );
  INV_X1 _43903_ (
    .A(_09489_),
    .ZN(_09490_)
  );
  AND2_X1 _43904_ (
    .A1(_21862_),
    .A2(_00007_[2]),
    .ZN(_09491_)
  );
  INV_X1 _43905_ (
    .A(_09491_),
    .ZN(_09492_)
  );
  AND2_X1 _43906_ (
    .A1(_09490_),
    .A2(_09492_),
    .ZN(_09493_)
  );
  AND2_X1 _43907_ (
    .A1(_22152_),
    .A2(_09493_),
    .ZN(_09494_)
  );
  INV_X1 _43908_ (
    .A(_09494_),
    .ZN(_09495_)
  );
  AND2_X1 _43909_ (
    .A1(_09488_),
    .A2(_09495_),
    .ZN(_09496_)
  );
  AND2_X1 _43910_ (
    .A1(_00007_[1]),
    .A2(_09496_),
    .ZN(_09497_)
  );
  INV_X1 _43911_ (
    .A(_09497_),
    .ZN(_09498_)
  );
  AND2_X1 _43912_ (
    .A1(_21846_),
    .A2(_22077_),
    .ZN(_09499_)
  );
  INV_X1 _43913_ (
    .A(_09499_),
    .ZN(_09500_)
  );
  AND2_X1 _43914_ (
    .A1(_21902_),
    .A2(_00007_[2]),
    .ZN(_09501_)
  );
  INV_X1 _43915_ (
    .A(_09501_),
    .ZN(_09502_)
  );
  AND2_X1 _43916_ (
    .A1(_00007_[0]),
    .A2(_09502_),
    .ZN(_09503_)
  );
  AND2_X1 _43917_ (
    .A1(_09500_),
    .A2(_09503_),
    .ZN(_09504_)
  );
  INV_X1 _43918_ (
    .A(_09504_),
    .ZN(_09505_)
  );
  AND2_X1 _43919_ (
    .A1(_21580_),
    .A2(_22077_),
    .ZN(_09506_)
  );
  INV_X1 _43920_ (
    .A(_09506_),
    .ZN(_09507_)
  );
  AND2_X1 _43921_ (
    .A1(_21918_),
    .A2(_00007_[2]),
    .ZN(_09508_)
  );
  INV_X1 _43922_ (
    .A(_09508_),
    .ZN(_09509_)
  );
  AND2_X1 _43923_ (
    .A1(_09507_),
    .A2(_09509_),
    .ZN(_09510_)
  );
  AND2_X1 _43924_ (
    .A1(_22152_),
    .A2(_09510_),
    .ZN(_09511_)
  );
  INV_X1 _43925_ (
    .A(_09511_),
    .ZN(_09512_)
  );
  AND2_X1 _43926_ (
    .A1(_09505_),
    .A2(_09512_),
    .ZN(_09513_)
  );
  AND2_X1 _43927_ (
    .A1(_22078_),
    .A2(_09513_),
    .ZN(_09514_)
  );
  INV_X1 _43928_ (
    .A(_09514_),
    .ZN(_09515_)
  );
  AND2_X1 _43929_ (
    .A1(_00007_[3]),
    .A2(_09515_),
    .ZN(_09516_)
  );
  AND2_X1 _43930_ (
    .A1(_09498_),
    .A2(_09516_),
    .ZN(_09517_)
  );
  INV_X1 _43931_ (
    .A(_09517_),
    .ZN(_09518_)
  );
  AND2_X1 _43932_ (
    .A1(_00007_[4]),
    .A2(_09518_),
    .ZN(_09519_)
  );
  AND2_X1 _43933_ (
    .A1(_09481_),
    .A2(_09519_),
    .ZN(_09520_)
  );
  INV_X1 _43934_ (
    .A(_09520_),
    .ZN(_09521_)
  );
  AND2_X1 _43935_ (
    .A1(_00007_[1]),
    .A2(_09420_),
    .ZN(_09522_)
  );
  INV_X1 _43936_ (
    .A(_09522_),
    .ZN(_09523_)
  );
  AND2_X1 _43937_ (
    .A1(_22078_),
    .A2(_09461_),
    .ZN(_09524_)
  );
  INV_X1 _43938_ (
    .A(_09524_),
    .ZN(_09525_)
  );
  AND2_X1 _43939_ (
    .A1(_22109_),
    .A2(_09525_),
    .ZN(_09526_)
  );
  AND2_X1 _43940_ (
    .A1(_09523_),
    .A2(_09526_),
    .ZN(_09527_)
  );
  INV_X1 _43941_ (
    .A(_09527_),
    .ZN(_09528_)
  );
  AND2_X1 _43942_ (
    .A1(_00007_[1]),
    .A2(_09405_),
    .ZN(_09529_)
  );
  INV_X1 _43943_ (
    .A(_09529_),
    .ZN(_09530_)
  );
  AND2_X1 _43944_ (
    .A1(_22078_),
    .A2(_09446_),
    .ZN(_09531_)
  );
  INV_X1 _43945_ (
    .A(_09531_),
    .ZN(_09532_)
  );
  AND2_X1 _43946_ (
    .A1(_00007_[3]),
    .A2(_09532_),
    .ZN(_09533_)
  );
  AND2_X1 _43947_ (
    .A1(_09530_),
    .A2(_09533_),
    .ZN(_09534_)
  );
  INV_X1 _43948_ (
    .A(_09534_),
    .ZN(_09535_)
  );
  AND2_X1 _43949_ (
    .A1(_09528_),
    .A2(_09535_),
    .ZN(_09536_)
  );
  AND2_X1 _43950_ (
    .A1(_22144_),
    .A2(_09536_),
    .ZN(_09537_)
  );
  INV_X1 _43951_ (
    .A(_09537_),
    .ZN(_09538_)
  );
  AND2_X1 _43952_ (
    .A1(_09521_),
    .A2(_09538_),
    .ZN(_09539_)
  );
  AND2_X1 _43953_ (
    .A1(_05842_),
    .A2(_09539_),
    .ZN(_09540_)
  );
  INV_X1 _43954_ (
    .A(_09540_),
    .ZN(_09541_)
  );
  AND2_X1 _43955_ (
    .A1(decoded_imm[26]),
    .A2(_04966_),
    .ZN(_09542_)
  );
  INV_X1 _43956_ (
    .A(_09542_),
    .ZN(_09543_)
  );
  AND2_X1 _43957_ (
    .A1(_21226_),
    .A2(_04963_),
    .ZN(_09544_)
  );
  INV_X1 _43958_ (
    .A(_09544_),
    .ZN(_09545_)
  );
  AND2_X1 _43959_ (
    .A1(_04962_),
    .A2(_09543_),
    .ZN(_09546_)
  );
  AND2_X1 _43960_ (
    .A1(_09541_),
    .A2(_09546_),
    .ZN(_09547_)
  );
  INV_X1 _43961_ (
    .A(_09547_),
    .ZN(_09548_)
  );
  AND2_X1 _43962_ (
    .A1(_09545_),
    .A2(_09548_),
    .ZN(_00307_)
  );
  AND2_X1 _43963_ (
    .A1(decoded_imm[27]),
    .A2(_04966_),
    .ZN(_09549_)
  );
  INV_X1 _43964_ (
    .A(_09549_),
    .ZN(_09550_)
  );
  AND2_X1 _43965_ (
    .A1(\cpuregs[19] [27]),
    .A2(_22077_),
    .ZN(_09551_)
  );
  INV_X1 _43966_ (
    .A(_09551_),
    .ZN(_09552_)
  );
  AND2_X1 _43967_ (
    .A1(\cpuregs[23] [27]),
    .A2(_00007_[2]),
    .ZN(_09553_)
  );
  INV_X1 _43968_ (
    .A(_09553_),
    .ZN(_09554_)
  );
  AND2_X1 _43969_ (
    .A1(_09552_),
    .A2(_09554_),
    .ZN(_09555_)
  );
  INV_X1 _43970_ (
    .A(_09555_),
    .ZN(_09556_)
  );
  AND2_X1 _43971_ (
    .A1(_00007_[0]),
    .A2(_09556_),
    .ZN(_09557_)
  );
  INV_X1 _43972_ (
    .A(_09557_),
    .ZN(_09558_)
  );
  AND2_X1 _43973_ (
    .A1(_21612_),
    .A2(_22077_),
    .ZN(_09559_)
  );
  INV_X1 _43974_ (
    .A(_09559_),
    .ZN(_09560_)
  );
  AND2_X1 _43975_ (
    .A1(_21432_),
    .A2(_00007_[2]),
    .ZN(_09561_)
  );
  INV_X1 _43976_ (
    .A(_09561_),
    .ZN(_09562_)
  );
  AND2_X1 _43977_ (
    .A1(_22152_),
    .A2(_09562_),
    .ZN(_09563_)
  );
  AND2_X1 _43978_ (
    .A1(_09560_),
    .A2(_09563_),
    .ZN(_09564_)
  );
  INV_X1 _43979_ (
    .A(_09564_),
    .ZN(_09565_)
  );
  AND2_X1 _43980_ (
    .A1(_21508_),
    .A2(_22077_),
    .ZN(_09566_)
  );
  INV_X1 _43981_ (
    .A(_09566_),
    .ZN(_09567_)
  );
  AND2_X1 _43982_ (
    .A1(_21800_),
    .A2(_00007_[2]),
    .ZN(_09568_)
  );
  INV_X1 _43983_ (
    .A(_09568_),
    .ZN(_09569_)
  );
  AND2_X1 _43984_ (
    .A1(_00007_[0]),
    .A2(_09569_),
    .ZN(_09570_)
  );
  AND2_X1 _43985_ (
    .A1(_09567_),
    .A2(_09570_),
    .ZN(_09571_)
  );
  INV_X1 _43986_ (
    .A(_09571_),
    .ZN(_09572_)
  );
  AND2_X1 _43987_ (
    .A1(_21829_),
    .A2(_00007_[2]),
    .ZN(_09573_)
  );
  INV_X1 _43988_ (
    .A(_09573_),
    .ZN(_09574_)
  );
  AND2_X1 _43989_ (
    .A1(_21563_),
    .A2(_22077_),
    .ZN(_09575_)
  );
  INV_X1 _43990_ (
    .A(_09575_),
    .ZN(_09576_)
  );
  AND2_X1 _43991_ (
    .A1(_22152_),
    .A2(_09576_),
    .ZN(_09577_)
  );
  AND2_X1 _43992_ (
    .A1(_09574_),
    .A2(_09577_),
    .ZN(_09578_)
  );
  INV_X1 _43993_ (
    .A(_09578_),
    .ZN(_09579_)
  );
  AND2_X1 _43994_ (
    .A1(\cpuregs[17] [27]),
    .A2(_22077_),
    .ZN(_09580_)
  );
  INV_X1 _43995_ (
    .A(_09580_),
    .ZN(_09581_)
  );
  AND2_X1 _43996_ (
    .A1(\cpuregs[21] [27]),
    .A2(_00007_[2]),
    .ZN(_09582_)
  );
  INV_X1 _43997_ (
    .A(_09582_),
    .ZN(_09583_)
  );
  AND2_X1 _43998_ (
    .A1(_09581_),
    .A2(_09583_),
    .ZN(_09584_)
  );
  INV_X1 _43999_ (
    .A(_09584_),
    .ZN(_09585_)
  );
  AND2_X1 _44000_ (
    .A1(_00007_[0]),
    .A2(_09585_),
    .ZN(_09586_)
  );
  INV_X1 _44001_ (
    .A(_09586_),
    .ZN(_09587_)
  );
  AND2_X1 _44002_ (
    .A1(\cpuregs[16] [27]),
    .A2(_22077_),
    .ZN(_09588_)
  );
  INV_X1 _44003_ (
    .A(_09588_),
    .ZN(_09589_)
  );
  AND2_X1 _44004_ (
    .A1(\cpuregs[20] [27]),
    .A2(_00007_[2]),
    .ZN(_09590_)
  );
  INV_X1 _44005_ (
    .A(_09590_),
    .ZN(_09591_)
  );
  AND2_X1 _44006_ (
    .A1(_09589_),
    .A2(_09591_),
    .ZN(_09592_)
  );
  INV_X1 _44007_ (
    .A(_09592_),
    .ZN(_09593_)
  );
  AND2_X1 _44008_ (
    .A1(_22152_),
    .A2(_09593_),
    .ZN(_09594_)
  );
  INV_X1 _44009_ (
    .A(_09594_),
    .ZN(_09595_)
  );
  AND2_X1 _44010_ (
    .A1(_09587_),
    .A2(_09595_),
    .ZN(_09596_)
  );
  AND2_X1 _44011_ (
    .A1(_21533_),
    .A2(_22077_),
    .ZN(_09597_)
  );
  INV_X1 _44012_ (
    .A(_09597_),
    .ZN(_09598_)
  );
  AND2_X1 _44013_ (
    .A1(_21753_),
    .A2(_00007_[2]),
    .ZN(_09599_)
  );
  INV_X1 _44014_ (
    .A(_09599_),
    .ZN(_09600_)
  );
  AND2_X1 _44015_ (
    .A1(_00007_[0]),
    .A2(_09600_),
    .ZN(_09601_)
  );
  AND2_X1 _44016_ (
    .A1(_09598_),
    .A2(_09601_),
    .ZN(_09602_)
  );
  INV_X1 _44017_ (
    .A(_09602_),
    .ZN(_09603_)
  );
  AND2_X1 _44018_ (
    .A1(_21974_),
    .A2(_22077_),
    .ZN(_09604_)
  );
  INV_X1 _44019_ (
    .A(_09604_),
    .ZN(_09605_)
  );
  AND2_X1 _44020_ (
    .A1(_21690_),
    .A2(_00007_[2]),
    .ZN(_09606_)
  );
  INV_X1 _44021_ (
    .A(_09606_),
    .ZN(_09607_)
  );
  AND2_X1 _44022_ (
    .A1(_09605_),
    .A2(_09607_),
    .ZN(_09608_)
  );
  AND2_X1 _44023_ (
    .A1(_22152_),
    .A2(_09608_),
    .ZN(_09609_)
  );
  INV_X1 _44024_ (
    .A(_09609_),
    .ZN(_09610_)
  );
  AND2_X1 _44025_ (
    .A1(_09603_),
    .A2(_09610_),
    .ZN(_09611_)
  );
  AND2_X1 _44026_ (
    .A1(_22078_),
    .A2(_09611_),
    .ZN(_09612_)
  );
  INV_X1 _44027_ (
    .A(_09612_),
    .ZN(_09613_)
  );
  AND2_X1 _44028_ (
    .A1(_00007_[1]),
    .A2(_09579_),
    .ZN(_09614_)
  );
  AND2_X1 _44029_ (
    .A1(_09572_),
    .A2(_09614_),
    .ZN(_09615_)
  );
  INV_X1 _44030_ (
    .A(_09615_),
    .ZN(_09616_)
  );
  AND2_X1 _44031_ (
    .A1(_09613_),
    .A2(_09616_),
    .ZN(_09617_)
  );
  AND2_X1 _44032_ (
    .A1(_22144_),
    .A2(_09617_),
    .ZN(_09618_)
  );
  INV_X1 _44033_ (
    .A(_09618_),
    .ZN(_09619_)
  );
  AND2_X1 _44034_ (
    .A1(_00007_[1]),
    .A2(_09565_),
    .ZN(_09620_)
  );
  AND2_X1 _44035_ (
    .A1(_09558_),
    .A2(_09620_),
    .ZN(_09621_)
  );
  INV_X1 _44036_ (
    .A(_09621_),
    .ZN(_09622_)
  );
  AND2_X1 _44037_ (
    .A1(_22078_),
    .A2(_09596_),
    .ZN(_09623_)
  );
  INV_X1 _44038_ (
    .A(_09623_),
    .ZN(_09624_)
  );
  AND2_X1 _44039_ (
    .A1(_09622_),
    .A2(_09624_),
    .ZN(_09625_)
  );
  AND2_X1 _44040_ (
    .A1(_00007_[4]),
    .A2(_09625_),
    .ZN(_09626_)
  );
  INV_X1 _44041_ (
    .A(_09626_),
    .ZN(_09627_)
  );
  AND2_X1 _44042_ (
    .A1(_09619_),
    .A2(_09627_),
    .ZN(_09628_)
  );
  AND2_X1 _44043_ (
    .A1(\cpuregs[26] [27]),
    .A2(_22077_),
    .ZN(_09629_)
  );
  INV_X1 _44044_ (
    .A(_09629_),
    .ZN(_09630_)
  );
  AND2_X1 _44045_ (
    .A1(\cpuregs[30] [27]),
    .A2(_00007_[2]),
    .ZN(_09631_)
  );
  INV_X1 _44046_ (
    .A(_09631_),
    .ZN(_09632_)
  );
  AND2_X1 _44047_ (
    .A1(_00007_[1]),
    .A2(_09632_),
    .ZN(_09633_)
  );
  AND2_X1 _44048_ (
    .A1(_09630_),
    .A2(_09633_),
    .ZN(_09634_)
  );
  INV_X1 _44049_ (
    .A(_09634_),
    .ZN(_09635_)
  );
  AND2_X1 _44050_ (
    .A1(\cpuregs[28] [27]),
    .A2(_00007_[2]),
    .ZN(_09636_)
  );
  INV_X1 _44051_ (
    .A(_09636_),
    .ZN(_09637_)
  );
  AND2_X1 _44052_ (
    .A1(\cpuregs[24] [27]),
    .A2(_22077_),
    .ZN(_09638_)
  );
  INV_X1 _44053_ (
    .A(_09638_),
    .ZN(_09639_)
  );
  AND2_X1 _44054_ (
    .A1(_22078_),
    .A2(_09639_),
    .ZN(_09640_)
  );
  AND2_X1 _44055_ (
    .A1(_09637_),
    .A2(_09640_),
    .ZN(_09641_)
  );
  INV_X1 _44056_ (
    .A(_09641_),
    .ZN(_09642_)
  );
  AND2_X1 _44057_ (
    .A1(_22152_),
    .A2(_09642_),
    .ZN(_09643_)
  );
  AND2_X1 _44058_ (
    .A1(_09635_),
    .A2(_09643_),
    .ZN(_09644_)
  );
  INV_X1 _44059_ (
    .A(_09644_),
    .ZN(_09645_)
  );
  AND2_X1 _44060_ (
    .A1(\cpuregs[27] [27]),
    .A2(_22077_),
    .ZN(_09646_)
  );
  INV_X1 _44061_ (
    .A(_09646_),
    .ZN(_09647_)
  );
  AND2_X1 _44062_ (
    .A1(\cpuregs[31] [27]),
    .A2(_00007_[2]),
    .ZN(_09648_)
  );
  INV_X1 _44063_ (
    .A(_09648_),
    .ZN(_09649_)
  );
  AND2_X1 _44064_ (
    .A1(_00007_[1]),
    .A2(_09649_),
    .ZN(_09650_)
  );
  AND2_X1 _44065_ (
    .A1(_09647_),
    .A2(_09650_),
    .ZN(_09651_)
  );
  INV_X1 _44066_ (
    .A(_09651_),
    .ZN(_09652_)
  );
  AND2_X1 _44067_ (
    .A1(\cpuregs[29] [27]),
    .A2(_00007_[2]),
    .ZN(_09653_)
  );
  INV_X1 _44068_ (
    .A(_09653_),
    .ZN(_09654_)
  );
  AND2_X1 _44069_ (
    .A1(\cpuregs[25] [27]),
    .A2(_22077_),
    .ZN(_09655_)
  );
  INV_X1 _44070_ (
    .A(_09655_),
    .ZN(_09656_)
  );
  AND2_X1 _44071_ (
    .A1(_22078_),
    .A2(_09656_),
    .ZN(_09657_)
  );
  AND2_X1 _44072_ (
    .A1(_09654_),
    .A2(_09657_),
    .ZN(_09658_)
  );
  INV_X1 _44073_ (
    .A(_09658_),
    .ZN(_09659_)
  );
  AND2_X1 _44074_ (
    .A1(_00007_[0]),
    .A2(_09659_),
    .ZN(_09660_)
  );
  AND2_X1 _44075_ (
    .A1(_09652_),
    .A2(_09660_),
    .ZN(_09661_)
  );
  INV_X1 _44076_ (
    .A(_09661_),
    .ZN(_09662_)
  );
  AND2_X1 _44077_ (
    .A1(_09645_),
    .A2(_09662_),
    .ZN(_09663_)
  );
  INV_X1 _44078_ (
    .A(_09663_),
    .ZN(_09664_)
  );
  AND2_X1 _44079_ (
    .A1(_00007_[4]),
    .A2(_09664_),
    .ZN(_09665_)
  );
  INV_X1 _44080_ (
    .A(_09665_),
    .ZN(_09666_)
  );
  AND2_X1 _44081_ (
    .A1(\cpuregs[12] [27]),
    .A2(_22078_),
    .ZN(_09667_)
  );
  INV_X1 _44082_ (
    .A(_09667_),
    .ZN(_09668_)
  );
  AND2_X1 _44083_ (
    .A1(\cpuregs[14] [27]),
    .A2(_00007_[1]),
    .ZN(_09669_)
  );
  INV_X1 _44084_ (
    .A(_09669_),
    .ZN(_09670_)
  );
  AND2_X1 _44085_ (
    .A1(_00007_[2]),
    .A2(_09670_),
    .ZN(_09671_)
  );
  AND2_X1 _44086_ (
    .A1(_09668_),
    .A2(_09671_),
    .ZN(_09672_)
  );
  INV_X1 _44087_ (
    .A(_09672_),
    .ZN(_09673_)
  );
  AND2_X1 _44088_ (
    .A1(\cpuregs[8] [27]),
    .A2(_22078_),
    .ZN(_09674_)
  );
  INV_X1 _44089_ (
    .A(_09674_),
    .ZN(_09675_)
  );
  AND2_X1 _44090_ (
    .A1(\cpuregs[10] [27]),
    .A2(_00007_[1]),
    .ZN(_09676_)
  );
  INV_X1 _44091_ (
    .A(_09676_),
    .ZN(_09677_)
  );
  AND2_X1 _44092_ (
    .A1(_22077_),
    .A2(_09677_),
    .ZN(_09678_)
  );
  AND2_X1 _44093_ (
    .A1(_09675_),
    .A2(_09678_),
    .ZN(_09679_)
  );
  INV_X1 _44094_ (
    .A(_09679_),
    .ZN(_09680_)
  );
  AND2_X1 _44095_ (
    .A1(_22152_),
    .A2(_09680_),
    .ZN(_09681_)
  );
  AND2_X1 _44096_ (
    .A1(_09673_),
    .A2(_09681_),
    .ZN(_09682_)
  );
  INV_X1 _44097_ (
    .A(_09682_),
    .ZN(_09683_)
  );
  AND2_X1 _44098_ (
    .A1(\cpuregs[13] [27]),
    .A2(_22078_),
    .ZN(_09684_)
  );
  INV_X1 _44099_ (
    .A(_09684_),
    .ZN(_09685_)
  );
  AND2_X1 _44100_ (
    .A1(\cpuregs[15] [27]),
    .A2(_00007_[1]),
    .ZN(_09686_)
  );
  INV_X1 _44101_ (
    .A(_09686_),
    .ZN(_09687_)
  );
  AND2_X1 _44102_ (
    .A1(_00007_[2]),
    .A2(_09687_),
    .ZN(_09688_)
  );
  AND2_X1 _44103_ (
    .A1(_09685_),
    .A2(_09688_),
    .ZN(_09689_)
  );
  INV_X1 _44104_ (
    .A(_09689_),
    .ZN(_09690_)
  );
  AND2_X1 _44105_ (
    .A1(\cpuregs[9] [27]),
    .A2(_22078_),
    .ZN(_09691_)
  );
  INV_X1 _44106_ (
    .A(_09691_),
    .ZN(_09692_)
  );
  AND2_X1 _44107_ (
    .A1(\cpuregs[11] [27]),
    .A2(_00007_[1]),
    .ZN(_09693_)
  );
  INV_X1 _44108_ (
    .A(_09693_),
    .ZN(_09694_)
  );
  AND2_X1 _44109_ (
    .A1(_22077_),
    .A2(_09694_),
    .ZN(_09695_)
  );
  AND2_X1 _44110_ (
    .A1(_09692_),
    .A2(_09695_),
    .ZN(_09696_)
  );
  INV_X1 _44111_ (
    .A(_09696_),
    .ZN(_09697_)
  );
  AND2_X1 _44112_ (
    .A1(_00007_[0]),
    .A2(_09697_),
    .ZN(_09698_)
  );
  AND2_X1 _44113_ (
    .A1(_09690_),
    .A2(_09698_),
    .ZN(_09699_)
  );
  INV_X1 _44114_ (
    .A(_09699_),
    .ZN(_09700_)
  );
  AND2_X1 _44115_ (
    .A1(_09683_),
    .A2(_09700_),
    .ZN(_09701_)
  );
  INV_X1 _44116_ (
    .A(_09701_),
    .ZN(_09702_)
  );
  AND2_X1 _44117_ (
    .A1(_22144_),
    .A2(_09702_),
    .ZN(_09703_)
  );
  INV_X1 _44118_ (
    .A(_09703_),
    .ZN(_09704_)
  );
  AND2_X1 _44119_ (
    .A1(_00007_[3]),
    .A2(_09704_),
    .ZN(_09705_)
  );
  AND2_X1 _44120_ (
    .A1(_09666_),
    .A2(_09705_),
    .ZN(_09706_)
  );
  INV_X1 _44121_ (
    .A(_09706_),
    .ZN(_09707_)
  );
  AND2_X1 _44122_ (
    .A1(_22109_),
    .A2(_09628_),
    .ZN(_09708_)
  );
  INV_X1 _44123_ (
    .A(_09708_),
    .ZN(_09709_)
  );
  AND2_X1 _44124_ (
    .A1(_09707_),
    .A2(_09709_),
    .ZN(_09710_)
  );
  AND2_X1 _44125_ (
    .A1(_05842_),
    .A2(_09710_),
    .ZN(_09711_)
  );
  INV_X1 _44126_ (
    .A(_09711_),
    .ZN(_09712_)
  );
  AND2_X1 _44127_ (
    .A1(_21227_),
    .A2(_04963_),
    .ZN(_09713_)
  );
  INV_X1 _44128_ (
    .A(_09713_),
    .ZN(_09714_)
  );
  AND2_X1 _44129_ (
    .A1(_04962_),
    .A2(_09712_),
    .ZN(_09715_)
  );
  AND2_X1 _44130_ (
    .A1(_09550_),
    .A2(_09715_),
    .ZN(_09716_)
  );
  INV_X1 _44131_ (
    .A(_09716_),
    .ZN(_09717_)
  );
  AND2_X1 _44132_ (
    .A1(_09714_),
    .A2(_09717_),
    .ZN(_00308_)
  );
  AND2_X1 _44133_ (
    .A1(decoded_imm[28]),
    .A2(_04966_),
    .ZN(_09718_)
  );
  INV_X1 _44134_ (
    .A(_09718_),
    .ZN(_09719_)
  );
  AND2_X1 _44135_ (
    .A1(_21613_),
    .A2(_22077_),
    .ZN(_09720_)
  );
  INV_X1 _44136_ (
    .A(_09720_),
    .ZN(_09721_)
  );
  AND2_X1 _44137_ (
    .A1(_21433_),
    .A2(_00007_[2]),
    .ZN(_09722_)
  );
  INV_X1 _44138_ (
    .A(_09722_),
    .ZN(_09723_)
  );
  AND2_X1 _44139_ (
    .A1(_21391_),
    .A2(_00007_[2]),
    .ZN(_09724_)
  );
  INV_X1 _44140_ (
    .A(_09724_),
    .ZN(_09725_)
  );
  AND2_X1 _44141_ (
    .A1(_21637_),
    .A2(_22077_),
    .ZN(_09726_)
  );
  INV_X1 _44142_ (
    .A(_09726_),
    .ZN(_09727_)
  );
  AND2_X1 _44143_ (
    .A1(\cpuregs[11] [28]),
    .A2(_22077_),
    .ZN(_09728_)
  );
  INV_X1 _44144_ (
    .A(_09728_),
    .ZN(_09729_)
  );
  AND2_X1 _44145_ (
    .A1(\cpuregs[15] [28]),
    .A2(_00007_[2]),
    .ZN(_09730_)
  );
  INV_X1 _44146_ (
    .A(_09730_),
    .ZN(_09731_)
  );
  AND2_X1 _44147_ (
    .A1(_09729_),
    .A2(_09731_),
    .ZN(_09732_)
  );
  INV_X1 _44148_ (
    .A(_09732_),
    .ZN(_09733_)
  );
  AND2_X1 _44149_ (
    .A1(_00007_[0]),
    .A2(_09733_),
    .ZN(_09734_)
  );
  INV_X1 _44150_ (
    .A(_09734_),
    .ZN(_09735_)
  );
  AND2_X1 _44151_ (
    .A1(\cpuregs[14] [28]),
    .A2(_00007_[2]),
    .ZN(_09736_)
  );
  INV_X1 _44152_ (
    .A(_09736_),
    .ZN(_09737_)
  );
  AND2_X1 _44153_ (
    .A1(\cpuregs[10] [28]),
    .A2(_22077_),
    .ZN(_09738_)
  );
  INV_X1 _44154_ (
    .A(_09738_),
    .ZN(_09739_)
  );
  AND2_X1 _44155_ (
    .A1(_09737_),
    .A2(_09739_),
    .ZN(_09740_)
  );
  INV_X1 _44156_ (
    .A(_09740_),
    .ZN(_09741_)
  );
  AND2_X1 _44157_ (
    .A1(_22152_),
    .A2(_09741_),
    .ZN(_09742_)
  );
  INV_X1 _44158_ (
    .A(_09742_),
    .ZN(_09743_)
  );
  AND2_X1 _44159_ (
    .A1(_09735_),
    .A2(_09743_),
    .ZN(_09744_)
  );
  AND2_X1 _44160_ (
    .A1(_21564_),
    .A2(_22077_),
    .ZN(_09745_)
  );
  INV_X1 _44161_ (
    .A(_09745_),
    .ZN(_09746_)
  );
  AND2_X1 _44162_ (
    .A1(_21830_),
    .A2(_00007_[2]),
    .ZN(_09747_)
  );
  INV_X1 _44163_ (
    .A(_09747_),
    .ZN(_09748_)
  );
  AND2_X1 _44164_ (
    .A1(_22152_),
    .A2(_09748_),
    .ZN(_09749_)
  );
  AND2_X1 _44165_ (
    .A1(_09746_),
    .A2(_09749_),
    .ZN(_09750_)
  );
  INV_X1 _44166_ (
    .A(_09750_),
    .ZN(_09751_)
  );
  AND2_X1 _44167_ (
    .A1(_21801_),
    .A2(_00007_[2]),
    .ZN(_09752_)
  );
  INV_X1 _44168_ (
    .A(_09752_),
    .ZN(_09753_)
  );
  AND2_X1 _44169_ (
    .A1(_21509_),
    .A2(_22077_),
    .ZN(_09754_)
  );
  INV_X1 _44170_ (
    .A(_09754_),
    .ZN(_09755_)
  );
  AND2_X1 _44171_ (
    .A1(_00007_[0]),
    .A2(_09755_),
    .ZN(_09756_)
  );
  AND2_X1 _44172_ (
    .A1(_09753_),
    .A2(_09756_),
    .ZN(_09757_)
  );
  INV_X1 _44173_ (
    .A(_09757_),
    .ZN(_09758_)
  );
  AND2_X1 _44174_ (
    .A1(_09751_),
    .A2(_09758_),
    .ZN(_09759_)
  );
  AND2_X1 _44175_ (
    .A1(_21456_),
    .A2(_22077_),
    .ZN(_09760_)
  );
  INV_X1 _44176_ (
    .A(_09760_),
    .ZN(_09761_)
  );
  AND2_X1 _44177_ (
    .A1(_21667_),
    .A2(_00007_[2]),
    .ZN(_09762_)
  );
  INV_X1 _44178_ (
    .A(_09762_),
    .ZN(_09763_)
  );
  AND2_X1 _44179_ (
    .A1(_09761_),
    .A2(_09763_),
    .ZN(_09764_)
  );
  AND2_X1 _44180_ (
    .A1(_21478_),
    .A2(_22077_),
    .ZN(_09765_)
  );
  INV_X1 _44181_ (
    .A(_09765_),
    .ZN(_09766_)
  );
  AND2_X1 _44182_ (
    .A1(_21777_),
    .A2(_00007_[2]),
    .ZN(_09767_)
  );
  INV_X1 _44183_ (
    .A(_09767_),
    .ZN(_09768_)
  );
  AND2_X1 _44184_ (
    .A1(\cpuregs[9] [28]),
    .A2(_22077_),
    .ZN(_09769_)
  );
  INV_X1 _44185_ (
    .A(_09769_),
    .ZN(_09770_)
  );
  AND2_X1 _44186_ (
    .A1(\cpuregs[13] [28]),
    .A2(_00007_[2]),
    .ZN(_09771_)
  );
  INV_X1 _44187_ (
    .A(_09771_),
    .ZN(_09772_)
  );
  AND2_X1 _44188_ (
    .A1(_09770_),
    .A2(_09772_),
    .ZN(_09773_)
  );
  INV_X1 _44189_ (
    .A(_09773_),
    .ZN(_09774_)
  );
  AND2_X1 _44190_ (
    .A1(_00007_[0]),
    .A2(_09774_),
    .ZN(_09775_)
  );
  INV_X1 _44191_ (
    .A(_09775_),
    .ZN(_09776_)
  );
  AND2_X1 _44192_ (
    .A1(\cpuregs[12] [28]),
    .A2(_00007_[2]),
    .ZN(_09777_)
  );
  INV_X1 _44193_ (
    .A(_09777_),
    .ZN(_09778_)
  );
  AND2_X1 _44194_ (
    .A1(\cpuregs[8] [28]),
    .A2(_22077_),
    .ZN(_09779_)
  );
  INV_X1 _44195_ (
    .A(_09779_),
    .ZN(_09780_)
  );
  AND2_X1 _44196_ (
    .A1(_09778_),
    .A2(_09780_),
    .ZN(_09781_)
  );
  INV_X1 _44197_ (
    .A(_09781_),
    .ZN(_09782_)
  );
  AND2_X1 _44198_ (
    .A1(_22152_),
    .A2(_09782_),
    .ZN(_09783_)
  );
  INV_X1 _44199_ (
    .A(_09783_),
    .ZN(_09784_)
  );
  AND2_X1 _44200_ (
    .A1(_09776_),
    .A2(_09784_),
    .ZN(_09785_)
  );
  AND2_X1 _44201_ (
    .A1(_21691_),
    .A2(_00007_[2]),
    .ZN(_09786_)
  );
  INV_X1 _44202_ (
    .A(_09786_),
    .ZN(_09787_)
  );
  AND2_X1 _44203_ (
    .A1(_21975_),
    .A2(_22077_),
    .ZN(_09788_)
  );
  INV_X1 _44204_ (
    .A(_09788_),
    .ZN(_09789_)
  );
  AND2_X1 _44205_ (
    .A1(_09787_),
    .A2(_09789_),
    .ZN(_09790_)
  );
  AND2_X1 _44206_ (
    .A1(_22152_),
    .A2(_09790_),
    .ZN(_09791_)
  );
  INV_X1 _44207_ (
    .A(_09791_),
    .ZN(_09792_)
  );
  AND2_X1 _44208_ (
    .A1(_21534_),
    .A2(_22077_),
    .ZN(_09793_)
  );
  INV_X1 _44209_ (
    .A(_09793_),
    .ZN(_09794_)
  );
  AND2_X1 _44210_ (
    .A1(_21754_),
    .A2(_00007_[2]),
    .ZN(_09795_)
  );
  INV_X1 _44211_ (
    .A(_09795_),
    .ZN(_09796_)
  );
  AND2_X1 _44212_ (
    .A1(_00007_[0]),
    .A2(_09796_),
    .ZN(_09797_)
  );
  AND2_X1 _44213_ (
    .A1(_09794_),
    .A2(_09797_),
    .ZN(_09798_)
  );
  INV_X1 _44214_ (
    .A(_09798_),
    .ZN(_09799_)
  );
  AND2_X1 _44215_ (
    .A1(_09792_),
    .A2(_09799_),
    .ZN(_09800_)
  );
  AND2_X1 _44216_ (
    .A1(_22152_),
    .A2(_09723_),
    .ZN(_09801_)
  );
  AND2_X1 _44217_ (
    .A1(_09721_),
    .A2(_09801_),
    .ZN(_09802_)
  );
  INV_X1 _44218_ (
    .A(_09802_),
    .ZN(_09803_)
  );
  AND2_X1 _44219_ (
    .A1(_00007_[0]),
    .A2(_09725_),
    .ZN(_09804_)
  );
  AND2_X1 _44220_ (
    .A1(_09727_),
    .A2(_09804_),
    .ZN(_09805_)
  );
  INV_X1 _44221_ (
    .A(_09805_),
    .ZN(_09806_)
  );
  AND2_X1 _44222_ (
    .A1(_09803_),
    .A2(_09806_),
    .ZN(_09807_)
  );
  AND2_X1 _44223_ (
    .A1(_00007_[1]),
    .A2(_09807_),
    .ZN(_09808_)
  );
  INV_X1 _44224_ (
    .A(_09808_),
    .ZN(_09809_)
  );
  AND2_X1 _44225_ (
    .A1(_00007_[0]),
    .A2(_09768_),
    .ZN(_09810_)
  );
  AND2_X1 _44226_ (
    .A1(_09766_),
    .A2(_09810_),
    .ZN(_09811_)
  );
  INV_X1 _44227_ (
    .A(_09811_),
    .ZN(_09812_)
  );
  AND2_X1 _44228_ (
    .A1(_22152_),
    .A2(_09764_),
    .ZN(_09813_)
  );
  INV_X1 _44229_ (
    .A(_09813_),
    .ZN(_09814_)
  );
  AND2_X1 _44230_ (
    .A1(_09812_),
    .A2(_09814_),
    .ZN(_09815_)
  );
  AND2_X1 _44231_ (
    .A1(_22078_),
    .A2(_09815_),
    .ZN(_09816_)
  );
  INV_X1 _44232_ (
    .A(_09816_),
    .ZN(_09817_)
  );
  AND2_X1 _44233_ (
    .A1(_22109_),
    .A2(_09817_),
    .ZN(_09818_)
  );
  AND2_X1 _44234_ (
    .A1(_09809_),
    .A2(_09818_),
    .ZN(_09819_)
  );
  INV_X1 _44235_ (
    .A(_09819_),
    .ZN(_09820_)
  );
  AND2_X1 _44236_ (
    .A1(_21935_),
    .A2(_22077_),
    .ZN(_09821_)
  );
  INV_X1 _44237_ (
    .A(_09821_),
    .ZN(_09822_)
  );
  AND2_X1 _44238_ (
    .A1(_21951_),
    .A2(_00007_[2]),
    .ZN(_09823_)
  );
  INV_X1 _44239_ (
    .A(_09823_),
    .ZN(_09824_)
  );
  AND2_X1 _44240_ (
    .A1(_00007_[0]),
    .A2(_09824_),
    .ZN(_09825_)
  );
  AND2_X1 _44241_ (
    .A1(_09822_),
    .A2(_09825_),
    .ZN(_09826_)
  );
  INV_X1 _44242_ (
    .A(_09826_),
    .ZN(_09827_)
  );
  AND2_X1 _44243_ (
    .A1(_21886_),
    .A2(_22077_),
    .ZN(_09828_)
  );
  INV_X1 _44244_ (
    .A(_09828_),
    .ZN(_09829_)
  );
  AND2_X1 _44245_ (
    .A1(_21863_),
    .A2(_00007_[2]),
    .ZN(_09830_)
  );
  INV_X1 _44246_ (
    .A(_09830_),
    .ZN(_09831_)
  );
  AND2_X1 _44247_ (
    .A1(_09829_),
    .A2(_09831_),
    .ZN(_09832_)
  );
  AND2_X1 _44248_ (
    .A1(_22152_),
    .A2(_09832_),
    .ZN(_09833_)
  );
  INV_X1 _44249_ (
    .A(_09833_),
    .ZN(_09834_)
  );
  AND2_X1 _44250_ (
    .A1(_09827_),
    .A2(_09834_),
    .ZN(_09835_)
  );
  AND2_X1 _44251_ (
    .A1(_00007_[1]),
    .A2(_09835_),
    .ZN(_09836_)
  );
  INV_X1 _44252_ (
    .A(_09836_),
    .ZN(_09837_)
  );
  AND2_X1 _44253_ (
    .A1(_21847_),
    .A2(_22077_),
    .ZN(_09838_)
  );
  INV_X1 _44254_ (
    .A(_09838_),
    .ZN(_09839_)
  );
  AND2_X1 _44255_ (
    .A1(_21903_),
    .A2(_00007_[2]),
    .ZN(_09840_)
  );
  INV_X1 _44256_ (
    .A(_09840_),
    .ZN(_09841_)
  );
  AND2_X1 _44257_ (
    .A1(_00007_[0]),
    .A2(_09841_),
    .ZN(_09842_)
  );
  AND2_X1 _44258_ (
    .A1(_09839_),
    .A2(_09842_),
    .ZN(_09843_)
  );
  INV_X1 _44259_ (
    .A(_09843_),
    .ZN(_09844_)
  );
  AND2_X1 _44260_ (
    .A1(_21581_),
    .A2(_22077_),
    .ZN(_09845_)
  );
  INV_X1 _44261_ (
    .A(_09845_),
    .ZN(_09846_)
  );
  AND2_X1 _44262_ (
    .A1(_21919_),
    .A2(_00007_[2]),
    .ZN(_09847_)
  );
  INV_X1 _44263_ (
    .A(_09847_),
    .ZN(_09848_)
  );
  AND2_X1 _44264_ (
    .A1(_09846_),
    .A2(_09848_),
    .ZN(_09849_)
  );
  AND2_X1 _44265_ (
    .A1(_22152_),
    .A2(_09849_),
    .ZN(_09850_)
  );
  INV_X1 _44266_ (
    .A(_09850_),
    .ZN(_09851_)
  );
  AND2_X1 _44267_ (
    .A1(_09844_),
    .A2(_09851_),
    .ZN(_09852_)
  );
  AND2_X1 _44268_ (
    .A1(_22078_),
    .A2(_09852_),
    .ZN(_09853_)
  );
  INV_X1 _44269_ (
    .A(_09853_),
    .ZN(_09854_)
  );
  AND2_X1 _44270_ (
    .A1(_00007_[3]),
    .A2(_09854_),
    .ZN(_09855_)
  );
  AND2_X1 _44271_ (
    .A1(_09837_),
    .A2(_09855_),
    .ZN(_09856_)
  );
  INV_X1 _44272_ (
    .A(_09856_),
    .ZN(_09857_)
  );
  AND2_X1 _44273_ (
    .A1(_00007_[4]),
    .A2(_09857_),
    .ZN(_09858_)
  );
  AND2_X1 _44274_ (
    .A1(_09820_),
    .A2(_09858_),
    .ZN(_09859_)
  );
  INV_X1 _44275_ (
    .A(_09859_),
    .ZN(_09860_)
  );
  AND2_X1 _44276_ (
    .A1(_00007_[1]),
    .A2(_09759_),
    .ZN(_09861_)
  );
  INV_X1 _44277_ (
    .A(_09861_),
    .ZN(_09862_)
  );
  AND2_X1 _44278_ (
    .A1(_22078_),
    .A2(_09800_),
    .ZN(_09863_)
  );
  INV_X1 _44279_ (
    .A(_09863_),
    .ZN(_09864_)
  );
  AND2_X1 _44280_ (
    .A1(_22109_),
    .A2(_09864_),
    .ZN(_09865_)
  );
  AND2_X1 _44281_ (
    .A1(_09862_),
    .A2(_09865_),
    .ZN(_09866_)
  );
  INV_X1 _44282_ (
    .A(_09866_),
    .ZN(_09867_)
  );
  AND2_X1 _44283_ (
    .A1(_00007_[1]),
    .A2(_09744_),
    .ZN(_09868_)
  );
  INV_X1 _44284_ (
    .A(_09868_),
    .ZN(_09869_)
  );
  AND2_X1 _44285_ (
    .A1(_22078_),
    .A2(_09785_),
    .ZN(_09870_)
  );
  INV_X1 _44286_ (
    .A(_09870_),
    .ZN(_09871_)
  );
  AND2_X1 _44287_ (
    .A1(_00007_[3]),
    .A2(_09871_),
    .ZN(_09872_)
  );
  AND2_X1 _44288_ (
    .A1(_09869_),
    .A2(_09872_),
    .ZN(_09873_)
  );
  INV_X1 _44289_ (
    .A(_09873_),
    .ZN(_09874_)
  );
  AND2_X1 _44290_ (
    .A1(_09867_),
    .A2(_09874_),
    .ZN(_09875_)
  );
  AND2_X1 _44291_ (
    .A1(_22144_),
    .A2(_09875_),
    .ZN(_09876_)
  );
  INV_X1 _44292_ (
    .A(_09876_),
    .ZN(_09877_)
  );
  AND2_X1 _44293_ (
    .A1(_09860_),
    .A2(_09877_),
    .ZN(_09878_)
  );
  AND2_X1 _44294_ (
    .A1(_05842_),
    .A2(_09878_),
    .ZN(_09879_)
  );
  INV_X1 _44295_ (
    .A(_09879_),
    .ZN(_09880_)
  );
  AND2_X1 _44296_ (
    .A1(_21228_),
    .A2(_04963_),
    .ZN(_09881_)
  );
  INV_X1 _44297_ (
    .A(_09881_),
    .ZN(_09882_)
  );
  AND2_X1 _44298_ (
    .A1(_04962_),
    .A2(_09880_),
    .ZN(_09883_)
  );
  AND2_X1 _44299_ (
    .A1(_09719_),
    .A2(_09883_),
    .ZN(_09884_)
  );
  INV_X1 _44300_ (
    .A(_09884_),
    .ZN(_09885_)
  );
  AND2_X1 _44301_ (
    .A1(_09882_),
    .A2(_09885_),
    .ZN(_00309_)
  );
  AND2_X1 _44302_ (
    .A1(_21614_),
    .A2(_22077_),
    .ZN(_09886_)
  );
  INV_X1 _44303_ (
    .A(_09886_),
    .ZN(_09887_)
  );
  AND2_X1 _44304_ (
    .A1(_21434_),
    .A2(_00007_[2]),
    .ZN(_09888_)
  );
  INV_X1 _44305_ (
    .A(_09888_),
    .ZN(_09889_)
  );
  AND2_X1 _44306_ (
    .A1(_21392_),
    .A2(_00007_[2]),
    .ZN(_09890_)
  );
  INV_X1 _44307_ (
    .A(_09890_),
    .ZN(_09891_)
  );
  AND2_X1 _44308_ (
    .A1(_21638_),
    .A2(_22077_),
    .ZN(_09892_)
  );
  INV_X1 _44309_ (
    .A(_09892_),
    .ZN(_09893_)
  );
  AND2_X1 _44310_ (
    .A1(_21588_),
    .A2(_22077_),
    .ZN(_09894_)
  );
  INV_X1 _44311_ (
    .A(_09894_),
    .ZN(_09895_)
  );
  AND2_X1 _44312_ (
    .A1(_21406_),
    .A2(_00007_[2]),
    .ZN(_09896_)
  );
  INV_X1 _44313_ (
    .A(_09896_),
    .ZN(_09897_)
  );
  AND2_X1 _44314_ (
    .A1(_00007_[0]),
    .A2(_09897_),
    .ZN(_09898_)
  );
  AND2_X1 _44315_ (
    .A1(_09895_),
    .A2(_09898_),
    .ZN(_09899_)
  );
  INV_X1 _44316_ (
    .A(_09899_),
    .ZN(_09900_)
  );
  AND2_X1 _44317_ (
    .A1(\cpuregs[14] [29]),
    .A2(_00007_[2]),
    .ZN(_09901_)
  );
  INV_X1 _44318_ (
    .A(_09901_),
    .ZN(_09902_)
  );
  AND2_X1 _44319_ (
    .A1(\cpuregs[10] [29]),
    .A2(_22077_),
    .ZN(_09903_)
  );
  INV_X1 _44320_ (
    .A(_09903_),
    .ZN(_09904_)
  );
  AND2_X1 _44321_ (
    .A1(_09902_),
    .A2(_09904_),
    .ZN(_09905_)
  );
  INV_X1 _44322_ (
    .A(_09905_),
    .ZN(_09906_)
  );
  AND2_X1 _44323_ (
    .A1(_22152_),
    .A2(_09906_),
    .ZN(_09907_)
  );
  INV_X1 _44324_ (
    .A(_09907_),
    .ZN(_09908_)
  );
  AND2_X1 _44325_ (
    .A1(_09900_),
    .A2(_09908_),
    .ZN(_09909_)
  );
  AND2_X1 _44326_ (
    .A1(_21565_),
    .A2(_22077_),
    .ZN(_09910_)
  );
  INV_X1 _44327_ (
    .A(_09910_),
    .ZN(_09911_)
  );
  AND2_X1 _44328_ (
    .A1(_21831_),
    .A2(_00007_[2]),
    .ZN(_09912_)
  );
  INV_X1 _44329_ (
    .A(_09912_),
    .ZN(_09913_)
  );
  AND2_X1 _44330_ (
    .A1(_22152_),
    .A2(_09913_),
    .ZN(_09914_)
  );
  AND2_X1 _44331_ (
    .A1(_09911_),
    .A2(_09914_),
    .ZN(_09915_)
  );
  INV_X1 _44332_ (
    .A(_09915_),
    .ZN(_09916_)
  );
  AND2_X1 _44333_ (
    .A1(_21802_),
    .A2(_00007_[2]),
    .ZN(_09917_)
  );
  INV_X1 _44334_ (
    .A(_09917_),
    .ZN(_09918_)
  );
  AND2_X1 _44335_ (
    .A1(_21510_),
    .A2(_22077_),
    .ZN(_09919_)
  );
  INV_X1 _44336_ (
    .A(_09919_),
    .ZN(_09920_)
  );
  AND2_X1 _44337_ (
    .A1(_00007_[0]),
    .A2(_09920_),
    .ZN(_09921_)
  );
  AND2_X1 _44338_ (
    .A1(_09918_),
    .A2(_09921_),
    .ZN(_09922_)
  );
  INV_X1 _44339_ (
    .A(_09922_),
    .ZN(_09923_)
  );
  AND2_X1 _44340_ (
    .A1(_09916_),
    .A2(_09923_),
    .ZN(_09924_)
  );
  AND2_X1 _44341_ (
    .A1(_21457_),
    .A2(_22077_),
    .ZN(_09925_)
  );
  INV_X1 _44342_ (
    .A(_09925_),
    .ZN(_09926_)
  );
  AND2_X1 _44343_ (
    .A1(_21668_),
    .A2(_00007_[2]),
    .ZN(_09927_)
  );
  INV_X1 _44344_ (
    .A(_09927_),
    .ZN(_09928_)
  );
  AND2_X1 _44345_ (
    .A1(_09926_),
    .A2(_09928_),
    .ZN(_09929_)
  );
  AND2_X1 _44346_ (
    .A1(_21479_),
    .A2(_22077_),
    .ZN(_09930_)
  );
  INV_X1 _44347_ (
    .A(_09930_),
    .ZN(_09931_)
  );
  AND2_X1 _44348_ (
    .A1(_21778_),
    .A2(_00007_[2]),
    .ZN(_09932_)
  );
  INV_X1 _44349_ (
    .A(_09932_),
    .ZN(_09933_)
  );
  AND2_X1 _44350_ (
    .A1(_21723_),
    .A2(_22077_),
    .ZN(_09934_)
  );
  INV_X1 _44351_ (
    .A(_09934_),
    .ZN(_09935_)
  );
  AND2_X1 _44352_ (
    .A1(_21645_),
    .A2(_00007_[2]),
    .ZN(_09936_)
  );
  INV_X1 _44353_ (
    .A(_09936_),
    .ZN(_09937_)
  );
  AND2_X1 _44354_ (
    .A1(_00007_[0]),
    .A2(_09937_),
    .ZN(_09938_)
  );
  AND2_X1 _44355_ (
    .A1(_09935_),
    .A2(_09938_),
    .ZN(_09939_)
  );
  INV_X1 _44356_ (
    .A(_09939_),
    .ZN(_09940_)
  );
  AND2_X1 _44357_ (
    .A1(\cpuregs[12] [29]),
    .A2(_00007_[2]),
    .ZN(_09941_)
  );
  INV_X1 _44358_ (
    .A(_09941_),
    .ZN(_09942_)
  );
  AND2_X1 _44359_ (
    .A1(\cpuregs[8] [29]),
    .A2(_22077_),
    .ZN(_09943_)
  );
  INV_X1 _44360_ (
    .A(_09943_),
    .ZN(_09944_)
  );
  AND2_X1 _44361_ (
    .A1(_09942_),
    .A2(_09944_),
    .ZN(_09945_)
  );
  INV_X1 _44362_ (
    .A(_09945_),
    .ZN(_09946_)
  );
  AND2_X1 _44363_ (
    .A1(_22152_),
    .A2(_09946_),
    .ZN(_09947_)
  );
  INV_X1 _44364_ (
    .A(_09947_),
    .ZN(_09948_)
  );
  AND2_X1 _44365_ (
    .A1(_09940_),
    .A2(_09948_),
    .ZN(_09949_)
  );
  AND2_X1 _44366_ (
    .A1(_21692_),
    .A2(_00007_[2]),
    .ZN(_09950_)
  );
  INV_X1 _44367_ (
    .A(_09950_),
    .ZN(_09951_)
  );
  AND2_X1 _44368_ (
    .A1(_21976_),
    .A2(_22077_),
    .ZN(_09952_)
  );
  INV_X1 _44369_ (
    .A(_09952_),
    .ZN(_09953_)
  );
  AND2_X1 _44370_ (
    .A1(_09951_),
    .A2(_09953_),
    .ZN(_09954_)
  );
  AND2_X1 _44371_ (
    .A1(_22152_),
    .A2(_09954_),
    .ZN(_09955_)
  );
  INV_X1 _44372_ (
    .A(_09955_),
    .ZN(_09956_)
  );
  AND2_X1 _44373_ (
    .A1(_21535_),
    .A2(_22077_),
    .ZN(_09957_)
  );
  INV_X1 _44374_ (
    .A(_09957_),
    .ZN(_09958_)
  );
  AND2_X1 _44375_ (
    .A1(_21755_),
    .A2(_00007_[2]),
    .ZN(_09959_)
  );
  INV_X1 _44376_ (
    .A(_09959_),
    .ZN(_09960_)
  );
  AND2_X1 _44377_ (
    .A1(_00007_[0]),
    .A2(_09960_),
    .ZN(_09961_)
  );
  AND2_X1 _44378_ (
    .A1(_09958_),
    .A2(_09961_),
    .ZN(_09962_)
  );
  INV_X1 _44379_ (
    .A(_09962_),
    .ZN(_09963_)
  );
  AND2_X1 _44380_ (
    .A1(_09956_),
    .A2(_09963_),
    .ZN(_09964_)
  );
  AND2_X1 _44381_ (
    .A1(_22152_),
    .A2(_09889_),
    .ZN(_09965_)
  );
  AND2_X1 _44382_ (
    .A1(_09887_),
    .A2(_09965_),
    .ZN(_09966_)
  );
  INV_X1 _44383_ (
    .A(_09966_),
    .ZN(_09967_)
  );
  AND2_X1 _44384_ (
    .A1(_00007_[0]),
    .A2(_09891_),
    .ZN(_09968_)
  );
  AND2_X1 _44385_ (
    .A1(_09893_),
    .A2(_09968_),
    .ZN(_09969_)
  );
  INV_X1 _44386_ (
    .A(_09969_),
    .ZN(_09970_)
  );
  AND2_X1 _44387_ (
    .A1(_09967_),
    .A2(_09970_),
    .ZN(_09971_)
  );
  AND2_X1 _44388_ (
    .A1(_00007_[1]),
    .A2(_09971_),
    .ZN(_09972_)
  );
  INV_X1 _44389_ (
    .A(_09972_),
    .ZN(_09973_)
  );
  AND2_X1 _44390_ (
    .A1(_00007_[0]),
    .A2(_09933_),
    .ZN(_09974_)
  );
  AND2_X1 _44391_ (
    .A1(_09931_),
    .A2(_09974_),
    .ZN(_09975_)
  );
  INV_X1 _44392_ (
    .A(_09975_),
    .ZN(_09976_)
  );
  AND2_X1 _44393_ (
    .A1(_22152_),
    .A2(_09929_),
    .ZN(_09977_)
  );
  INV_X1 _44394_ (
    .A(_09977_),
    .ZN(_09978_)
  );
  AND2_X1 _44395_ (
    .A1(_09976_),
    .A2(_09978_),
    .ZN(_09979_)
  );
  AND2_X1 _44396_ (
    .A1(_22078_),
    .A2(_09979_),
    .ZN(_09980_)
  );
  INV_X1 _44397_ (
    .A(_09980_),
    .ZN(_09981_)
  );
  AND2_X1 _44398_ (
    .A1(_22109_),
    .A2(_09981_),
    .ZN(_09982_)
  );
  AND2_X1 _44399_ (
    .A1(_09973_),
    .A2(_09982_),
    .ZN(_09983_)
  );
  INV_X1 _44400_ (
    .A(_09983_),
    .ZN(_09984_)
  );
  AND2_X1 _44401_ (
    .A1(_21936_),
    .A2(_22077_),
    .ZN(_09985_)
  );
  INV_X1 _44402_ (
    .A(_09985_),
    .ZN(_09986_)
  );
  AND2_X1 _44403_ (
    .A1(_21952_),
    .A2(_00007_[2]),
    .ZN(_09987_)
  );
  INV_X1 _44404_ (
    .A(_09987_),
    .ZN(_09988_)
  );
  AND2_X1 _44405_ (
    .A1(_00007_[0]),
    .A2(_09988_),
    .ZN(_09989_)
  );
  AND2_X1 _44406_ (
    .A1(_09986_),
    .A2(_09989_),
    .ZN(_09990_)
  );
  INV_X1 _44407_ (
    .A(_09990_),
    .ZN(_09991_)
  );
  AND2_X1 _44408_ (
    .A1(_21887_),
    .A2(_22077_),
    .ZN(_09992_)
  );
  INV_X1 _44409_ (
    .A(_09992_),
    .ZN(_09993_)
  );
  AND2_X1 _44410_ (
    .A1(_21864_),
    .A2(_00007_[2]),
    .ZN(_09994_)
  );
  INV_X1 _44411_ (
    .A(_09994_),
    .ZN(_09995_)
  );
  AND2_X1 _44412_ (
    .A1(_09993_),
    .A2(_09995_),
    .ZN(_09996_)
  );
  AND2_X1 _44413_ (
    .A1(_22152_),
    .A2(_09996_),
    .ZN(_09997_)
  );
  INV_X1 _44414_ (
    .A(_09997_),
    .ZN(_09998_)
  );
  AND2_X1 _44415_ (
    .A1(_09991_),
    .A2(_09998_),
    .ZN(_09999_)
  );
  AND2_X1 _44416_ (
    .A1(_00007_[1]),
    .A2(_09999_),
    .ZN(_10000_)
  );
  INV_X1 _44417_ (
    .A(_10000_),
    .ZN(_10001_)
  );
  AND2_X1 _44418_ (
    .A1(_21848_),
    .A2(_22077_),
    .ZN(_10002_)
  );
  INV_X1 _44419_ (
    .A(_10002_),
    .ZN(_10003_)
  );
  AND2_X1 _44420_ (
    .A1(_21904_),
    .A2(_00007_[2]),
    .ZN(_10004_)
  );
  INV_X1 _44421_ (
    .A(_10004_),
    .ZN(_10005_)
  );
  AND2_X1 _44422_ (
    .A1(_00007_[0]),
    .A2(_10005_),
    .ZN(_10006_)
  );
  AND2_X1 _44423_ (
    .A1(_10003_),
    .A2(_10006_),
    .ZN(_10007_)
  );
  INV_X1 _44424_ (
    .A(_10007_),
    .ZN(_10008_)
  );
  AND2_X1 _44425_ (
    .A1(_21582_),
    .A2(_22077_),
    .ZN(_10009_)
  );
  INV_X1 _44426_ (
    .A(_10009_),
    .ZN(_10010_)
  );
  AND2_X1 _44427_ (
    .A1(_21920_),
    .A2(_00007_[2]),
    .ZN(_10011_)
  );
  INV_X1 _44428_ (
    .A(_10011_),
    .ZN(_10012_)
  );
  AND2_X1 _44429_ (
    .A1(_10010_),
    .A2(_10012_),
    .ZN(_10013_)
  );
  AND2_X1 _44430_ (
    .A1(_22152_),
    .A2(_10013_),
    .ZN(_10014_)
  );
  INV_X1 _44431_ (
    .A(_10014_),
    .ZN(_10015_)
  );
  AND2_X1 _44432_ (
    .A1(_10008_),
    .A2(_10015_),
    .ZN(_10016_)
  );
  AND2_X1 _44433_ (
    .A1(_22078_),
    .A2(_10016_),
    .ZN(_10017_)
  );
  INV_X1 _44434_ (
    .A(_10017_),
    .ZN(_10018_)
  );
  AND2_X1 _44435_ (
    .A1(_00007_[3]),
    .A2(_10018_),
    .ZN(_10019_)
  );
  AND2_X1 _44436_ (
    .A1(_10001_),
    .A2(_10019_),
    .ZN(_10020_)
  );
  INV_X1 _44437_ (
    .A(_10020_),
    .ZN(_10021_)
  );
  AND2_X1 _44438_ (
    .A1(_00007_[4]),
    .A2(_10021_),
    .ZN(_10022_)
  );
  AND2_X1 _44439_ (
    .A1(_09984_),
    .A2(_10022_),
    .ZN(_10023_)
  );
  INV_X1 _44440_ (
    .A(_10023_),
    .ZN(_10024_)
  );
  AND2_X1 _44441_ (
    .A1(_00007_[1]),
    .A2(_09924_),
    .ZN(_10025_)
  );
  INV_X1 _44442_ (
    .A(_10025_),
    .ZN(_10026_)
  );
  AND2_X1 _44443_ (
    .A1(_22078_),
    .A2(_09964_),
    .ZN(_10027_)
  );
  INV_X1 _44444_ (
    .A(_10027_),
    .ZN(_10028_)
  );
  AND2_X1 _44445_ (
    .A1(_22109_),
    .A2(_10028_),
    .ZN(_10029_)
  );
  AND2_X1 _44446_ (
    .A1(_10026_),
    .A2(_10029_),
    .ZN(_10030_)
  );
  INV_X1 _44447_ (
    .A(_10030_),
    .ZN(_10031_)
  );
  AND2_X1 _44448_ (
    .A1(_00007_[1]),
    .A2(_09909_),
    .ZN(_10032_)
  );
  INV_X1 _44449_ (
    .A(_10032_),
    .ZN(_10033_)
  );
  AND2_X1 _44450_ (
    .A1(_22078_),
    .A2(_09949_),
    .ZN(_10034_)
  );
  INV_X1 _44451_ (
    .A(_10034_),
    .ZN(_10035_)
  );
  AND2_X1 _44452_ (
    .A1(_00007_[3]),
    .A2(_10035_),
    .ZN(_10036_)
  );
  AND2_X1 _44453_ (
    .A1(_10033_),
    .A2(_10036_),
    .ZN(_10037_)
  );
  INV_X1 _44454_ (
    .A(_10037_),
    .ZN(_10038_)
  );
  AND2_X1 _44455_ (
    .A1(_10031_),
    .A2(_10038_),
    .ZN(_10039_)
  );
  AND2_X1 _44456_ (
    .A1(_22144_),
    .A2(_10039_),
    .ZN(_10040_)
  );
  INV_X1 _44457_ (
    .A(_10040_),
    .ZN(_10041_)
  );
  AND2_X1 _44458_ (
    .A1(_10024_),
    .A2(_10041_),
    .ZN(_10042_)
  );
  AND2_X1 _44459_ (
    .A1(_05842_),
    .A2(_10042_),
    .ZN(_10043_)
  );
  INV_X1 _44460_ (
    .A(_10043_),
    .ZN(_10044_)
  );
  AND2_X1 _44461_ (
    .A1(decoded_imm[29]),
    .A2(_04966_),
    .ZN(_10045_)
  );
  INV_X1 _44462_ (
    .A(_10045_),
    .ZN(_10046_)
  );
  AND2_X1 _44463_ (
    .A1(_21229_),
    .A2(_04963_),
    .ZN(_10047_)
  );
  INV_X1 _44464_ (
    .A(_10047_),
    .ZN(_10048_)
  );
  AND2_X1 _44465_ (
    .A1(_04962_),
    .A2(_10046_),
    .ZN(_10049_)
  );
  AND2_X1 _44466_ (
    .A1(_10044_),
    .A2(_10049_),
    .ZN(_10050_)
  );
  INV_X1 _44467_ (
    .A(_10050_),
    .ZN(_10051_)
  );
  AND2_X1 _44468_ (
    .A1(_10048_),
    .A2(_10051_),
    .ZN(_00310_)
  );
  AND2_X1 _44469_ (
    .A1(decoded_imm[30]),
    .A2(_04966_),
    .ZN(_10052_)
  );
  INV_X1 _44470_ (
    .A(_10052_),
    .ZN(_10053_)
  );
  AND2_X1 _44471_ (
    .A1(\cpuregs[19] [30]),
    .A2(_22077_),
    .ZN(_10054_)
  );
  INV_X1 _44472_ (
    .A(_10054_),
    .ZN(_10055_)
  );
  AND2_X1 _44473_ (
    .A1(\cpuregs[23] [30]),
    .A2(_00007_[2]),
    .ZN(_10056_)
  );
  INV_X1 _44474_ (
    .A(_10056_),
    .ZN(_10057_)
  );
  AND2_X1 _44475_ (
    .A1(_10055_),
    .A2(_10057_),
    .ZN(_10058_)
  );
  INV_X1 _44476_ (
    .A(_10058_),
    .ZN(_10059_)
  );
  AND2_X1 _44477_ (
    .A1(_00007_[0]),
    .A2(_10059_),
    .ZN(_10060_)
  );
  INV_X1 _44478_ (
    .A(_10060_),
    .ZN(_10061_)
  );
  AND2_X1 _44479_ (
    .A1(_21615_),
    .A2(_22077_),
    .ZN(_10062_)
  );
  INV_X1 _44480_ (
    .A(_10062_),
    .ZN(_10063_)
  );
  AND2_X1 _44481_ (
    .A1(_21435_),
    .A2(_00007_[2]),
    .ZN(_10064_)
  );
  INV_X1 _44482_ (
    .A(_10064_),
    .ZN(_10065_)
  );
  AND2_X1 _44483_ (
    .A1(_22152_),
    .A2(_10065_),
    .ZN(_10066_)
  );
  AND2_X1 _44484_ (
    .A1(_10063_),
    .A2(_10066_),
    .ZN(_10067_)
  );
  INV_X1 _44485_ (
    .A(_10067_),
    .ZN(_10068_)
  );
  AND2_X1 _44486_ (
    .A1(_21511_),
    .A2(_22077_),
    .ZN(_10069_)
  );
  INV_X1 _44487_ (
    .A(_10069_),
    .ZN(_10070_)
  );
  AND2_X1 _44488_ (
    .A1(_21803_),
    .A2(_00007_[2]),
    .ZN(_10071_)
  );
  INV_X1 _44489_ (
    .A(_10071_),
    .ZN(_10072_)
  );
  AND2_X1 _44490_ (
    .A1(_00007_[0]),
    .A2(_10072_),
    .ZN(_10073_)
  );
  AND2_X1 _44491_ (
    .A1(_10070_),
    .A2(_10073_),
    .ZN(_10074_)
  );
  INV_X1 _44492_ (
    .A(_10074_),
    .ZN(_10075_)
  );
  AND2_X1 _44493_ (
    .A1(_21832_),
    .A2(_00007_[2]),
    .ZN(_10076_)
  );
  INV_X1 _44494_ (
    .A(_10076_),
    .ZN(_10077_)
  );
  AND2_X1 _44495_ (
    .A1(_21566_),
    .A2(_22077_),
    .ZN(_10078_)
  );
  INV_X1 _44496_ (
    .A(_10078_),
    .ZN(_10079_)
  );
  AND2_X1 _44497_ (
    .A1(_22152_),
    .A2(_10079_),
    .ZN(_10080_)
  );
  AND2_X1 _44498_ (
    .A1(_10077_),
    .A2(_10080_),
    .ZN(_10081_)
  );
  INV_X1 _44499_ (
    .A(_10081_),
    .ZN(_10082_)
  );
  AND2_X1 _44500_ (
    .A1(\cpuregs[17] [30]),
    .A2(_22077_),
    .ZN(_10083_)
  );
  INV_X1 _44501_ (
    .A(_10083_),
    .ZN(_10084_)
  );
  AND2_X1 _44502_ (
    .A1(\cpuregs[21] [30]),
    .A2(_00007_[2]),
    .ZN(_10085_)
  );
  INV_X1 _44503_ (
    .A(_10085_),
    .ZN(_10086_)
  );
  AND2_X1 _44504_ (
    .A1(_10084_),
    .A2(_10086_),
    .ZN(_10087_)
  );
  INV_X1 _44505_ (
    .A(_10087_),
    .ZN(_10088_)
  );
  AND2_X1 _44506_ (
    .A1(_00007_[0]),
    .A2(_10088_),
    .ZN(_10089_)
  );
  INV_X1 _44507_ (
    .A(_10089_),
    .ZN(_10090_)
  );
  AND2_X1 _44508_ (
    .A1(\cpuregs[16] [30]),
    .A2(_22077_),
    .ZN(_10091_)
  );
  INV_X1 _44509_ (
    .A(_10091_),
    .ZN(_10092_)
  );
  AND2_X1 _44510_ (
    .A1(\cpuregs[20] [30]),
    .A2(_00007_[2]),
    .ZN(_10093_)
  );
  INV_X1 _44511_ (
    .A(_10093_),
    .ZN(_10094_)
  );
  AND2_X1 _44512_ (
    .A1(_10092_),
    .A2(_10094_),
    .ZN(_10095_)
  );
  INV_X1 _44513_ (
    .A(_10095_),
    .ZN(_10096_)
  );
  AND2_X1 _44514_ (
    .A1(_22152_),
    .A2(_10096_),
    .ZN(_10097_)
  );
  INV_X1 _44515_ (
    .A(_10097_),
    .ZN(_10098_)
  );
  AND2_X1 _44516_ (
    .A1(_10090_),
    .A2(_10098_),
    .ZN(_10099_)
  );
  AND2_X1 _44517_ (
    .A1(_21536_),
    .A2(_22077_),
    .ZN(_10100_)
  );
  INV_X1 _44518_ (
    .A(_10100_),
    .ZN(_10101_)
  );
  AND2_X1 _44519_ (
    .A1(_21756_),
    .A2(_00007_[2]),
    .ZN(_10102_)
  );
  INV_X1 _44520_ (
    .A(_10102_),
    .ZN(_10103_)
  );
  AND2_X1 _44521_ (
    .A1(_00007_[0]),
    .A2(_10103_),
    .ZN(_10104_)
  );
  AND2_X1 _44522_ (
    .A1(_10101_),
    .A2(_10104_),
    .ZN(_10105_)
  );
  INV_X1 _44523_ (
    .A(_10105_),
    .ZN(_10106_)
  );
  AND2_X1 _44524_ (
    .A1(_21977_),
    .A2(_22077_),
    .ZN(_10107_)
  );
  INV_X1 _44525_ (
    .A(_10107_),
    .ZN(_10108_)
  );
  AND2_X1 _44526_ (
    .A1(_21693_),
    .A2(_00007_[2]),
    .ZN(_10109_)
  );
  INV_X1 _44527_ (
    .A(_10109_),
    .ZN(_10110_)
  );
  AND2_X1 _44528_ (
    .A1(_10108_),
    .A2(_10110_),
    .ZN(_10111_)
  );
  AND2_X1 _44529_ (
    .A1(_22152_),
    .A2(_10111_),
    .ZN(_10112_)
  );
  INV_X1 _44530_ (
    .A(_10112_),
    .ZN(_10113_)
  );
  AND2_X1 _44531_ (
    .A1(_10106_),
    .A2(_10113_),
    .ZN(_10114_)
  );
  AND2_X1 _44532_ (
    .A1(_22078_),
    .A2(_10114_),
    .ZN(_10115_)
  );
  INV_X1 _44533_ (
    .A(_10115_),
    .ZN(_10116_)
  );
  AND2_X1 _44534_ (
    .A1(_00007_[1]),
    .A2(_10082_),
    .ZN(_10117_)
  );
  AND2_X1 _44535_ (
    .A1(_10075_),
    .A2(_10117_),
    .ZN(_10118_)
  );
  INV_X1 _44536_ (
    .A(_10118_),
    .ZN(_10119_)
  );
  AND2_X1 _44537_ (
    .A1(_10116_),
    .A2(_10119_),
    .ZN(_10120_)
  );
  AND2_X1 _44538_ (
    .A1(_22144_),
    .A2(_10120_),
    .ZN(_10121_)
  );
  INV_X1 _44539_ (
    .A(_10121_),
    .ZN(_10122_)
  );
  AND2_X1 _44540_ (
    .A1(_00007_[1]),
    .A2(_10068_),
    .ZN(_10123_)
  );
  AND2_X1 _44541_ (
    .A1(_10061_),
    .A2(_10123_),
    .ZN(_10124_)
  );
  INV_X1 _44542_ (
    .A(_10124_),
    .ZN(_10125_)
  );
  AND2_X1 _44543_ (
    .A1(_22078_),
    .A2(_10099_),
    .ZN(_10126_)
  );
  INV_X1 _44544_ (
    .A(_10126_),
    .ZN(_10127_)
  );
  AND2_X1 _44545_ (
    .A1(_10125_),
    .A2(_10127_),
    .ZN(_10128_)
  );
  AND2_X1 _44546_ (
    .A1(_00007_[4]),
    .A2(_10128_),
    .ZN(_10129_)
  );
  INV_X1 _44547_ (
    .A(_10129_),
    .ZN(_10130_)
  );
  AND2_X1 _44548_ (
    .A1(_10122_),
    .A2(_10130_),
    .ZN(_10131_)
  );
  AND2_X1 _44549_ (
    .A1(\cpuregs[26] [30]),
    .A2(_22077_),
    .ZN(_10132_)
  );
  INV_X1 _44550_ (
    .A(_10132_),
    .ZN(_10133_)
  );
  AND2_X1 _44551_ (
    .A1(\cpuregs[30] [30]),
    .A2(_00007_[2]),
    .ZN(_10134_)
  );
  INV_X1 _44552_ (
    .A(_10134_),
    .ZN(_10135_)
  );
  AND2_X1 _44553_ (
    .A1(_00007_[1]),
    .A2(_10135_),
    .ZN(_10136_)
  );
  AND2_X1 _44554_ (
    .A1(_10133_),
    .A2(_10136_),
    .ZN(_10137_)
  );
  INV_X1 _44555_ (
    .A(_10137_),
    .ZN(_10138_)
  );
  AND2_X1 _44556_ (
    .A1(\cpuregs[28] [30]),
    .A2(_00007_[2]),
    .ZN(_10139_)
  );
  INV_X1 _44557_ (
    .A(_10139_),
    .ZN(_10140_)
  );
  AND2_X1 _44558_ (
    .A1(\cpuregs[24] [30]),
    .A2(_22077_),
    .ZN(_10141_)
  );
  INV_X1 _44559_ (
    .A(_10141_),
    .ZN(_10142_)
  );
  AND2_X1 _44560_ (
    .A1(_22078_),
    .A2(_10142_),
    .ZN(_10143_)
  );
  AND2_X1 _44561_ (
    .A1(_10140_),
    .A2(_10143_),
    .ZN(_10144_)
  );
  INV_X1 _44562_ (
    .A(_10144_),
    .ZN(_10145_)
  );
  AND2_X1 _44563_ (
    .A1(_22152_),
    .A2(_10145_),
    .ZN(_10146_)
  );
  AND2_X1 _44564_ (
    .A1(_10138_),
    .A2(_10146_),
    .ZN(_10147_)
  );
  INV_X1 _44565_ (
    .A(_10147_),
    .ZN(_10148_)
  );
  AND2_X1 _44566_ (
    .A1(\cpuregs[27] [30]),
    .A2(_22077_),
    .ZN(_10149_)
  );
  INV_X1 _44567_ (
    .A(_10149_),
    .ZN(_10150_)
  );
  AND2_X1 _44568_ (
    .A1(\cpuregs[31] [30]),
    .A2(_00007_[2]),
    .ZN(_10151_)
  );
  INV_X1 _44569_ (
    .A(_10151_),
    .ZN(_10152_)
  );
  AND2_X1 _44570_ (
    .A1(_00007_[1]),
    .A2(_10152_),
    .ZN(_10153_)
  );
  AND2_X1 _44571_ (
    .A1(_10150_),
    .A2(_10153_),
    .ZN(_10154_)
  );
  INV_X1 _44572_ (
    .A(_10154_),
    .ZN(_10155_)
  );
  AND2_X1 _44573_ (
    .A1(\cpuregs[29] [30]),
    .A2(_00007_[2]),
    .ZN(_10156_)
  );
  INV_X1 _44574_ (
    .A(_10156_),
    .ZN(_10157_)
  );
  AND2_X1 _44575_ (
    .A1(\cpuregs[25] [30]),
    .A2(_22077_),
    .ZN(_10158_)
  );
  INV_X1 _44576_ (
    .A(_10158_),
    .ZN(_10159_)
  );
  AND2_X1 _44577_ (
    .A1(_22078_),
    .A2(_10159_),
    .ZN(_10160_)
  );
  AND2_X1 _44578_ (
    .A1(_10157_),
    .A2(_10160_),
    .ZN(_10161_)
  );
  INV_X1 _44579_ (
    .A(_10161_),
    .ZN(_10162_)
  );
  AND2_X1 _44580_ (
    .A1(_00007_[0]),
    .A2(_10162_),
    .ZN(_10163_)
  );
  AND2_X1 _44581_ (
    .A1(_10155_),
    .A2(_10163_),
    .ZN(_10164_)
  );
  INV_X1 _44582_ (
    .A(_10164_),
    .ZN(_10165_)
  );
  AND2_X1 _44583_ (
    .A1(_10148_),
    .A2(_10165_),
    .ZN(_10166_)
  );
  INV_X1 _44584_ (
    .A(_10166_),
    .ZN(_10167_)
  );
  AND2_X1 _44585_ (
    .A1(_00007_[4]),
    .A2(_10167_),
    .ZN(_10168_)
  );
  INV_X1 _44586_ (
    .A(_10168_),
    .ZN(_10169_)
  );
  AND2_X1 _44587_ (
    .A1(_21646_),
    .A2(_00007_[2]),
    .ZN(_10170_)
  );
  INV_X1 _44588_ (
    .A(_10170_),
    .ZN(_10171_)
  );
  AND2_X1 _44589_ (
    .A1(_21724_),
    .A2(_22077_),
    .ZN(_10172_)
  );
  INV_X1 _44590_ (
    .A(_10172_),
    .ZN(_10173_)
  );
  AND2_X1 _44591_ (
    .A1(_00007_[0]),
    .A2(_10173_),
    .ZN(_10174_)
  );
  AND2_X1 _44592_ (
    .A1(_10171_),
    .A2(_10174_),
    .ZN(_10175_)
  );
  INV_X1 _44593_ (
    .A(_10175_),
    .ZN(_10176_)
  );
  AND2_X1 _44594_ (
    .A1(_21731_),
    .A2(_22077_),
    .ZN(_10177_)
  );
  INV_X1 _44595_ (
    .A(_10177_),
    .ZN(_10178_)
  );
  AND2_X1 _44596_ (
    .A1(_21486_),
    .A2(_00007_[2]),
    .ZN(_10179_)
  );
  INV_X1 _44597_ (
    .A(_10179_),
    .ZN(_10180_)
  );
  AND2_X1 _44598_ (
    .A1(_10178_),
    .A2(_10180_),
    .ZN(_10181_)
  );
  AND2_X1 _44599_ (
    .A1(_22152_),
    .A2(_10181_),
    .ZN(_10182_)
  );
  INV_X1 _44600_ (
    .A(_10182_),
    .ZN(_10183_)
  );
  AND2_X1 _44601_ (
    .A1(_10176_),
    .A2(_10183_),
    .ZN(_10184_)
  );
  AND2_X1 _44602_ (
    .A1(_22078_),
    .A2(_10184_),
    .ZN(_10185_)
  );
  INV_X1 _44603_ (
    .A(_10185_),
    .ZN(_10186_)
  );
  AND2_X1 _44604_ (
    .A1(_21400_),
    .A2(_00007_[2]),
    .ZN(_10187_)
  );
  INV_X1 _44605_ (
    .A(_10187_),
    .ZN(_10188_)
  );
  AND2_X1 _44606_ (
    .A1(_21716_),
    .A2(_22077_),
    .ZN(_10189_)
  );
  INV_X1 _44607_ (
    .A(_10189_),
    .ZN(_10190_)
  );
  AND2_X1 _44608_ (
    .A1(_10188_),
    .A2(_10190_),
    .ZN(_10191_)
  );
  AND2_X1 _44609_ (
    .A1(_22152_),
    .A2(_10191_),
    .ZN(_10192_)
  );
  INV_X1 _44610_ (
    .A(_10192_),
    .ZN(_10193_)
  );
  AND2_X1 _44611_ (
    .A1(_21589_),
    .A2(_22077_),
    .ZN(_10194_)
  );
  INV_X1 _44612_ (
    .A(_10194_),
    .ZN(_10195_)
  );
  AND2_X1 _44613_ (
    .A1(_21407_),
    .A2(_00007_[2]),
    .ZN(_10196_)
  );
  INV_X1 _44614_ (
    .A(_10196_),
    .ZN(_10197_)
  );
  AND2_X1 _44615_ (
    .A1(_00007_[0]),
    .A2(_10197_),
    .ZN(_10198_)
  );
  AND2_X1 _44616_ (
    .A1(_10195_),
    .A2(_10198_),
    .ZN(_10199_)
  );
  INV_X1 _44617_ (
    .A(_10199_),
    .ZN(_10200_)
  );
  AND2_X1 _44618_ (
    .A1(_00007_[1]),
    .A2(_10200_),
    .ZN(_10201_)
  );
  AND2_X1 _44619_ (
    .A1(_10193_),
    .A2(_10201_),
    .ZN(_10202_)
  );
  INV_X1 _44620_ (
    .A(_10202_),
    .ZN(_10203_)
  );
  AND2_X1 _44621_ (
    .A1(_10186_),
    .A2(_10203_),
    .ZN(_10204_)
  );
  AND2_X1 _44622_ (
    .A1(_22144_),
    .A2(_10204_),
    .ZN(_10205_)
  );
  INV_X1 _44623_ (
    .A(_10205_),
    .ZN(_10206_)
  );
  AND2_X1 _44624_ (
    .A1(_00007_[3]),
    .A2(_10206_),
    .ZN(_10207_)
  );
  AND2_X1 _44625_ (
    .A1(_10169_),
    .A2(_10207_),
    .ZN(_10208_)
  );
  INV_X1 _44626_ (
    .A(_10208_),
    .ZN(_10209_)
  );
  AND2_X1 _44627_ (
    .A1(_22109_),
    .A2(_10131_),
    .ZN(_10210_)
  );
  INV_X1 _44628_ (
    .A(_10210_),
    .ZN(_10211_)
  );
  AND2_X1 _44629_ (
    .A1(_10209_),
    .A2(_10211_),
    .ZN(_10212_)
  );
  AND2_X1 _44630_ (
    .A1(_05842_),
    .A2(_10212_),
    .ZN(_10213_)
  );
  INV_X1 _44631_ (
    .A(_10213_),
    .ZN(_10214_)
  );
  AND2_X1 _44632_ (
    .A1(_21230_),
    .A2(_04963_),
    .ZN(_10215_)
  );
  INV_X1 _44633_ (
    .A(_10215_),
    .ZN(_10216_)
  );
  AND2_X1 _44634_ (
    .A1(_04962_),
    .A2(_10214_),
    .ZN(_10217_)
  );
  AND2_X1 _44635_ (
    .A1(_10053_),
    .A2(_10217_),
    .ZN(_10218_)
  );
  INV_X1 _44636_ (
    .A(_10218_),
    .ZN(_10219_)
  );
  AND2_X1 _44637_ (
    .A1(_10216_),
    .A2(_10219_),
    .ZN(_00311_)
  );
  AND2_X1 _44638_ (
    .A1(\cpuregs[29] [31]),
    .A2(_00007_[2]),
    .ZN(_10220_)
  );
  INV_X1 _44639_ (
    .A(_10220_),
    .ZN(_10221_)
  );
  AND2_X1 _44640_ (
    .A1(\cpuregs[25] [31]),
    .A2(_22077_),
    .ZN(_10222_)
  );
  INV_X1 _44641_ (
    .A(_10222_),
    .ZN(_10223_)
  );
  AND2_X1 _44642_ (
    .A1(_00007_[0]),
    .A2(_10223_),
    .ZN(_10224_)
  );
  AND2_X1 _44643_ (
    .A1(_10221_),
    .A2(_10224_),
    .ZN(_10225_)
  );
  INV_X1 _44644_ (
    .A(_10225_),
    .ZN(_10226_)
  );
  AND2_X1 _44645_ (
    .A1(\cpuregs[24] [31]),
    .A2(_22077_),
    .ZN(_10227_)
  );
  INV_X1 _44646_ (
    .A(_10227_),
    .ZN(_10228_)
  );
  AND2_X1 _44647_ (
    .A1(\cpuregs[28] [31]),
    .A2(_00007_[2]),
    .ZN(_10229_)
  );
  INV_X1 _44648_ (
    .A(_10229_),
    .ZN(_10230_)
  );
  AND2_X1 _44649_ (
    .A1(_22152_),
    .A2(_10230_),
    .ZN(_10231_)
  );
  AND2_X1 _44650_ (
    .A1(_10228_),
    .A2(_10231_),
    .ZN(_10232_)
  );
  INV_X1 _44651_ (
    .A(_10232_),
    .ZN(_10233_)
  );
  AND2_X1 _44652_ (
    .A1(_22078_),
    .A2(_10233_),
    .ZN(_10234_)
  );
  AND2_X1 _44653_ (
    .A1(_10226_),
    .A2(_10234_),
    .ZN(_10235_)
  );
  INV_X1 _44654_ (
    .A(_10235_),
    .ZN(_10236_)
  );
  AND2_X1 _44655_ (
    .A1(\cpuregs[31] [31]),
    .A2(_00007_[2]),
    .ZN(_10237_)
  );
  INV_X1 _44656_ (
    .A(_10237_),
    .ZN(_10238_)
  );
  AND2_X1 _44657_ (
    .A1(\cpuregs[27] [31]),
    .A2(_22077_),
    .ZN(_10239_)
  );
  INV_X1 _44658_ (
    .A(_10239_),
    .ZN(_10240_)
  );
  AND2_X1 _44659_ (
    .A1(_00007_[0]),
    .A2(_10240_),
    .ZN(_10241_)
  );
  AND2_X1 _44660_ (
    .A1(_10238_),
    .A2(_10241_),
    .ZN(_10242_)
  );
  INV_X1 _44661_ (
    .A(_10242_),
    .ZN(_10243_)
  );
  AND2_X1 _44662_ (
    .A1(\cpuregs[26] [31]),
    .A2(_22077_),
    .ZN(_10244_)
  );
  INV_X1 _44663_ (
    .A(_10244_),
    .ZN(_10245_)
  );
  AND2_X1 _44664_ (
    .A1(\cpuregs[30] [31]),
    .A2(_00007_[2]),
    .ZN(_10246_)
  );
  INV_X1 _44665_ (
    .A(_10246_),
    .ZN(_10247_)
  );
  AND2_X1 _44666_ (
    .A1(_22152_),
    .A2(_10247_),
    .ZN(_10248_)
  );
  AND2_X1 _44667_ (
    .A1(_10245_),
    .A2(_10248_),
    .ZN(_10249_)
  );
  INV_X1 _44668_ (
    .A(_10249_),
    .ZN(_10250_)
  );
  AND2_X1 _44669_ (
    .A1(_00007_[1]),
    .A2(_10250_),
    .ZN(_10251_)
  );
  AND2_X1 _44670_ (
    .A1(_10243_),
    .A2(_10251_),
    .ZN(_10252_)
  );
  INV_X1 _44671_ (
    .A(_10252_),
    .ZN(_10253_)
  );
  AND2_X1 _44672_ (
    .A1(_10236_),
    .A2(_10253_),
    .ZN(_10254_)
  );
  INV_X1 _44673_ (
    .A(_10254_),
    .ZN(_10255_)
  );
  AND2_X1 _44674_ (
    .A1(\cpuregs[11] [31]),
    .A2(_22077_),
    .ZN(_10256_)
  );
  INV_X1 _44675_ (
    .A(_10256_),
    .ZN(_10257_)
  );
  AND2_X1 _44676_ (
    .A1(\cpuregs[15] [31]),
    .A2(_00007_[2]),
    .ZN(_10258_)
  );
  INV_X1 _44677_ (
    .A(_10258_),
    .ZN(_10259_)
  );
  AND2_X1 _44678_ (
    .A1(_10257_),
    .A2(_10259_),
    .ZN(_10260_)
  );
  INV_X1 _44679_ (
    .A(_10260_),
    .ZN(_10261_)
  );
  AND2_X1 _44680_ (
    .A1(_00007_[0]),
    .A2(_10261_),
    .ZN(_10262_)
  );
  INV_X1 _44681_ (
    .A(_10262_),
    .ZN(_10263_)
  );
  AND2_X1 _44682_ (
    .A1(\cpuregs[14] [31]),
    .A2(_00007_[2]),
    .ZN(_10264_)
  );
  INV_X1 _44683_ (
    .A(_10264_),
    .ZN(_10265_)
  );
  AND2_X1 _44684_ (
    .A1(\cpuregs[10] [31]),
    .A2(_22077_),
    .ZN(_10266_)
  );
  INV_X1 _44685_ (
    .A(_10266_),
    .ZN(_10267_)
  );
  AND2_X1 _44686_ (
    .A1(_10265_),
    .A2(_10267_),
    .ZN(_10268_)
  );
  INV_X1 _44687_ (
    .A(_10268_),
    .ZN(_10269_)
  );
  AND2_X1 _44688_ (
    .A1(_22152_),
    .A2(_10269_),
    .ZN(_10270_)
  );
  INV_X1 _44689_ (
    .A(_10270_),
    .ZN(_10271_)
  );
  AND2_X1 _44690_ (
    .A1(_10263_),
    .A2(_10271_),
    .ZN(_10272_)
  );
  AND2_X1 _44691_ (
    .A1(\cpuregs[9] [31]),
    .A2(_22077_),
    .ZN(_10273_)
  );
  INV_X1 _44692_ (
    .A(_10273_),
    .ZN(_10274_)
  );
  AND2_X1 _44693_ (
    .A1(\cpuregs[13] [31]),
    .A2(_00007_[2]),
    .ZN(_10275_)
  );
  INV_X1 _44694_ (
    .A(_10275_),
    .ZN(_10276_)
  );
  AND2_X1 _44695_ (
    .A1(_10274_),
    .A2(_10276_),
    .ZN(_10277_)
  );
  INV_X1 _44696_ (
    .A(_10277_),
    .ZN(_10278_)
  );
  AND2_X1 _44697_ (
    .A1(_00007_[0]),
    .A2(_10278_),
    .ZN(_10279_)
  );
  INV_X1 _44698_ (
    .A(_10279_),
    .ZN(_10280_)
  );
  AND2_X1 _44699_ (
    .A1(\cpuregs[12] [31]),
    .A2(_00007_[2]),
    .ZN(_10281_)
  );
  INV_X1 _44700_ (
    .A(_10281_),
    .ZN(_10282_)
  );
  AND2_X1 _44701_ (
    .A1(\cpuregs[8] [31]),
    .A2(_22077_),
    .ZN(_10283_)
  );
  INV_X1 _44702_ (
    .A(_10283_),
    .ZN(_10284_)
  );
  AND2_X1 _44703_ (
    .A1(_10282_),
    .A2(_10284_),
    .ZN(_10285_)
  );
  INV_X1 _44704_ (
    .A(_10285_),
    .ZN(_10286_)
  );
  AND2_X1 _44705_ (
    .A1(_22152_),
    .A2(_10286_),
    .ZN(_10287_)
  );
  INV_X1 _44706_ (
    .A(_10287_),
    .ZN(_10288_)
  );
  AND2_X1 _44707_ (
    .A1(_10280_),
    .A2(_10288_),
    .ZN(_10289_)
  );
  AND2_X1 _44708_ (
    .A1(_21369_),
    .A2(_22077_),
    .ZN(_10290_)
  );
  INV_X1 _44709_ (
    .A(_10290_),
    .ZN(_10291_)
  );
  AND2_X1 _44710_ (
    .A1(_21365_),
    .A2(_00007_[2]),
    .ZN(_10292_)
  );
  INV_X1 _44711_ (
    .A(_10292_),
    .ZN(_10293_)
  );
  AND2_X1 _44712_ (
    .A1(_10291_),
    .A2(_10293_),
    .ZN(_10294_)
  );
  AND2_X1 _44713_ (
    .A1(_21368_),
    .A2(_22077_),
    .ZN(_10295_)
  );
  INV_X1 _44714_ (
    .A(_10295_),
    .ZN(_10296_)
  );
  AND2_X1 _44715_ (
    .A1(_21364_),
    .A2(_00007_[2]),
    .ZN(_10297_)
  );
  INV_X1 _44716_ (
    .A(_10297_),
    .ZN(_10298_)
  );
  AND2_X1 _44717_ (
    .A1(_00007_[0]),
    .A2(_10298_),
    .ZN(_10299_)
  );
  AND2_X1 _44718_ (
    .A1(_10296_),
    .A2(_10299_),
    .ZN(_10300_)
  );
  INV_X1 _44719_ (
    .A(_10300_),
    .ZN(_10301_)
  );
  AND2_X1 _44720_ (
    .A1(_22152_),
    .A2(_10294_),
    .ZN(_10302_)
  );
  INV_X1 _44721_ (
    .A(_10302_),
    .ZN(_10303_)
  );
  AND2_X1 _44722_ (
    .A1(_10301_),
    .A2(_10303_),
    .ZN(_10304_)
  );
  AND2_X1 _44723_ (
    .A1(_21367_),
    .A2(_22077_),
    .ZN(_10305_)
  );
  INV_X1 _44724_ (
    .A(_10305_),
    .ZN(_10306_)
  );
  AND2_X1 _44725_ (
    .A1(_21363_),
    .A2(_00007_[2]),
    .ZN(_10307_)
  );
  INV_X1 _44726_ (
    .A(_10307_),
    .ZN(_10308_)
  );
  AND2_X1 _44727_ (
    .A1(_21362_),
    .A2(_00007_[2]),
    .ZN(_10309_)
  );
  INV_X1 _44728_ (
    .A(_10309_),
    .ZN(_10310_)
  );
  AND2_X1 _44729_ (
    .A1(_21366_),
    .A2(_22077_),
    .ZN(_10311_)
  );
  INV_X1 _44730_ (
    .A(_10311_),
    .ZN(_10312_)
  );
  AND2_X1 _44731_ (
    .A1(_22152_),
    .A2(_10308_),
    .ZN(_10313_)
  );
  AND2_X1 _44732_ (
    .A1(_10306_),
    .A2(_10313_),
    .ZN(_10314_)
  );
  INV_X1 _44733_ (
    .A(_10314_),
    .ZN(_10315_)
  );
  AND2_X1 _44734_ (
    .A1(_00007_[0]),
    .A2(_10310_),
    .ZN(_10316_)
  );
  AND2_X1 _44735_ (
    .A1(_10312_),
    .A2(_10316_),
    .ZN(_10317_)
  );
  INV_X1 _44736_ (
    .A(_10317_),
    .ZN(_10318_)
  );
  AND2_X1 _44737_ (
    .A1(_10315_),
    .A2(_10318_),
    .ZN(_10319_)
  );
  AND2_X1 _44738_ (
    .A1(_00007_[1]),
    .A2(_10319_),
    .ZN(_10320_)
  );
  INV_X1 _44739_ (
    .A(_10320_),
    .ZN(_10321_)
  );
  AND2_X1 _44740_ (
    .A1(_22078_),
    .A2(_10304_),
    .ZN(_10322_)
  );
  INV_X1 _44741_ (
    .A(_10322_),
    .ZN(_10323_)
  );
  AND2_X1 _44742_ (
    .A1(_10321_),
    .A2(_10323_),
    .ZN(_10324_)
  );
  AND2_X1 _44743_ (
    .A1(_21361_),
    .A2(_22077_),
    .ZN(_10325_)
  );
  INV_X1 _44744_ (
    .A(_10325_),
    .ZN(_10326_)
  );
  AND2_X1 _44745_ (
    .A1(_21360_),
    .A2(_00007_[2]),
    .ZN(_10327_)
  );
  INV_X1 _44746_ (
    .A(_10327_),
    .ZN(_10328_)
  );
  AND2_X1 _44747_ (
    .A1(_22152_),
    .A2(_10328_),
    .ZN(_10329_)
  );
  AND2_X1 _44748_ (
    .A1(_10326_),
    .A2(_10329_),
    .ZN(_10330_)
  );
  INV_X1 _44749_ (
    .A(_10330_),
    .ZN(_10331_)
  );
  AND2_X1 _44750_ (
    .A1(\cpuregs[7] [31]),
    .A2(_00007_[2]),
    .ZN(_10332_)
  );
  INV_X1 _44751_ (
    .A(_10332_),
    .ZN(_10333_)
  );
  AND2_X1 _44752_ (
    .A1(\cpuregs[3] [31]),
    .A2(_22077_),
    .ZN(_10334_)
  );
  INV_X1 _44753_ (
    .A(_10334_),
    .ZN(_10335_)
  );
  AND2_X1 _44754_ (
    .A1(_10333_),
    .A2(_10335_),
    .ZN(_10336_)
  );
  INV_X1 _44755_ (
    .A(_10336_),
    .ZN(_10337_)
  );
  AND2_X1 _44756_ (
    .A1(_00007_[0]),
    .A2(_10337_),
    .ZN(_10338_)
  );
  INV_X1 _44757_ (
    .A(_10338_),
    .ZN(_10339_)
  );
  AND2_X1 _44758_ (
    .A1(_10331_),
    .A2(_10339_),
    .ZN(_10340_)
  );
  AND2_X1 _44759_ (
    .A1(\cpuregs[1] [31]),
    .A2(_22077_),
    .ZN(_10341_)
  );
  INV_X1 _44760_ (
    .A(_10341_),
    .ZN(_10342_)
  );
  AND2_X1 _44761_ (
    .A1(\cpuregs[5] [31]),
    .A2(_00007_[2]),
    .ZN(_10343_)
  );
  INV_X1 _44762_ (
    .A(_10343_),
    .ZN(_10344_)
  );
  AND2_X1 _44763_ (
    .A1(_10342_),
    .A2(_10344_),
    .ZN(_10345_)
  );
  INV_X1 _44764_ (
    .A(_10345_),
    .ZN(_10346_)
  );
  AND2_X1 _44765_ (
    .A1(_00007_[0]),
    .A2(_10346_),
    .ZN(_10347_)
  );
  INV_X1 _44766_ (
    .A(_10347_),
    .ZN(_10348_)
  );
  AND2_X1 _44767_ (
    .A1(\cpuregs[4] [31]),
    .A2(_00007_[2]),
    .ZN(_10349_)
  );
  INV_X1 _44768_ (
    .A(_10349_),
    .ZN(_10350_)
  );
  AND2_X1 _44769_ (
    .A1(\cpuregs[0] [31]),
    .A2(_22077_),
    .ZN(_10351_)
  );
  INV_X1 _44770_ (
    .A(_10351_),
    .ZN(_10352_)
  );
  AND2_X1 _44771_ (
    .A1(_10350_),
    .A2(_10352_),
    .ZN(_10353_)
  );
  INV_X1 _44772_ (
    .A(_10353_),
    .ZN(_10354_)
  );
  AND2_X1 _44773_ (
    .A1(_22152_),
    .A2(_10354_),
    .ZN(_10355_)
  );
  INV_X1 _44774_ (
    .A(_10355_),
    .ZN(_10356_)
  );
  AND2_X1 _44775_ (
    .A1(_10348_),
    .A2(_10356_),
    .ZN(_10357_)
  );
  AND2_X1 _44776_ (
    .A1(_00007_[1]),
    .A2(_10340_),
    .ZN(_10358_)
  );
  INV_X1 _44777_ (
    .A(_10358_),
    .ZN(_10359_)
  );
  AND2_X1 _44778_ (
    .A1(_22078_),
    .A2(_10357_),
    .ZN(_10360_)
  );
  INV_X1 _44779_ (
    .A(_10360_),
    .ZN(_10361_)
  );
  AND2_X1 _44780_ (
    .A1(_10359_),
    .A2(_10361_),
    .ZN(_10362_)
  );
  AND2_X1 _44781_ (
    .A1(_22109_),
    .A2(_10324_),
    .ZN(_10363_)
  );
  INV_X1 _44782_ (
    .A(_10363_),
    .ZN(_10364_)
  );
  AND2_X1 _44783_ (
    .A1(_00007_[3]),
    .A2(_10255_),
    .ZN(_10365_)
  );
  INV_X1 _44784_ (
    .A(_10365_),
    .ZN(_10366_)
  );
  AND2_X1 _44785_ (
    .A1(_00007_[4]),
    .A2(_10366_),
    .ZN(_10367_)
  );
  AND2_X1 _44786_ (
    .A1(_10364_),
    .A2(_10367_),
    .ZN(_10368_)
  );
  INV_X1 _44787_ (
    .A(_10368_),
    .ZN(_10369_)
  );
  AND2_X1 _44788_ (
    .A1(_00007_[1]),
    .A2(_10272_),
    .ZN(_10370_)
  );
  INV_X1 _44789_ (
    .A(_10370_),
    .ZN(_10371_)
  );
  AND2_X1 _44790_ (
    .A1(_22078_),
    .A2(_10289_),
    .ZN(_10372_)
  );
  INV_X1 _44791_ (
    .A(_10372_),
    .ZN(_10373_)
  );
  AND2_X1 _44792_ (
    .A1(_00007_[3]),
    .A2(_10373_),
    .ZN(_10374_)
  );
  AND2_X1 _44793_ (
    .A1(_10371_),
    .A2(_10374_),
    .ZN(_10375_)
  );
  INV_X1 _44794_ (
    .A(_10375_),
    .ZN(_10376_)
  );
  AND2_X1 _44795_ (
    .A1(_22109_),
    .A2(_10362_),
    .ZN(_10377_)
  );
  INV_X1 _44796_ (
    .A(_10377_),
    .ZN(_10378_)
  );
  AND2_X1 _44797_ (
    .A1(_10376_),
    .A2(_10378_),
    .ZN(_10379_)
  );
  AND2_X1 _44798_ (
    .A1(_22144_),
    .A2(_10379_),
    .ZN(_10380_)
  );
  INV_X1 _44799_ (
    .A(_10380_),
    .ZN(_10381_)
  );
  AND2_X1 _44800_ (
    .A1(_10369_),
    .A2(_10381_),
    .ZN(_10382_)
  );
  AND2_X1 _44801_ (
    .A1(_05842_),
    .A2(_10382_),
    .ZN(_10383_)
  );
  INV_X1 _44802_ (
    .A(_10383_),
    .ZN(_10384_)
  );
  AND2_X1 _44803_ (
    .A1(decoded_imm[31]),
    .A2(_04966_),
    .ZN(_10385_)
  );
  INV_X1 _44804_ (
    .A(_10385_),
    .ZN(_10386_)
  );
  AND2_X1 _44805_ (
    .A1(_21231_),
    .A2(_04963_),
    .ZN(_10387_)
  );
  INV_X1 _44806_ (
    .A(_10387_),
    .ZN(_10388_)
  );
  AND2_X1 _44807_ (
    .A1(_04962_),
    .A2(_10386_),
    .ZN(_10389_)
  );
  AND2_X1 _44808_ (
    .A1(_10384_),
    .A2(_10389_),
    .ZN(_10390_)
  );
  INV_X1 _44809_ (
    .A(_10390_),
    .ZN(_10391_)
  );
  AND2_X1 _44810_ (
    .A1(_10388_),
    .A2(_10391_),
    .ZN(_00312_)
  );
  AND2_X1 _44811_ (
    .A1(mem_rdata[7]),
    .A2(_22307_),
    .ZN(_10392_)
  );
  INV_X1 _44812_ (
    .A(_10392_),
    .ZN(_10393_)
  );
  AND2_X1 _44813_ (
    .A1(mem_rdata_q[7]),
    .A2(_22308_),
    .ZN(_10394_)
  );
  INV_X1 _44814_ (
    .A(_10394_),
    .ZN(_10395_)
  );
  AND2_X1 _44815_ (
    .A1(_10393_),
    .A2(_10395_),
    .ZN(_10396_)
  );
  INV_X1 _44816_ (
    .A(_10396_),
    .ZN(_00313_)
  );
  AND2_X1 _44817_ (
    .A1(mem_rdata[8]),
    .A2(_22307_),
    .ZN(_10397_)
  );
  INV_X1 _44818_ (
    .A(_10397_),
    .ZN(_10398_)
  );
  AND2_X1 _44819_ (
    .A1(mem_rdata_q[8]),
    .A2(_22308_),
    .ZN(_10399_)
  );
  INV_X1 _44820_ (
    .A(_10399_),
    .ZN(_10400_)
  );
  AND2_X1 _44821_ (
    .A1(_10398_),
    .A2(_10400_),
    .ZN(_10401_)
  );
  INV_X1 _44822_ (
    .A(_10401_),
    .ZN(_00314_)
  );
  AND2_X1 _44823_ (
    .A1(mem_rdata[9]),
    .A2(_22307_),
    .ZN(_10402_)
  );
  INV_X1 _44824_ (
    .A(_10402_),
    .ZN(_10403_)
  );
  AND2_X1 _44825_ (
    .A1(mem_rdata_q[9]),
    .A2(_22308_),
    .ZN(_10404_)
  );
  INV_X1 _44826_ (
    .A(_10404_),
    .ZN(_10405_)
  );
  AND2_X1 _44827_ (
    .A1(_10403_),
    .A2(_10405_),
    .ZN(_10406_)
  );
  INV_X1 _44828_ (
    .A(_10406_),
    .ZN(_00315_)
  );
  AND2_X1 _44829_ (
    .A1(mem_rdata[10]),
    .A2(_22307_),
    .ZN(_10407_)
  );
  INV_X1 _44830_ (
    .A(_10407_),
    .ZN(_10408_)
  );
  AND2_X1 _44831_ (
    .A1(mem_rdata_q[10]),
    .A2(_22308_),
    .ZN(_10409_)
  );
  INV_X1 _44832_ (
    .A(_10409_),
    .ZN(_10410_)
  );
  AND2_X1 _44833_ (
    .A1(_10408_),
    .A2(_10410_),
    .ZN(_10411_)
  );
  INV_X1 _44834_ (
    .A(_10411_),
    .ZN(_00316_)
  );
  AND2_X1 _44835_ (
    .A1(mem_rdata[11]),
    .A2(_22307_),
    .ZN(_10412_)
  );
  INV_X1 _44836_ (
    .A(_10412_),
    .ZN(_10413_)
  );
  AND2_X1 _44837_ (
    .A1(mem_rdata_q[11]),
    .A2(_22308_),
    .ZN(_10414_)
  );
  INV_X1 _44838_ (
    .A(_10414_),
    .ZN(_10415_)
  );
  AND2_X1 _44839_ (
    .A1(_10413_),
    .A2(_10415_),
    .ZN(_10416_)
  );
  INV_X1 _44840_ (
    .A(_10416_),
    .ZN(_00317_)
  );
  AND2_X1 _44841_ (
    .A1(mem_rdata[12]),
    .A2(_22307_),
    .ZN(_10417_)
  );
  INV_X1 _44842_ (
    .A(_10417_),
    .ZN(_10418_)
  );
  AND2_X1 _44843_ (
    .A1(mem_rdata_q[12]),
    .A2(_22308_),
    .ZN(_10419_)
  );
  INV_X1 _44844_ (
    .A(_10419_),
    .ZN(_10420_)
  );
  AND2_X1 _44845_ (
    .A1(_10418_),
    .A2(_10420_),
    .ZN(_10421_)
  );
  INV_X1 _44846_ (
    .A(_10421_),
    .ZN(_00318_)
  );
  AND2_X1 _44847_ (
    .A1(mem_rdata[13]),
    .A2(_22307_),
    .ZN(_10422_)
  );
  INV_X1 _44848_ (
    .A(_10422_),
    .ZN(_10423_)
  );
  AND2_X1 _44849_ (
    .A1(mem_rdata_q[13]),
    .A2(_22308_),
    .ZN(_10424_)
  );
  INV_X1 _44850_ (
    .A(_10424_),
    .ZN(_10425_)
  );
  AND2_X1 _44851_ (
    .A1(_10423_),
    .A2(_10425_),
    .ZN(_10426_)
  );
  INV_X1 _44852_ (
    .A(_10426_),
    .ZN(_00319_)
  );
  AND2_X1 _44853_ (
    .A1(mem_rdata[14]),
    .A2(_22307_),
    .ZN(_10427_)
  );
  INV_X1 _44854_ (
    .A(_10427_),
    .ZN(_10428_)
  );
  AND2_X1 _44855_ (
    .A1(mem_rdata_q[14]),
    .A2(_22308_),
    .ZN(_10429_)
  );
  INV_X1 _44856_ (
    .A(_10429_),
    .ZN(_10430_)
  );
  AND2_X1 _44857_ (
    .A1(_10428_),
    .A2(_10430_),
    .ZN(_10431_)
  );
  INV_X1 _44858_ (
    .A(_10431_),
    .ZN(_00320_)
  );
  AND2_X1 _44859_ (
    .A1(mem_rdata[15]),
    .A2(_22307_),
    .ZN(_10432_)
  );
  INV_X1 _44860_ (
    .A(_10432_),
    .ZN(_10433_)
  );
  AND2_X1 _44861_ (
    .A1(mem_rdata_q[15]),
    .A2(_22308_),
    .ZN(_10434_)
  );
  INV_X1 _44862_ (
    .A(_10434_),
    .ZN(_10435_)
  );
  AND2_X1 _44863_ (
    .A1(_10433_),
    .A2(_10435_),
    .ZN(_10436_)
  );
  INV_X1 _44864_ (
    .A(_10436_),
    .ZN(_00321_)
  );
  AND2_X1 _44865_ (
    .A1(mem_rdata[16]),
    .A2(_22307_),
    .ZN(_10437_)
  );
  INV_X1 _44866_ (
    .A(_10437_),
    .ZN(_10438_)
  );
  AND2_X1 _44867_ (
    .A1(mem_rdata_q[16]),
    .A2(_22308_),
    .ZN(_10439_)
  );
  INV_X1 _44868_ (
    .A(_10439_),
    .ZN(_10440_)
  );
  AND2_X1 _44869_ (
    .A1(_10438_),
    .A2(_10440_),
    .ZN(_10441_)
  );
  INV_X1 _44870_ (
    .A(_10441_),
    .ZN(_00322_)
  );
  AND2_X1 _44871_ (
    .A1(mem_rdata[17]),
    .A2(_22307_),
    .ZN(_10442_)
  );
  INV_X1 _44872_ (
    .A(_10442_),
    .ZN(_10443_)
  );
  AND2_X1 _44873_ (
    .A1(mem_rdata_q[17]),
    .A2(_22308_),
    .ZN(_10444_)
  );
  INV_X1 _44874_ (
    .A(_10444_),
    .ZN(_10445_)
  );
  AND2_X1 _44875_ (
    .A1(_10443_),
    .A2(_10445_),
    .ZN(_10446_)
  );
  INV_X1 _44876_ (
    .A(_10446_),
    .ZN(_00323_)
  );
  AND2_X1 _44877_ (
    .A1(mem_rdata[18]),
    .A2(_22307_),
    .ZN(_10447_)
  );
  INV_X1 _44878_ (
    .A(_10447_),
    .ZN(_10448_)
  );
  AND2_X1 _44879_ (
    .A1(mem_rdata_q[18]),
    .A2(_22308_),
    .ZN(_10449_)
  );
  INV_X1 _44880_ (
    .A(_10449_),
    .ZN(_10450_)
  );
  AND2_X1 _44881_ (
    .A1(_10448_),
    .A2(_10450_),
    .ZN(_10451_)
  );
  INV_X1 _44882_ (
    .A(_10451_),
    .ZN(_00324_)
  );
  AND2_X1 _44883_ (
    .A1(mem_rdata[19]),
    .A2(_22307_),
    .ZN(_10452_)
  );
  INV_X1 _44884_ (
    .A(_10452_),
    .ZN(_10453_)
  );
  AND2_X1 _44885_ (
    .A1(mem_rdata_q[19]),
    .A2(_22308_),
    .ZN(_10454_)
  );
  INV_X1 _44886_ (
    .A(_10454_),
    .ZN(_10455_)
  );
  AND2_X1 _44887_ (
    .A1(_10453_),
    .A2(_10455_),
    .ZN(_10456_)
  );
  INV_X1 _44888_ (
    .A(_10456_),
    .ZN(_00325_)
  );
  AND2_X1 _44889_ (
    .A1(mem_rdata[20]),
    .A2(_22307_),
    .ZN(_10457_)
  );
  INV_X1 _44890_ (
    .A(_10457_),
    .ZN(_10458_)
  );
  AND2_X1 _44891_ (
    .A1(mem_rdata_q[20]),
    .A2(_22308_),
    .ZN(_10459_)
  );
  INV_X1 _44892_ (
    .A(_10459_),
    .ZN(_10460_)
  );
  AND2_X1 _44893_ (
    .A1(_10458_),
    .A2(_10460_),
    .ZN(_10461_)
  );
  INV_X1 _44894_ (
    .A(_10461_),
    .ZN(_00326_)
  );
  AND2_X1 _44895_ (
    .A1(mem_rdata[21]),
    .A2(_22307_),
    .ZN(_10462_)
  );
  INV_X1 _44896_ (
    .A(_10462_),
    .ZN(_10463_)
  );
  AND2_X1 _44897_ (
    .A1(mem_rdata_q[21]),
    .A2(_22308_),
    .ZN(_10464_)
  );
  INV_X1 _44898_ (
    .A(_10464_),
    .ZN(_10465_)
  );
  AND2_X1 _44899_ (
    .A1(_10463_),
    .A2(_10465_),
    .ZN(_10466_)
  );
  INV_X1 _44900_ (
    .A(_10466_),
    .ZN(_00327_)
  );
  AND2_X1 _44901_ (
    .A1(mem_rdata[22]),
    .A2(_22307_),
    .ZN(_10467_)
  );
  INV_X1 _44902_ (
    .A(_10467_),
    .ZN(_10468_)
  );
  AND2_X1 _44903_ (
    .A1(mem_rdata_q[22]),
    .A2(_22308_),
    .ZN(_10469_)
  );
  INV_X1 _44904_ (
    .A(_10469_),
    .ZN(_10470_)
  );
  AND2_X1 _44905_ (
    .A1(_10468_),
    .A2(_10470_),
    .ZN(_10471_)
  );
  INV_X1 _44906_ (
    .A(_10471_),
    .ZN(_00328_)
  );
  AND2_X1 _44907_ (
    .A1(mem_rdata[23]),
    .A2(_22307_),
    .ZN(_10472_)
  );
  INV_X1 _44908_ (
    .A(_10472_),
    .ZN(_10473_)
  );
  AND2_X1 _44909_ (
    .A1(mem_rdata_q[23]),
    .A2(_22308_),
    .ZN(_10474_)
  );
  INV_X1 _44910_ (
    .A(_10474_),
    .ZN(_10475_)
  );
  AND2_X1 _44911_ (
    .A1(_10473_),
    .A2(_10475_),
    .ZN(_10476_)
  );
  INV_X1 _44912_ (
    .A(_10476_),
    .ZN(_00329_)
  );
  AND2_X1 _44913_ (
    .A1(mem_rdata[24]),
    .A2(_22307_),
    .ZN(_10477_)
  );
  INV_X1 _44914_ (
    .A(_10477_),
    .ZN(_10478_)
  );
  AND2_X1 _44915_ (
    .A1(mem_rdata_q[24]),
    .A2(_22308_),
    .ZN(_10479_)
  );
  INV_X1 _44916_ (
    .A(_10479_),
    .ZN(_10480_)
  );
  AND2_X1 _44917_ (
    .A1(_10478_),
    .A2(_10480_),
    .ZN(_10481_)
  );
  INV_X1 _44918_ (
    .A(_10481_),
    .ZN(_00330_)
  );
  AND2_X1 _44919_ (
    .A1(mem_rdata[25]),
    .A2(_22307_),
    .ZN(_10482_)
  );
  INV_X1 _44920_ (
    .A(_10482_),
    .ZN(_10483_)
  );
  AND2_X1 _44921_ (
    .A1(mem_rdata_q[25]),
    .A2(_22308_),
    .ZN(_10484_)
  );
  INV_X1 _44922_ (
    .A(_10484_),
    .ZN(_10485_)
  );
  AND2_X1 _44923_ (
    .A1(_10483_),
    .A2(_10485_),
    .ZN(_10486_)
  );
  INV_X1 _44924_ (
    .A(_10486_),
    .ZN(_00331_)
  );
  AND2_X1 _44925_ (
    .A1(mem_rdata[26]),
    .A2(_22307_),
    .ZN(_10487_)
  );
  INV_X1 _44926_ (
    .A(_10487_),
    .ZN(_10488_)
  );
  AND2_X1 _44927_ (
    .A1(mem_rdata_q[26]),
    .A2(_22308_),
    .ZN(_10489_)
  );
  INV_X1 _44928_ (
    .A(_10489_),
    .ZN(_10490_)
  );
  AND2_X1 _44929_ (
    .A1(_10488_),
    .A2(_10490_),
    .ZN(_10491_)
  );
  INV_X1 _44930_ (
    .A(_10491_),
    .ZN(_00332_)
  );
  AND2_X1 _44931_ (
    .A1(mem_rdata[27]),
    .A2(_22307_),
    .ZN(_10492_)
  );
  INV_X1 _44932_ (
    .A(_10492_),
    .ZN(_10493_)
  );
  AND2_X1 _44933_ (
    .A1(mem_rdata_q[27]),
    .A2(_22308_),
    .ZN(_10494_)
  );
  INV_X1 _44934_ (
    .A(_10494_),
    .ZN(_10495_)
  );
  AND2_X1 _44935_ (
    .A1(_10493_),
    .A2(_10495_),
    .ZN(_10496_)
  );
  INV_X1 _44936_ (
    .A(_10496_),
    .ZN(_00333_)
  );
  AND2_X1 _44937_ (
    .A1(mem_rdata[28]),
    .A2(_22307_),
    .ZN(_10497_)
  );
  INV_X1 _44938_ (
    .A(_10497_),
    .ZN(_10498_)
  );
  AND2_X1 _44939_ (
    .A1(mem_rdata_q[28]),
    .A2(_22308_),
    .ZN(_10499_)
  );
  INV_X1 _44940_ (
    .A(_10499_),
    .ZN(_10500_)
  );
  AND2_X1 _44941_ (
    .A1(_10498_),
    .A2(_10500_),
    .ZN(_10501_)
  );
  INV_X1 _44942_ (
    .A(_10501_),
    .ZN(_00334_)
  );
  AND2_X1 _44943_ (
    .A1(mem_rdata[29]),
    .A2(_22307_),
    .ZN(_10502_)
  );
  INV_X1 _44944_ (
    .A(_10502_),
    .ZN(_10503_)
  );
  AND2_X1 _44945_ (
    .A1(mem_rdata_q[29]),
    .A2(_22308_),
    .ZN(_10504_)
  );
  INV_X1 _44946_ (
    .A(_10504_),
    .ZN(_10505_)
  );
  AND2_X1 _44947_ (
    .A1(_10503_),
    .A2(_10505_),
    .ZN(_10506_)
  );
  INV_X1 _44948_ (
    .A(_10506_),
    .ZN(_00335_)
  );
  AND2_X1 _44949_ (
    .A1(mem_rdata[30]),
    .A2(_22307_),
    .ZN(_10507_)
  );
  INV_X1 _44950_ (
    .A(_10507_),
    .ZN(_10508_)
  );
  AND2_X1 _44951_ (
    .A1(mem_rdata_q[30]),
    .A2(_22308_),
    .ZN(_10509_)
  );
  INV_X1 _44952_ (
    .A(_10509_),
    .ZN(_10510_)
  );
  AND2_X1 _44953_ (
    .A1(_10508_),
    .A2(_10510_),
    .ZN(_10511_)
  );
  INV_X1 _44954_ (
    .A(_10511_),
    .ZN(_00336_)
  );
  AND2_X1 _44955_ (
    .A1(mem_rdata[31]),
    .A2(_22307_),
    .ZN(_10512_)
  );
  INV_X1 _44956_ (
    .A(_10512_),
    .ZN(_10513_)
  );
  AND2_X1 _44957_ (
    .A1(mem_rdata_q[31]),
    .A2(_22308_),
    .ZN(_10514_)
  );
  INV_X1 _44958_ (
    .A(_10514_),
    .ZN(_10515_)
  );
  AND2_X1 _44959_ (
    .A1(_10513_),
    .A2(_10515_),
    .ZN(_10516_)
  );
  INV_X1 _44960_ (
    .A(_10516_),
    .ZN(_00337_)
  );
  AND2_X1 _44961_ (
    .A1(_00029_),
    .A2(_02469_),
    .ZN(_10517_)
  );
  INV_X1 _44962_ (
    .A(_10517_),
    .ZN(_10518_)
  );
  AND2_X1 _44963_ (
    .A1(_21072_),
    .A2(_10517_),
    .ZN(_10519_)
  );
  INV_X1 _44964_ (
    .A(_10519_),
    .ZN(_10520_)
  );
  AND2_X1 _44965_ (
    .A1(resetn),
    .A2(_22316_),
    .ZN(_10521_)
  );
  AND2_X1 _44966_ (
    .A1(_21071_),
    .A2(_10518_),
    .ZN(_10522_)
  );
  INV_X1 _44967_ (
    .A(_10522_),
    .ZN(_10523_)
  );
  AND2_X1 _44968_ (
    .A1(_10520_),
    .A2(_10521_),
    .ZN(_10524_)
  );
  AND2_X1 _44969_ (
    .A1(_10523_),
    .A2(_10524_),
    .ZN(_00338_)
  );
  AND2_X1 _44970_ (
    .A1(reg_op1[31]),
    .A2(_29151_[31]),
    .ZN(_10525_)
  );
  INV_X1 _44971_ (
    .A(_10525_),
    .ZN(_10526_)
  );
  AND2_X1 _44972_ (
    .A1(_21199_),
    .A2(_22249_),
    .ZN(_10527_)
  );
  INV_X1 _44973_ (
    .A(_10527_),
    .ZN(_10528_)
  );
  AND2_X1 _44974_ (
    .A1(_10526_),
    .A2(_10528_),
    .ZN(_10529_)
  );
  INV_X1 _44975_ (
    .A(_10529_),
    .ZN(_10530_)
  );
  AND2_X1 _44976_ (
    .A1(reg_op1[30]),
    .A2(_29151_[30]),
    .ZN(_10531_)
  );
  INV_X1 _44977_ (
    .A(_10531_),
    .ZN(_10532_)
  );
  AND2_X1 _44978_ (
    .A1(_21197_),
    .A2(_22231_),
    .ZN(_10533_)
  );
  INV_X1 _44979_ (
    .A(_10533_),
    .ZN(_10534_)
  );
  AND2_X1 _44980_ (
    .A1(_10532_),
    .A2(_10534_),
    .ZN(_10535_)
  );
  INV_X1 _44981_ (
    .A(_10535_),
    .ZN(_10536_)
  );
  AND2_X1 _44982_ (
    .A1(_21196_),
    .A2(_22219_),
    .ZN(_10537_)
  );
  INV_X1 _44983_ (
    .A(_10537_),
    .ZN(_10538_)
  );
  AND2_X1 _44984_ (
    .A1(reg_op1[28]),
    .A2(_29151_[28]),
    .ZN(_10539_)
  );
  INV_X1 _44985_ (
    .A(_10539_),
    .ZN(_10540_)
  );
  AND2_X1 _44986_ (
    .A1(_21195_),
    .A2(_22218_),
    .ZN(_10541_)
  );
  INV_X1 _44987_ (
    .A(_10541_),
    .ZN(_10542_)
  );
  AND2_X1 _44988_ (
    .A1(_10540_),
    .A2(_10542_),
    .ZN(_10543_)
  );
  INV_X1 _44989_ (
    .A(_10543_),
    .ZN(_10544_)
  );
  AND2_X1 _44990_ (
    .A1(reg_op1[27]),
    .A2(_29151_[27]),
    .ZN(_10545_)
  );
  INV_X1 _44991_ (
    .A(_10545_),
    .ZN(_10546_)
  );
  AND2_X1 _44992_ (
    .A1(_21194_),
    .A2(_22241_),
    .ZN(_10547_)
  );
  INV_X1 _44993_ (
    .A(_10547_),
    .ZN(_10548_)
  );
  AND2_X1 _44994_ (
    .A1(reg_op1[26]),
    .A2(_29151_[26]),
    .ZN(_10549_)
  );
  INV_X1 _44995_ (
    .A(_10549_),
    .ZN(_10550_)
  );
  AND2_X1 _44996_ (
    .A1(_21193_),
    .A2(_22248_),
    .ZN(_10551_)
  );
  INV_X1 _44997_ (
    .A(_10551_),
    .ZN(_10552_)
  );
  AND2_X1 _44998_ (
    .A1(_10550_),
    .A2(_10552_),
    .ZN(_10553_)
  );
  INV_X1 _44999_ (
    .A(_10553_),
    .ZN(_10554_)
  );
  AND2_X1 _45000_ (
    .A1(reg_op1[25]),
    .A2(_29151_[25]),
    .ZN(_10555_)
  );
  INV_X1 _45001_ (
    .A(_10555_),
    .ZN(_10556_)
  );
  AND2_X1 _45002_ (
    .A1(_21192_),
    .A2(_22230_),
    .ZN(_10557_)
  );
  INV_X1 _45003_ (
    .A(_10557_),
    .ZN(_10558_)
  );
  AND2_X1 _45004_ (
    .A1(reg_op1[24]),
    .A2(_29151_[24]),
    .ZN(_10559_)
  );
  INV_X1 _45005_ (
    .A(_10559_),
    .ZN(_10560_)
  );
  AND2_X1 _45006_ (
    .A1(_21191_),
    .A2(_22240_),
    .ZN(_10561_)
  );
  INV_X1 _45007_ (
    .A(_10561_),
    .ZN(_10562_)
  );
  AND2_X1 _45008_ (
    .A1(_10560_),
    .A2(_10562_),
    .ZN(_10563_)
  );
  INV_X1 _45009_ (
    .A(_10563_),
    .ZN(_10564_)
  );
  AND2_X1 _45010_ (
    .A1(reg_op1[23]),
    .A2(_29151_[23]),
    .ZN(_10565_)
  );
  INV_X1 _45011_ (
    .A(_10565_),
    .ZN(_10566_)
  );
  AND2_X1 _45012_ (
    .A1(_21190_),
    .A2(_22229_),
    .ZN(_10567_)
  );
  INV_X1 _45013_ (
    .A(_10567_),
    .ZN(_10568_)
  );
  AND2_X1 _45014_ (
    .A1(reg_op1[22]),
    .A2(_29151_[22]),
    .ZN(_10569_)
  );
  INV_X1 _45015_ (
    .A(_10569_),
    .ZN(_10570_)
  );
  AND2_X1 _45016_ (
    .A1(_21189_),
    .A2(_22242_),
    .ZN(_10571_)
  );
  INV_X1 _45017_ (
    .A(_10571_),
    .ZN(_10572_)
  );
  AND2_X1 _45018_ (
    .A1(_10570_),
    .A2(_10572_),
    .ZN(_10573_)
  );
  INV_X1 _45019_ (
    .A(_10573_),
    .ZN(_10574_)
  );
  AND2_X1 _45020_ (
    .A1(reg_op1[21]),
    .A2(_29151_[21]),
    .ZN(_10575_)
  );
  INV_X1 _45021_ (
    .A(_10575_),
    .ZN(_10576_)
  );
  AND2_X1 _45022_ (
    .A1(_21188_),
    .A2(_22247_),
    .ZN(_10577_)
  );
  INV_X1 _45023_ (
    .A(_10577_),
    .ZN(_10578_)
  );
  AND2_X1 _45024_ (
    .A1(reg_op1[20]),
    .A2(_29151_[20]),
    .ZN(_10579_)
  );
  INV_X1 _45025_ (
    .A(_10579_),
    .ZN(_10580_)
  );
  AND2_X1 _45026_ (
    .A1(_21187_),
    .A2(_22228_),
    .ZN(_10581_)
  );
  INV_X1 _45027_ (
    .A(_10581_),
    .ZN(_10582_)
  );
  AND2_X1 _45028_ (
    .A1(_10580_),
    .A2(_10582_),
    .ZN(_10583_)
  );
  INV_X1 _45029_ (
    .A(_10583_),
    .ZN(_10584_)
  );
  AND2_X1 _45030_ (
    .A1(reg_op1[19]),
    .A2(_29151_[19]),
    .ZN(_10585_)
  );
  INV_X1 _45031_ (
    .A(_10585_),
    .ZN(_10586_)
  );
  AND2_X1 _45032_ (
    .A1(_21186_),
    .A2(_22227_),
    .ZN(_10587_)
  );
  INV_X1 _45033_ (
    .A(_10587_),
    .ZN(_10588_)
  );
  AND2_X1 _45034_ (
    .A1(reg_op1[18]),
    .A2(_29151_[18]),
    .ZN(_10589_)
  );
  INV_X1 _45035_ (
    .A(_10589_),
    .ZN(_10590_)
  );
  AND2_X1 _45036_ (
    .A1(_21185_),
    .A2(_22226_),
    .ZN(_10591_)
  );
  INV_X1 _45037_ (
    .A(_10591_),
    .ZN(_10592_)
  );
  AND2_X1 _45038_ (
    .A1(_10590_),
    .A2(_10592_),
    .ZN(_10593_)
  );
  INV_X1 _45039_ (
    .A(_10593_),
    .ZN(_10594_)
  );
  AND2_X1 _45040_ (
    .A1(reg_op1[17]),
    .A2(_29151_[17]),
    .ZN(_10595_)
  );
  INV_X1 _45041_ (
    .A(_10595_),
    .ZN(_10596_)
  );
  AND2_X1 _45042_ (
    .A1(_21184_),
    .A2(_22239_),
    .ZN(_10597_)
  );
  INV_X1 _45043_ (
    .A(_10597_),
    .ZN(_10598_)
  );
  AND2_X1 _45044_ (
    .A1(reg_op1[16]),
    .A2(_29151_[16]),
    .ZN(_10599_)
  );
  INV_X1 _45045_ (
    .A(_10599_),
    .ZN(_10600_)
  );
  AND2_X1 _45046_ (
    .A1(_21183_),
    .A2(_22225_),
    .ZN(_10601_)
  );
  INV_X1 _45047_ (
    .A(_10601_),
    .ZN(_10602_)
  );
  AND2_X1 _45048_ (
    .A1(_10600_),
    .A2(_10602_),
    .ZN(_10603_)
  );
  INV_X1 _45049_ (
    .A(_10603_),
    .ZN(_10604_)
  );
  AND2_X1 _45050_ (
    .A1(reg_op1[15]),
    .A2(_29151_[15]),
    .ZN(_10605_)
  );
  INV_X1 _45051_ (
    .A(_10605_),
    .ZN(_10606_)
  );
  AND2_X1 _45052_ (
    .A1(_21182_),
    .A2(_22224_),
    .ZN(_10607_)
  );
  INV_X1 _45053_ (
    .A(_10607_),
    .ZN(_10608_)
  );
  AND2_X1 _45054_ (
    .A1(reg_op1[14]),
    .A2(_29151_[14]),
    .ZN(_10609_)
  );
  INV_X1 _45055_ (
    .A(_10609_),
    .ZN(_10610_)
  );
  AND2_X1 _45056_ (
    .A1(_21181_),
    .A2(_22223_),
    .ZN(_10611_)
  );
  INV_X1 _45057_ (
    .A(_10611_),
    .ZN(_10612_)
  );
  AND2_X1 _45058_ (
    .A1(_10610_),
    .A2(_10612_),
    .ZN(_10613_)
  );
  INV_X1 _45059_ (
    .A(_10613_),
    .ZN(_10614_)
  );
  AND2_X1 _45060_ (
    .A1(reg_op1[13]),
    .A2(_29151_[13]),
    .ZN(_10615_)
  );
  INV_X1 _45061_ (
    .A(_10615_),
    .ZN(_10616_)
  );
  AND2_X1 _45062_ (
    .A1(_21180_),
    .A2(_22246_),
    .ZN(_10617_)
  );
  INV_X1 _45063_ (
    .A(_10617_),
    .ZN(_10618_)
  );
  AND2_X1 _45064_ (
    .A1(reg_op1[12]),
    .A2(_29151_[12]),
    .ZN(_10619_)
  );
  INV_X1 _45065_ (
    .A(_10619_),
    .ZN(_10620_)
  );
  AND2_X1 _45066_ (
    .A1(_21179_),
    .A2(_22245_),
    .ZN(_10621_)
  );
  INV_X1 _45067_ (
    .A(_10621_),
    .ZN(_10622_)
  );
  AND2_X1 _45068_ (
    .A1(_10620_),
    .A2(_10622_),
    .ZN(_10623_)
  );
  INV_X1 _45069_ (
    .A(_10623_),
    .ZN(_10624_)
  );
  AND2_X1 _45070_ (
    .A1(reg_op1[11]),
    .A2(_29151_[11]),
    .ZN(_10625_)
  );
  INV_X1 _45071_ (
    .A(_10625_),
    .ZN(_10626_)
  );
  AND2_X1 _45072_ (
    .A1(_21178_),
    .A2(_22222_),
    .ZN(_10627_)
  );
  INV_X1 _45073_ (
    .A(_10627_),
    .ZN(_10628_)
  );
  AND2_X1 _45074_ (
    .A1(reg_op1[10]),
    .A2(_29151_[10]),
    .ZN(_10629_)
  );
  INV_X1 _45075_ (
    .A(_10629_),
    .ZN(_10630_)
  );
  AND2_X1 _45076_ (
    .A1(_21177_),
    .A2(_22221_),
    .ZN(_10631_)
  );
  INV_X1 _45077_ (
    .A(_10631_),
    .ZN(_10632_)
  );
  AND2_X1 _45078_ (
    .A1(_10630_),
    .A2(_10632_),
    .ZN(_10633_)
  );
  INV_X1 _45079_ (
    .A(_10633_),
    .ZN(_10634_)
  );
  AND2_X1 _45080_ (
    .A1(reg_op1[9]),
    .A2(_29151_[9]),
    .ZN(_10635_)
  );
  INV_X1 _45081_ (
    .A(_10635_),
    .ZN(_10636_)
  );
  AND2_X1 _45082_ (
    .A1(_21176_),
    .A2(_22220_),
    .ZN(_10637_)
  );
  INV_X1 _45083_ (
    .A(_10637_),
    .ZN(_10638_)
  );
  AND2_X1 _45084_ (
    .A1(reg_op1[8]),
    .A2(_29151_[8]),
    .ZN(_10639_)
  );
  INV_X1 _45085_ (
    .A(_10639_),
    .ZN(_10640_)
  );
  AND2_X1 _45086_ (
    .A1(_21175_),
    .A2(_22244_),
    .ZN(_10641_)
  );
  INV_X1 _45087_ (
    .A(_10641_),
    .ZN(_10642_)
  );
  AND2_X1 _45088_ (
    .A1(_10640_),
    .A2(_10642_),
    .ZN(_10643_)
  );
  INV_X1 _45089_ (
    .A(_10643_),
    .ZN(_10644_)
  );
  AND2_X1 _45090_ (
    .A1(reg_op1[7]),
    .A2(_29151_[7]),
    .ZN(_10645_)
  );
  INV_X1 _45091_ (
    .A(_10645_),
    .ZN(_10646_)
  );
  AND2_X1 _45092_ (
    .A1(_21174_),
    .A2(_22243_),
    .ZN(_10647_)
  );
  INV_X1 _45093_ (
    .A(_10647_),
    .ZN(_10648_)
  );
  AND2_X1 _45094_ (
    .A1(reg_op1[6]),
    .A2(_29151_[6]),
    .ZN(_10649_)
  );
  INV_X1 _45095_ (
    .A(_10649_),
    .ZN(_10650_)
  );
  AND2_X1 _45096_ (
    .A1(_21173_),
    .A2(_22238_),
    .ZN(_10651_)
  );
  INV_X1 _45097_ (
    .A(_10651_),
    .ZN(_10652_)
  );
  AND2_X1 _45098_ (
    .A1(_10650_),
    .A2(_10652_),
    .ZN(_10653_)
  );
  INV_X1 _45099_ (
    .A(_10653_),
    .ZN(_10654_)
  );
  AND2_X1 _45100_ (
    .A1(reg_op1[5]),
    .A2(_29151_[5]),
    .ZN(_10655_)
  );
  INV_X1 _45101_ (
    .A(_10655_),
    .ZN(_10656_)
  );
  AND2_X1 _45102_ (
    .A1(_21172_),
    .A2(_22237_),
    .ZN(_10657_)
  );
  INV_X1 _45103_ (
    .A(_10657_),
    .ZN(_10658_)
  );
  AND2_X1 _45104_ (
    .A1(reg_op1[4]),
    .A2(_29151_[4]),
    .ZN(_10659_)
  );
  INV_X1 _45105_ (
    .A(_10659_),
    .ZN(_10660_)
  );
  AND2_X1 _45106_ (
    .A1(_21171_),
    .A2(_22236_),
    .ZN(_10661_)
  );
  INV_X1 _45107_ (
    .A(_10661_),
    .ZN(_10662_)
  );
  AND2_X1 _45108_ (
    .A1(_10660_),
    .A2(_10662_),
    .ZN(_10663_)
  );
  INV_X1 _45109_ (
    .A(_10663_),
    .ZN(_10664_)
  );
  AND2_X1 _45110_ (
    .A1(reg_op1[3]),
    .A2(_29151_[3]),
    .ZN(_10665_)
  );
  INV_X1 _45111_ (
    .A(_10665_),
    .ZN(_10666_)
  );
  AND2_X1 _45112_ (
    .A1(_21170_),
    .A2(_22235_),
    .ZN(_10667_)
  );
  INV_X1 _45113_ (
    .A(_10667_),
    .ZN(_10668_)
  );
  AND2_X1 _45114_ (
    .A1(reg_op1[2]),
    .A2(_29151_[2]),
    .ZN(_10669_)
  );
  INV_X1 _45115_ (
    .A(_10669_),
    .ZN(_10670_)
  );
  AND2_X1 _45116_ (
    .A1(reg_op1[1]),
    .A2(_29151_[1]),
    .ZN(_10671_)
  );
  INV_X1 _45117_ (
    .A(_10671_),
    .ZN(_10672_)
  );
  AND2_X1 _45118_ (
    .A1(_21168_),
    .A2(_22232_),
    .ZN(_10673_)
  );
  INV_X1 _45119_ (
    .A(_10673_),
    .ZN(_10674_)
  );
  AND2_X1 _45120_ (
    .A1(_22024_),
    .A2(_22233_),
    .ZN(_10675_)
  );
  INV_X1 _45121_ (
    .A(_10675_),
    .ZN(_10676_)
  );
  AND2_X1 _45122_ (
    .A1(_10672_),
    .A2(_10676_),
    .ZN(_10677_)
  );
  INV_X1 _45123_ (
    .A(_10677_),
    .ZN(_10678_)
  );
  AND2_X1 _45124_ (
    .A1(_10674_),
    .A2(_10677_),
    .ZN(_10679_)
  );
  INV_X1 _45125_ (
    .A(_10679_),
    .ZN(_10680_)
  );
  AND2_X1 _45126_ (
    .A1(_10672_),
    .A2(_10680_),
    .ZN(_10681_)
  );
  INV_X1 _45127_ (
    .A(_10681_),
    .ZN(_10682_)
  );
  AND2_X1 _45128_ (
    .A1(_21169_),
    .A2(_22234_),
    .ZN(_10683_)
  );
  INV_X1 _45129_ (
    .A(_10683_),
    .ZN(_10684_)
  );
  AND2_X1 _45130_ (
    .A1(_10670_),
    .A2(_10684_),
    .ZN(_10685_)
  );
  INV_X1 _45131_ (
    .A(_10685_),
    .ZN(_10686_)
  );
  AND2_X1 _45132_ (
    .A1(_10682_),
    .A2(_10685_),
    .ZN(_10687_)
  );
  INV_X1 _45133_ (
    .A(_10687_),
    .ZN(_10688_)
  );
  AND2_X1 _45134_ (
    .A1(_10670_),
    .A2(_10688_),
    .ZN(_10689_)
  );
  INV_X1 _45135_ (
    .A(_10689_),
    .ZN(_10690_)
  );
  AND2_X1 _45136_ (
    .A1(_10668_),
    .A2(_10690_),
    .ZN(_10691_)
  );
  INV_X1 _45137_ (
    .A(_10691_),
    .ZN(_10692_)
  );
  AND2_X1 _45138_ (
    .A1(_10666_),
    .A2(_10689_),
    .ZN(_10693_)
  );
  INV_X1 _45139_ (
    .A(_10693_),
    .ZN(_10694_)
  );
  AND2_X1 _45140_ (
    .A1(_10666_),
    .A2(_10692_),
    .ZN(_10695_)
  );
  AND2_X1 _45141_ (
    .A1(_10668_),
    .A2(_10694_),
    .ZN(_10696_)
  );
  AND2_X1 _45142_ (
    .A1(_10663_),
    .A2(_10696_),
    .ZN(_10697_)
  );
  INV_X1 _45143_ (
    .A(_10697_),
    .ZN(_10698_)
  );
  AND2_X1 _45144_ (
    .A1(_10660_),
    .A2(_10698_),
    .ZN(_10699_)
  );
  INV_X1 _45145_ (
    .A(_10699_),
    .ZN(_10700_)
  );
  AND2_X1 _45146_ (
    .A1(_10658_),
    .A2(_10700_),
    .ZN(_10701_)
  );
  INV_X1 _45147_ (
    .A(_10701_),
    .ZN(_10702_)
  );
  AND2_X1 _45148_ (
    .A1(_10656_),
    .A2(_10699_),
    .ZN(_10703_)
  );
  INV_X1 _45149_ (
    .A(_10703_),
    .ZN(_10704_)
  );
  AND2_X1 _45150_ (
    .A1(_10656_),
    .A2(_10702_),
    .ZN(_10705_)
  );
  AND2_X1 _45151_ (
    .A1(_10658_),
    .A2(_10704_),
    .ZN(_10706_)
  );
  AND2_X1 _45152_ (
    .A1(_10653_),
    .A2(_10706_),
    .ZN(_10707_)
  );
  INV_X1 _45153_ (
    .A(_10707_),
    .ZN(_10708_)
  );
  AND2_X1 _45154_ (
    .A1(_10650_),
    .A2(_10708_),
    .ZN(_10709_)
  );
  INV_X1 _45155_ (
    .A(_10709_),
    .ZN(_10710_)
  );
  AND2_X1 _45156_ (
    .A1(_10648_),
    .A2(_10710_),
    .ZN(_10711_)
  );
  INV_X1 _45157_ (
    .A(_10711_),
    .ZN(_10712_)
  );
  AND2_X1 _45158_ (
    .A1(_10646_),
    .A2(_10709_),
    .ZN(_10713_)
  );
  INV_X1 _45159_ (
    .A(_10713_),
    .ZN(_10714_)
  );
  AND2_X1 _45160_ (
    .A1(_10646_),
    .A2(_10712_),
    .ZN(_10715_)
  );
  AND2_X1 _45161_ (
    .A1(_10648_),
    .A2(_10714_),
    .ZN(_10716_)
  );
  AND2_X1 _45162_ (
    .A1(_10643_),
    .A2(_10716_),
    .ZN(_10717_)
  );
  INV_X1 _45163_ (
    .A(_10717_),
    .ZN(_10718_)
  );
  AND2_X1 _45164_ (
    .A1(_10640_),
    .A2(_10718_),
    .ZN(_10719_)
  );
  INV_X1 _45165_ (
    .A(_10719_),
    .ZN(_10720_)
  );
  AND2_X1 _45166_ (
    .A1(_10638_),
    .A2(_10720_),
    .ZN(_10721_)
  );
  INV_X1 _45167_ (
    .A(_10721_),
    .ZN(_10722_)
  );
  AND2_X1 _45168_ (
    .A1(_10636_),
    .A2(_10719_),
    .ZN(_10723_)
  );
  INV_X1 _45169_ (
    .A(_10723_),
    .ZN(_10724_)
  );
  AND2_X1 _45170_ (
    .A1(_10636_),
    .A2(_10722_),
    .ZN(_10725_)
  );
  AND2_X1 _45171_ (
    .A1(_10638_),
    .A2(_10724_),
    .ZN(_10726_)
  );
  AND2_X1 _45172_ (
    .A1(_10633_),
    .A2(_10726_),
    .ZN(_10727_)
  );
  INV_X1 _45173_ (
    .A(_10727_),
    .ZN(_10728_)
  );
  AND2_X1 _45174_ (
    .A1(_10630_),
    .A2(_10728_),
    .ZN(_10729_)
  );
  INV_X1 _45175_ (
    .A(_10729_),
    .ZN(_10730_)
  );
  AND2_X1 _45176_ (
    .A1(_10628_),
    .A2(_10730_),
    .ZN(_10731_)
  );
  INV_X1 _45177_ (
    .A(_10731_),
    .ZN(_10732_)
  );
  AND2_X1 _45178_ (
    .A1(_10626_),
    .A2(_10729_),
    .ZN(_10733_)
  );
  INV_X1 _45179_ (
    .A(_10733_),
    .ZN(_10734_)
  );
  AND2_X1 _45180_ (
    .A1(_10626_),
    .A2(_10732_),
    .ZN(_10735_)
  );
  AND2_X1 _45181_ (
    .A1(_10628_),
    .A2(_10734_),
    .ZN(_10736_)
  );
  AND2_X1 _45182_ (
    .A1(_10623_),
    .A2(_10736_),
    .ZN(_10737_)
  );
  INV_X1 _45183_ (
    .A(_10737_),
    .ZN(_10738_)
  );
  AND2_X1 _45184_ (
    .A1(_10620_),
    .A2(_10738_),
    .ZN(_10739_)
  );
  INV_X1 _45185_ (
    .A(_10739_),
    .ZN(_10740_)
  );
  AND2_X1 _45186_ (
    .A1(_10618_),
    .A2(_10740_),
    .ZN(_10741_)
  );
  INV_X1 _45187_ (
    .A(_10741_),
    .ZN(_10742_)
  );
  AND2_X1 _45188_ (
    .A1(_10616_),
    .A2(_10739_),
    .ZN(_10743_)
  );
  INV_X1 _45189_ (
    .A(_10743_),
    .ZN(_10744_)
  );
  AND2_X1 _45190_ (
    .A1(_10616_),
    .A2(_10742_),
    .ZN(_10745_)
  );
  AND2_X1 _45191_ (
    .A1(_10618_),
    .A2(_10744_),
    .ZN(_10746_)
  );
  AND2_X1 _45192_ (
    .A1(_10613_),
    .A2(_10746_),
    .ZN(_10747_)
  );
  INV_X1 _45193_ (
    .A(_10747_),
    .ZN(_10748_)
  );
  AND2_X1 _45194_ (
    .A1(_10610_),
    .A2(_10748_),
    .ZN(_10749_)
  );
  INV_X1 _45195_ (
    .A(_10749_),
    .ZN(_10750_)
  );
  AND2_X1 _45196_ (
    .A1(_10608_),
    .A2(_10750_),
    .ZN(_10751_)
  );
  INV_X1 _45197_ (
    .A(_10751_),
    .ZN(_10752_)
  );
  AND2_X1 _45198_ (
    .A1(_10606_),
    .A2(_10749_),
    .ZN(_10753_)
  );
  INV_X1 _45199_ (
    .A(_10753_),
    .ZN(_10754_)
  );
  AND2_X1 _45200_ (
    .A1(_10606_),
    .A2(_10752_),
    .ZN(_10755_)
  );
  AND2_X1 _45201_ (
    .A1(_10608_),
    .A2(_10754_),
    .ZN(_10756_)
  );
  AND2_X1 _45202_ (
    .A1(_10603_),
    .A2(_10756_),
    .ZN(_10757_)
  );
  INV_X1 _45203_ (
    .A(_10757_),
    .ZN(_10758_)
  );
  AND2_X1 _45204_ (
    .A1(_10600_),
    .A2(_10758_),
    .ZN(_10759_)
  );
  INV_X1 _45205_ (
    .A(_10759_),
    .ZN(_10760_)
  );
  AND2_X1 _45206_ (
    .A1(_10598_),
    .A2(_10760_),
    .ZN(_10761_)
  );
  INV_X1 _45207_ (
    .A(_10761_),
    .ZN(_10762_)
  );
  AND2_X1 _45208_ (
    .A1(_10596_),
    .A2(_10759_),
    .ZN(_10763_)
  );
  INV_X1 _45209_ (
    .A(_10763_),
    .ZN(_10764_)
  );
  AND2_X1 _45210_ (
    .A1(_10596_),
    .A2(_10762_),
    .ZN(_10765_)
  );
  AND2_X1 _45211_ (
    .A1(_10598_),
    .A2(_10764_),
    .ZN(_10766_)
  );
  AND2_X1 _45212_ (
    .A1(_10593_),
    .A2(_10766_),
    .ZN(_10767_)
  );
  INV_X1 _45213_ (
    .A(_10767_),
    .ZN(_10768_)
  );
  AND2_X1 _45214_ (
    .A1(_10590_),
    .A2(_10768_),
    .ZN(_10769_)
  );
  INV_X1 _45215_ (
    .A(_10769_),
    .ZN(_10770_)
  );
  AND2_X1 _45216_ (
    .A1(_10588_),
    .A2(_10770_),
    .ZN(_10771_)
  );
  INV_X1 _45217_ (
    .A(_10771_),
    .ZN(_10772_)
  );
  AND2_X1 _45218_ (
    .A1(_10586_),
    .A2(_10769_),
    .ZN(_10773_)
  );
  INV_X1 _45219_ (
    .A(_10773_),
    .ZN(_10774_)
  );
  AND2_X1 _45220_ (
    .A1(_10586_),
    .A2(_10772_),
    .ZN(_10775_)
  );
  AND2_X1 _45221_ (
    .A1(_10588_),
    .A2(_10774_),
    .ZN(_10776_)
  );
  AND2_X1 _45222_ (
    .A1(_10583_),
    .A2(_10776_),
    .ZN(_10777_)
  );
  INV_X1 _45223_ (
    .A(_10777_),
    .ZN(_10778_)
  );
  AND2_X1 _45224_ (
    .A1(_10580_),
    .A2(_10778_),
    .ZN(_10779_)
  );
  INV_X1 _45225_ (
    .A(_10779_),
    .ZN(_10780_)
  );
  AND2_X1 _45226_ (
    .A1(_10578_),
    .A2(_10780_),
    .ZN(_10781_)
  );
  INV_X1 _45227_ (
    .A(_10781_),
    .ZN(_10782_)
  );
  AND2_X1 _45228_ (
    .A1(_10576_),
    .A2(_10779_),
    .ZN(_10783_)
  );
  INV_X1 _45229_ (
    .A(_10783_),
    .ZN(_10784_)
  );
  AND2_X1 _45230_ (
    .A1(_10576_),
    .A2(_10782_),
    .ZN(_10785_)
  );
  AND2_X1 _45231_ (
    .A1(_10578_),
    .A2(_10784_),
    .ZN(_10786_)
  );
  AND2_X1 _45232_ (
    .A1(_10573_),
    .A2(_10786_),
    .ZN(_10787_)
  );
  INV_X1 _45233_ (
    .A(_10787_),
    .ZN(_10788_)
  );
  AND2_X1 _45234_ (
    .A1(_10570_),
    .A2(_10788_),
    .ZN(_10789_)
  );
  INV_X1 _45235_ (
    .A(_10789_),
    .ZN(_10790_)
  );
  AND2_X1 _45236_ (
    .A1(_10568_),
    .A2(_10790_),
    .ZN(_10791_)
  );
  INV_X1 _45237_ (
    .A(_10791_),
    .ZN(_10792_)
  );
  AND2_X1 _45238_ (
    .A1(_10566_),
    .A2(_10789_),
    .ZN(_10793_)
  );
  INV_X1 _45239_ (
    .A(_10793_),
    .ZN(_10794_)
  );
  AND2_X1 _45240_ (
    .A1(_10566_),
    .A2(_10792_),
    .ZN(_10795_)
  );
  AND2_X1 _45241_ (
    .A1(_10568_),
    .A2(_10794_),
    .ZN(_10796_)
  );
  AND2_X1 _45242_ (
    .A1(_10563_),
    .A2(_10796_),
    .ZN(_10797_)
  );
  INV_X1 _45243_ (
    .A(_10797_),
    .ZN(_10798_)
  );
  AND2_X1 _45244_ (
    .A1(_10560_),
    .A2(_10798_),
    .ZN(_10799_)
  );
  INV_X1 _45245_ (
    .A(_10799_),
    .ZN(_10800_)
  );
  AND2_X1 _45246_ (
    .A1(_10558_),
    .A2(_10800_),
    .ZN(_10801_)
  );
  INV_X1 _45247_ (
    .A(_10801_),
    .ZN(_10802_)
  );
  AND2_X1 _45248_ (
    .A1(_10556_),
    .A2(_10799_),
    .ZN(_10803_)
  );
  INV_X1 _45249_ (
    .A(_10803_),
    .ZN(_10804_)
  );
  AND2_X1 _45250_ (
    .A1(_10556_),
    .A2(_10802_),
    .ZN(_10805_)
  );
  AND2_X1 _45251_ (
    .A1(_10558_),
    .A2(_10804_),
    .ZN(_10806_)
  );
  AND2_X1 _45252_ (
    .A1(_10553_),
    .A2(_10806_),
    .ZN(_10807_)
  );
  INV_X1 _45253_ (
    .A(_10807_),
    .ZN(_10808_)
  );
  AND2_X1 _45254_ (
    .A1(_10550_),
    .A2(_10808_),
    .ZN(_10809_)
  );
  INV_X1 _45255_ (
    .A(_10809_),
    .ZN(_10810_)
  );
  AND2_X1 _45256_ (
    .A1(_10548_),
    .A2(_10810_),
    .ZN(_10811_)
  );
  INV_X1 _45257_ (
    .A(_10811_),
    .ZN(_10812_)
  );
  AND2_X1 _45258_ (
    .A1(_10546_),
    .A2(_10809_),
    .ZN(_10813_)
  );
  INV_X1 _45259_ (
    .A(_10813_),
    .ZN(_10814_)
  );
  AND2_X1 _45260_ (
    .A1(_10546_),
    .A2(_10812_),
    .ZN(_10815_)
  );
  AND2_X1 _45261_ (
    .A1(_10548_),
    .A2(_10814_),
    .ZN(_10816_)
  );
  AND2_X1 _45262_ (
    .A1(_10543_),
    .A2(_10816_),
    .ZN(_10817_)
  );
  INV_X1 _45263_ (
    .A(_10817_),
    .ZN(_10818_)
  );
  AND2_X1 _45264_ (
    .A1(reg_op1[29]),
    .A2(_29151_[29]),
    .ZN(_10819_)
  );
  INV_X1 _45265_ (
    .A(_10819_),
    .ZN(_10820_)
  );
  AND2_X1 _45266_ (
    .A1(_10540_),
    .A2(_10820_),
    .ZN(_10821_)
  );
  AND2_X1 _45267_ (
    .A1(_10818_),
    .A2(_10821_),
    .ZN(_10822_)
  );
  INV_X1 _45268_ (
    .A(_10822_),
    .ZN(_10823_)
  );
  AND2_X1 _45269_ (
    .A1(_10538_),
    .A2(_10820_),
    .ZN(_10824_)
  );
  INV_X1 _45270_ (
    .A(_10824_),
    .ZN(_10825_)
  );
  AND2_X1 _45271_ (
    .A1(_10538_),
    .A2(_10823_),
    .ZN(_10826_)
  );
  INV_X1 _45272_ (
    .A(_10826_),
    .ZN(_10827_)
  );
  AND2_X1 _45273_ (
    .A1(_10535_),
    .A2(_10826_),
    .ZN(_10828_)
  );
  INV_X1 _45274_ (
    .A(_10828_),
    .ZN(_10829_)
  );
  AND2_X1 _45275_ (
    .A1(_10532_),
    .A2(_10829_),
    .ZN(_10830_)
  );
  INV_X1 _45276_ (
    .A(_10830_),
    .ZN(_10831_)
  );
  AND2_X1 _45277_ (
    .A1(_10529_),
    .A2(_10830_),
    .ZN(_10832_)
  );
  INV_X1 _45278_ (
    .A(_10832_),
    .ZN(_10833_)
  );
  AND2_X1 _45279_ (
    .A1(_10526_),
    .A2(_10833_),
    .ZN(_10834_)
  );
  INV_X1 _45280_ (
    .A(_10834_),
    .ZN(_10835_)
  );
  AND2_X1 _45281_ (
    .A1(is_slti_blt_slt),
    .A2(_10835_),
    .ZN(_10836_)
  );
  INV_X1 _45282_ (
    .A(_10836_),
    .ZN(_10837_)
  );
  AND2_X1 _45283_ (
    .A1(instr_bge),
    .A2(_10834_),
    .ZN(_10838_)
  );
  INV_X1 _45284_ (
    .A(_10838_),
    .ZN(_10839_)
  );
  AND2_X1 _45285_ (
    .A1(_10526_),
    .A2(_10532_),
    .ZN(_10840_)
  );
  INV_X1 _45286_ (
    .A(_10840_),
    .ZN(_10841_)
  );
  AND2_X1 _45287_ (
    .A1(_10528_),
    .A2(_10841_),
    .ZN(_10842_)
  );
  INV_X1 _45288_ (
    .A(_10842_),
    .ZN(_10843_)
  );
  AND2_X1 _45289_ (
    .A1(_10529_),
    .A2(_10535_),
    .ZN(_10844_)
  );
  AND2_X1 _45290_ (
    .A1(_10826_),
    .A2(_10844_),
    .ZN(_10845_)
  );
  INV_X1 _45291_ (
    .A(_10845_),
    .ZN(_10846_)
  );
  AND2_X1 _45292_ (
    .A1(_10843_),
    .A2(_10846_),
    .ZN(_10847_)
  );
  INV_X1 _45293_ (
    .A(_10847_),
    .ZN(_10848_)
  );
  AND2_X1 _45294_ (
    .A1(instr_bgeu),
    .A2(_10848_),
    .ZN(_10849_)
  );
  INV_X1 _45295_ (
    .A(_10849_),
    .ZN(_10850_)
  );
  AND2_X1 _45296_ (
    .A1(reg_op2[1]),
    .A2(reg_op1[1]),
    .ZN(_10851_)
  );
  INV_X1 _45297_ (
    .A(_10851_),
    .ZN(_10852_)
  );
  AND2_X1 _45298_ (
    .A1(_21201_),
    .A2(_22024_),
    .ZN(_10853_)
  );
  INV_X1 _45299_ (
    .A(_10853_),
    .ZN(_10854_)
  );
  AND2_X1 _45300_ (
    .A1(_10852_),
    .A2(_10854_),
    .ZN(_10855_)
  );
  INV_X1 _45301_ (
    .A(_10855_),
    .ZN(_10856_)
  );
  AND2_X1 _45302_ (
    .A1(reg_op1[9]),
    .A2(reg_op2[9]),
    .ZN(_10857_)
  );
  INV_X1 _45303_ (
    .A(_10857_),
    .ZN(_10858_)
  );
  AND2_X1 _45304_ (
    .A1(_21176_),
    .A2(_21209_),
    .ZN(_10859_)
  );
  INV_X1 _45305_ (
    .A(_10859_),
    .ZN(_10860_)
  );
  AND2_X1 _45306_ (
    .A1(_10858_),
    .A2(_10860_),
    .ZN(_10861_)
  );
  INV_X1 _45307_ (
    .A(_10861_),
    .ZN(_10862_)
  );
  AND2_X1 _45308_ (
    .A1(reg_op1[15]),
    .A2(reg_op2[15]),
    .ZN(_10863_)
  );
  INV_X1 _45309_ (
    .A(_10863_),
    .ZN(_10864_)
  );
  AND2_X1 _45310_ (
    .A1(_21182_),
    .A2(_21215_),
    .ZN(_10865_)
  );
  INV_X1 _45311_ (
    .A(_10865_),
    .ZN(_10866_)
  );
  AND2_X1 _45312_ (
    .A1(_10864_),
    .A2(_10866_),
    .ZN(_10867_)
  );
  INV_X1 _45313_ (
    .A(_10867_),
    .ZN(_10868_)
  );
  AND2_X1 _45314_ (
    .A1(reg_op1[8]),
    .A2(reg_op2[8]),
    .ZN(_10869_)
  );
  INV_X1 _45315_ (
    .A(_10869_),
    .ZN(_10870_)
  );
  AND2_X1 _45316_ (
    .A1(_21175_),
    .A2(_21208_),
    .ZN(_10871_)
  );
  INV_X1 _45317_ (
    .A(_10871_),
    .ZN(_10872_)
  );
  AND2_X1 _45318_ (
    .A1(_10870_),
    .A2(_10872_),
    .ZN(_10873_)
  );
  INV_X1 _45319_ (
    .A(_10873_),
    .ZN(_10874_)
  );
  AND2_X1 _45320_ (
    .A1(reg_op1[30]),
    .A2(reg_op2[30]),
    .ZN(_10875_)
  );
  INV_X1 _45321_ (
    .A(_10875_),
    .ZN(_10876_)
  );
  AND2_X1 _45322_ (
    .A1(_21197_),
    .A2(_21230_),
    .ZN(_10877_)
  );
  INV_X1 _45323_ (
    .A(_10877_),
    .ZN(_10878_)
  );
  AND2_X1 _45324_ (
    .A1(_10876_),
    .A2(_10878_),
    .ZN(_10879_)
  );
  INV_X1 _45325_ (
    .A(_10879_),
    .ZN(_10880_)
  );
  AND2_X1 _45326_ (
    .A1(reg_op1[19]),
    .A2(reg_op2[19]),
    .ZN(_10881_)
  );
  INV_X1 _45327_ (
    .A(_10881_),
    .ZN(_10882_)
  );
  AND2_X1 _45328_ (
    .A1(_21186_),
    .A2(_21219_),
    .ZN(_10883_)
  );
  INV_X1 _45329_ (
    .A(_10883_),
    .ZN(_10884_)
  );
  AND2_X1 _45330_ (
    .A1(_10882_),
    .A2(_10884_),
    .ZN(_10885_)
  );
  INV_X1 _45331_ (
    .A(_10885_),
    .ZN(_10886_)
  );
  AND2_X1 _45332_ (
    .A1(reg_op1[14]),
    .A2(reg_op2[14]),
    .ZN(_10887_)
  );
  INV_X1 _45333_ (
    .A(_10887_),
    .ZN(_10888_)
  );
  AND2_X1 _45334_ (
    .A1(_21181_),
    .A2(_21214_),
    .ZN(_10889_)
  );
  INV_X1 _45335_ (
    .A(_10889_),
    .ZN(_10890_)
  );
  AND2_X1 _45336_ (
    .A1(_10888_),
    .A2(_10890_),
    .ZN(_10891_)
  );
  INV_X1 _45337_ (
    .A(_10891_),
    .ZN(_10892_)
  );
  AND2_X1 _45338_ (
    .A1(reg_op1[10]),
    .A2(reg_op2[10]),
    .ZN(_10893_)
  );
  INV_X1 _45339_ (
    .A(_10893_),
    .ZN(_10894_)
  );
  AND2_X1 _45340_ (
    .A1(_21177_),
    .A2(_21210_),
    .ZN(_10895_)
  );
  INV_X1 _45341_ (
    .A(_10895_),
    .ZN(_10896_)
  );
  AND2_X1 _45342_ (
    .A1(_10894_),
    .A2(_10896_),
    .ZN(_10897_)
  );
  INV_X1 _45343_ (
    .A(_10897_),
    .ZN(_10898_)
  );
  AND2_X1 _45344_ (
    .A1(reg_op1[23]),
    .A2(reg_op2[23]),
    .ZN(_10899_)
  );
  INV_X1 _45345_ (
    .A(_10899_),
    .ZN(_10900_)
  );
  AND2_X1 _45346_ (
    .A1(_21190_),
    .A2(_21223_),
    .ZN(_10901_)
  );
  INV_X1 _45347_ (
    .A(_10901_),
    .ZN(_10902_)
  );
  AND2_X1 _45348_ (
    .A1(_10900_),
    .A2(_10902_),
    .ZN(_10903_)
  );
  INV_X1 _45349_ (
    .A(_10903_),
    .ZN(_10904_)
  );
  AND2_X1 _45350_ (
    .A1(reg_op1[11]),
    .A2(reg_op2[11]),
    .ZN(_10905_)
  );
  INV_X1 _45351_ (
    .A(_10905_),
    .ZN(_10906_)
  );
  AND2_X1 _45352_ (
    .A1(_21178_),
    .A2(_21211_),
    .ZN(_10907_)
  );
  INV_X1 _45353_ (
    .A(_10907_),
    .ZN(_10908_)
  );
  AND2_X1 _45354_ (
    .A1(_10906_),
    .A2(_10908_),
    .ZN(_10909_)
  );
  INV_X1 _45355_ (
    .A(_10909_),
    .ZN(_10910_)
  );
  AND2_X1 _45356_ (
    .A1(reg_op1[18]),
    .A2(reg_op2[18]),
    .ZN(_10911_)
  );
  INV_X1 _45357_ (
    .A(_10911_),
    .ZN(_10912_)
  );
  AND2_X1 _45358_ (
    .A1(_21185_),
    .A2(_21218_),
    .ZN(_10913_)
  );
  INV_X1 _45359_ (
    .A(_10913_),
    .ZN(_10914_)
  );
  AND2_X1 _45360_ (
    .A1(_10912_),
    .A2(_10914_),
    .ZN(_10915_)
  );
  INV_X1 _45361_ (
    .A(_10915_),
    .ZN(_10916_)
  );
  AND2_X1 _45362_ (
    .A1(reg_op1[29]),
    .A2(reg_op2[29]),
    .ZN(_10917_)
  );
  INV_X1 _45363_ (
    .A(_10917_),
    .ZN(_10918_)
  );
  AND2_X1 _45364_ (
    .A1(_21196_),
    .A2(_21229_),
    .ZN(_10919_)
  );
  INV_X1 _45365_ (
    .A(_10919_),
    .ZN(_10920_)
  );
  AND2_X1 _45366_ (
    .A1(_10918_),
    .A2(_10920_),
    .ZN(_10921_)
  );
  INV_X1 _45367_ (
    .A(_10921_),
    .ZN(_10922_)
  );
  AND2_X1 _45368_ (
    .A1(reg_op1[3]),
    .A2(reg_op2[3]),
    .ZN(_10923_)
  );
  INV_X1 _45369_ (
    .A(_10923_),
    .ZN(_10924_)
  );
  AND2_X1 _45370_ (
    .A1(_21170_),
    .A2(_21203_),
    .ZN(_10925_)
  );
  INV_X1 _45371_ (
    .A(_10925_),
    .ZN(_10926_)
  );
  AND2_X1 _45372_ (
    .A1(_10924_),
    .A2(_10926_),
    .ZN(_10927_)
  );
  INV_X1 _45373_ (
    .A(_10927_),
    .ZN(_10928_)
  );
  AND2_X1 _45374_ (
    .A1(reg_op1[6]),
    .A2(reg_op2[6]),
    .ZN(_10929_)
  );
  INV_X1 _45375_ (
    .A(_10929_),
    .ZN(_10930_)
  );
  AND2_X1 _45376_ (
    .A1(_21173_),
    .A2(_21206_),
    .ZN(_10931_)
  );
  INV_X1 _45377_ (
    .A(_10931_),
    .ZN(_10932_)
  );
  AND2_X1 _45378_ (
    .A1(_10930_),
    .A2(_10932_),
    .ZN(_10933_)
  );
  INV_X1 _45379_ (
    .A(_10933_),
    .ZN(_10934_)
  );
  AND2_X1 _45380_ (
    .A1(reg_op1[27]),
    .A2(reg_op2[27]),
    .ZN(_10935_)
  );
  INV_X1 _45381_ (
    .A(_10935_),
    .ZN(_10936_)
  );
  AND2_X1 _45382_ (
    .A1(_21194_),
    .A2(_21227_),
    .ZN(_10937_)
  );
  INV_X1 _45383_ (
    .A(_10937_),
    .ZN(_10938_)
  );
  AND2_X1 _45384_ (
    .A1(_10936_),
    .A2(_10938_),
    .ZN(_10939_)
  );
  INV_X1 _45385_ (
    .A(_10939_),
    .ZN(_10940_)
  );
  AND2_X1 _45386_ (
    .A1(reg_op1[16]),
    .A2(reg_op2[16]),
    .ZN(_10941_)
  );
  INV_X1 _45387_ (
    .A(_10941_),
    .ZN(_10942_)
  );
  AND2_X1 _45388_ (
    .A1(_21183_),
    .A2(_21216_),
    .ZN(_10943_)
  );
  INV_X1 _45389_ (
    .A(_10943_),
    .ZN(_10944_)
  );
  AND2_X1 _45390_ (
    .A1(_10942_),
    .A2(_10944_),
    .ZN(_10945_)
  );
  INV_X1 _45391_ (
    .A(_10945_),
    .ZN(_10946_)
  );
  AND2_X1 _45392_ (
    .A1(reg_op1[24]),
    .A2(reg_op2[24]),
    .ZN(_10947_)
  );
  INV_X1 _45393_ (
    .A(_10947_),
    .ZN(_10948_)
  );
  AND2_X1 _45394_ (
    .A1(_21191_),
    .A2(_21224_),
    .ZN(_10949_)
  );
  INV_X1 _45395_ (
    .A(_10949_),
    .ZN(_10950_)
  );
  AND2_X1 _45396_ (
    .A1(_10948_),
    .A2(_10950_),
    .ZN(_10951_)
  );
  INV_X1 _45397_ (
    .A(_10951_),
    .ZN(_10952_)
  );
  AND2_X1 _45398_ (
    .A1(reg_op1[17]),
    .A2(reg_op2[17]),
    .ZN(_10953_)
  );
  INV_X1 _45399_ (
    .A(_10953_),
    .ZN(_10954_)
  );
  AND2_X1 _45400_ (
    .A1(_21184_),
    .A2(_21217_),
    .ZN(_10955_)
  );
  INV_X1 _45401_ (
    .A(_10955_),
    .ZN(_10956_)
  );
  AND2_X1 _45402_ (
    .A1(_10954_),
    .A2(_10956_),
    .ZN(_10957_)
  );
  INV_X1 _45403_ (
    .A(_10957_),
    .ZN(_10958_)
  );
  AND2_X1 _45404_ (
    .A1(reg_op1[7]),
    .A2(reg_op2[7]),
    .ZN(_10959_)
  );
  INV_X1 _45405_ (
    .A(_10959_),
    .ZN(_10960_)
  );
  AND2_X1 _45406_ (
    .A1(_21174_),
    .A2(_21207_),
    .ZN(_10961_)
  );
  INV_X1 _45407_ (
    .A(_10961_),
    .ZN(_10962_)
  );
  AND2_X1 _45408_ (
    .A1(_10960_),
    .A2(_10962_),
    .ZN(_10963_)
  );
  INV_X1 _45409_ (
    .A(_10963_),
    .ZN(_10964_)
  );
  AND2_X1 _45410_ (
    .A1(reg_op1[13]),
    .A2(reg_op2[13]),
    .ZN(_10965_)
  );
  INV_X1 _45411_ (
    .A(_10965_),
    .ZN(_10966_)
  );
  AND2_X1 _45412_ (
    .A1(_21180_),
    .A2(_21213_),
    .ZN(_10967_)
  );
  INV_X1 _45413_ (
    .A(_10967_),
    .ZN(_10968_)
  );
  AND2_X1 _45414_ (
    .A1(_10966_),
    .A2(_10968_),
    .ZN(_10969_)
  );
  INV_X1 _45415_ (
    .A(_10969_),
    .ZN(_10970_)
  );
  AND2_X1 _45416_ (
    .A1(reg_op1[0]),
    .A2(reg_op2[0]),
    .ZN(_10971_)
  );
  INV_X1 _45417_ (
    .A(_10971_),
    .ZN(_10972_)
  );
  AND2_X1 _45418_ (
    .A1(_21168_),
    .A2(_21200_),
    .ZN(_10973_)
  );
  INV_X1 _45419_ (
    .A(_10973_),
    .ZN(_10974_)
  );
  AND2_X1 _45420_ (
    .A1(_10972_),
    .A2(_10974_),
    .ZN(_10975_)
  );
  INV_X1 _45421_ (
    .A(_10975_),
    .ZN(_10976_)
  );
  AND2_X1 _45422_ (
    .A1(reg_op1[22]),
    .A2(reg_op2[22]),
    .ZN(_10977_)
  );
  INV_X1 _45423_ (
    .A(_10977_),
    .ZN(_10978_)
  );
  AND2_X1 _45424_ (
    .A1(_21189_),
    .A2(_21222_),
    .ZN(_10979_)
  );
  INV_X1 _45425_ (
    .A(_10979_),
    .ZN(_10980_)
  );
  AND2_X1 _45426_ (
    .A1(_10978_),
    .A2(_10980_),
    .ZN(_10981_)
  );
  INV_X1 _45427_ (
    .A(_10981_),
    .ZN(_10982_)
  );
  AND2_X1 _45428_ (
    .A1(reg_op1[28]),
    .A2(reg_op2[28]),
    .ZN(_10983_)
  );
  INV_X1 _45429_ (
    .A(_10983_),
    .ZN(_10984_)
  );
  AND2_X1 _45430_ (
    .A1(_21195_),
    .A2(_21228_),
    .ZN(_10985_)
  );
  INV_X1 _45431_ (
    .A(_10985_),
    .ZN(_10986_)
  );
  AND2_X1 _45432_ (
    .A1(_10984_),
    .A2(_10986_),
    .ZN(_10987_)
  );
  INV_X1 _45433_ (
    .A(_10987_),
    .ZN(_10988_)
  );
  AND2_X1 _45434_ (
    .A1(reg_op1[5]),
    .A2(reg_op2[5]),
    .ZN(_10989_)
  );
  INV_X1 _45435_ (
    .A(_10989_),
    .ZN(_10990_)
  );
  AND2_X1 _45436_ (
    .A1(_21172_),
    .A2(_21205_),
    .ZN(_10991_)
  );
  INV_X1 _45437_ (
    .A(_10991_),
    .ZN(_10992_)
  );
  AND2_X1 _45438_ (
    .A1(_10990_),
    .A2(_10992_),
    .ZN(_10993_)
  );
  INV_X1 _45439_ (
    .A(_10993_),
    .ZN(_10994_)
  );
  AND2_X1 _45440_ (
    .A1(reg_op1[31]),
    .A2(reg_op2[31]),
    .ZN(_10995_)
  );
  INV_X1 _45441_ (
    .A(_10995_),
    .ZN(_10996_)
  );
  AND2_X1 _45442_ (
    .A1(_21199_),
    .A2(_21231_),
    .ZN(_10997_)
  );
  INV_X1 _45443_ (
    .A(_10997_),
    .ZN(_10998_)
  );
  AND2_X1 _45444_ (
    .A1(_10996_),
    .A2(_10998_),
    .ZN(_10999_)
  );
  INV_X1 _45445_ (
    .A(_10999_),
    .ZN(_11000_)
  );
  AND2_X1 _45446_ (
    .A1(reg_op1[4]),
    .A2(reg_op2[4]),
    .ZN(_11001_)
  );
  INV_X1 _45447_ (
    .A(_11001_),
    .ZN(_11002_)
  );
  AND2_X1 _45448_ (
    .A1(_21171_),
    .A2(_21204_),
    .ZN(_11003_)
  );
  INV_X1 _45449_ (
    .A(_11003_),
    .ZN(_11004_)
  );
  AND2_X1 _45450_ (
    .A1(_11002_),
    .A2(_11004_),
    .ZN(_11005_)
  );
  INV_X1 _45451_ (
    .A(_11005_),
    .ZN(_11006_)
  );
  AND2_X1 _45452_ (
    .A1(reg_op1[12]),
    .A2(reg_op2[12]),
    .ZN(_11007_)
  );
  INV_X1 _45453_ (
    .A(_11007_),
    .ZN(_11008_)
  );
  AND2_X1 _45454_ (
    .A1(_21179_),
    .A2(_21212_),
    .ZN(_11009_)
  );
  INV_X1 _45455_ (
    .A(_11009_),
    .ZN(_11010_)
  );
  AND2_X1 _45456_ (
    .A1(_11008_),
    .A2(_11010_),
    .ZN(_11011_)
  );
  INV_X1 _45457_ (
    .A(_11011_),
    .ZN(_11012_)
  );
  AND2_X1 _45458_ (
    .A1(reg_op1[26]),
    .A2(reg_op2[26]),
    .ZN(_11013_)
  );
  INV_X1 _45459_ (
    .A(_11013_),
    .ZN(_11014_)
  );
  AND2_X1 _45460_ (
    .A1(_21193_),
    .A2(_21226_),
    .ZN(_11015_)
  );
  INV_X1 _45461_ (
    .A(_11015_),
    .ZN(_11016_)
  );
  AND2_X1 _45462_ (
    .A1(_11014_),
    .A2(_11016_),
    .ZN(_11017_)
  );
  INV_X1 _45463_ (
    .A(_11017_),
    .ZN(_11018_)
  );
  AND2_X1 _45464_ (
    .A1(reg_op1[25]),
    .A2(reg_op2[25]),
    .ZN(_11019_)
  );
  INV_X1 _45465_ (
    .A(_11019_),
    .ZN(_11020_)
  );
  AND2_X1 _45466_ (
    .A1(_21192_),
    .A2(_21225_),
    .ZN(_11021_)
  );
  INV_X1 _45467_ (
    .A(_11021_),
    .ZN(_11022_)
  );
  AND2_X1 _45468_ (
    .A1(_11020_),
    .A2(_11022_),
    .ZN(_11023_)
  );
  INV_X1 _45469_ (
    .A(_11023_),
    .ZN(_11024_)
  );
  AND2_X1 _45470_ (
    .A1(reg_op1[21]),
    .A2(reg_op2[21]),
    .ZN(_11025_)
  );
  INV_X1 _45471_ (
    .A(_11025_),
    .ZN(_11026_)
  );
  AND2_X1 _45472_ (
    .A1(_21188_),
    .A2(_21221_),
    .ZN(_11027_)
  );
  INV_X1 _45473_ (
    .A(_11027_),
    .ZN(_11028_)
  );
  AND2_X1 _45474_ (
    .A1(_11026_),
    .A2(_11028_),
    .ZN(_11029_)
  );
  INV_X1 _45475_ (
    .A(_11029_),
    .ZN(_11030_)
  );
  AND2_X1 _45476_ (
    .A1(reg_op1[2]),
    .A2(reg_op2[2]),
    .ZN(_11031_)
  );
  INV_X1 _45477_ (
    .A(_11031_),
    .ZN(_11032_)
  );
  AND2_X1 _45478_ (
    .A1(_21169_),
    .A2(_21202_),
    .ZN(_11033_)
  );
  INV_X1 _45479_ (
    .A(_11033_),
    .ZN(_11034_)
  );
  AND2_X1 _45480_ (
    .A1(_11032_),
    .A2(_11034_),
    .ZN(_11035_)
  );
  INV_X1 _45481_ (
    .A(_11035_),
    .ZN(_11036_)
  );
  AND2_X1 _45482_ (
    .A1(reg_op1[20]),
    .A2(reg_op2[20]),
    .ZN(_11037_)
  );
  INV_X1 _45483_ (
    .A(_11037_),
    .ZN(_11038_)
  );
  AND2_X1 _45484_ (
    .A1(_21187_),
    .A2(_21220_),
    .ZN(_11039_)
  );
  INV_X1 _45485_ (
    .A(_11039_),
    .ZN(_11040_)
  );
  AND2_X1 _45486_ (
    .A1(_11038_),
    .A2(_11040_),
    .ZN(_11041_)
  );
  INV_X1 _45487_ (
    .A(_11041_),
    .ZN(_11042_)
  );
  AND2_X1 _45488_ (
    .A1(_10874_),
    .A2(_11036_),
    .ZN(_11043_)
  );
  AND2_X1 _45489_ (
    .A1(_10868_),
    .A2(_11006_),
    .ZN(_11044_)
  );
  AND2_X1 _45490_ (
    .A1(_11043_),
    .A2(_11044_),
    .ZN(_11045_)
  );
  AND2_X1 _45491_ (
    .A1(_10898_),
    .A2(_11030_),
    .ZN(_11046_)
  );
  AND2_X1 _45492_ (
    .A1(_10892_),
    .A2(_11042_),
    .ZN(_11047_)
  );
  AND2_X1 _45493_ (
    .A1(_11046_),
    .A2(_11047_),
    .ZN(_11048_)
  );
  AND2_X1 _45494_ (
    .A1(_11045_),
    .A2(_11048_),
    .ZN(_11049_)
  );
  AND2_X1 _45495_ (
    .A1(_10922_),
    .A2(_10946_),
    .ZN(_11050_)
  );
  AND2_X1 _45496_ (
    .A1(_10916_),
    .A2(_10940_),
    .ZN(_11051_)
  );
  AND2_X1 _45497_ (
    .A1(_11050_),
    .A2(_11051_),
    .ZN(_11052_)
  );
  AND2_X1 _45498_ (
    .A1(_10928_),
    .A2(_11012_),
    .ZN(_11053_)
  );
  AND2_X1 _45499_ (
    .A1(_10934_),
    .A2(_11000_),
    .ZN(_11054_)
  );
  AND2_X1 _45500_ (
    .A1(_11053_),
    .A2(_11054_),
    .ZN(_11055_)
  );
  AND2_X1 _45501_ (
    .A1(_11052_),
    .A2(_11055_),
    .ZN(_11056_)
  );
  AND2_X1 _45502_ (
    .A1(_11049_),
    .A2(_11056_),
    .ZN(_11057_)
  );
  AND2_X1 _45503_ (
    .A1(_10970_),
    .A2(_10982_),
    .ZN(_11058_)
  );
  AND2_X1 _45504_ (
    .A1(_10964_),
    .A2(_10976_),
    .ZN(_11059_)
  );
  AND2_X1 _45505_ (
    .A1(_11058_),
    .A2(_11059_),
    .ZN(_11060_)
  );
  AND2_X1 _45506_ (
    .A1(_10862_),
    .A2(_10910_),
    .ZN(_11061_)
  );
  AND2_X1 _45507_ (
    .A1(_10856_),
    .A2(_10904_),
    .ZN(_11062_)
  );
  AND2_X1 _45508_ (
    .A1(_11061_),
    .A2(_11062_),
    .ZN(_11063_)
  );
  AND2_X1 _45509_ (
    .A1(_11060_),
    .A2(_11063_),
    .ZN(_11064_)
  );
  AND2_X1 _45510_ (
    .A1(_10880_),
    .A2(_10952_),
    .ZN(_11065_)
  );
  AND2_X1 _45511_ (
    .A1(_10886_),
    .A2(_10958_),
    .ZN(_11066_)
  );
  AND2_X1 _45512_ (
    .A1(_11065_),
    .A2(_11066_),
    .ZN(_11067_)
  );
  AND2_X1 _45513_ (
    .A1(_10994_),
    .A2(_11024_),
    .ZN(_11068_)
  );
  AND2_X1 _45514_ (
    .A1(_10988_),
    .A2(_11018_),
    .ZN(_11069_)
  );
  AND2_X1 _45515_ (
    .A1(_11068_),
    .A2(_11069_),
    .ZN(_11070_)
  );
  AND2_X1 _45516_ (
    .A1(_11067_),
    .A2(_11070_),
    .ZN(_11071_)
  );
  AND2_X1 _45517_ (
    .A1(_11064_),
    .A2(_11071_),
    .ZN(_11072_)
  );
  AND2_X1 _45518_ (
    .A1(_11057_),
    .A2(_11072_),
    .ZN(_11073_)
  );
  INV_X1 _45519_ (
    .A(_11073_),
    .ZN(_11074_)
  );
  AND2_X1 _45520_ (
    .A1(_21061_),
    .A2(_11074_),
    .ZN(_11075_)
  );
  INV_X1 _45521_ (
    .A(_11075_),
    .ZN(_11076_)
  );
  AND2_X1 _45522_ (
    .A1(_21062_),
    .A2(_11073_),
    .ZN(_11077_)
  );
  INV_X1 _45523_ (
    .A(_11077_),
    .ZN(_11078_)
  );
  AND2_X1 _45524_ (
    .A1(_11076_),
    .A2(_11078_),
    .ZN(_11079_)
  );
  INV_X1 _45525_ (
    .A(_11079_),
    .ZN(_11080_)
  );
  AND2_X1 _45526_ (
    .A1(is_sltiu_bltu_sltu),
    .A2(_10847_),
    .ZN(_11081_)
  );
  INV_X1 _45527_ (
    .A(_11081_),
    .ZN(_11082_)
  );
  AND2_X1 _45528_ (
    .A1(_11080_),
    .A2(_11082_),
    .ZN(_11083_)
  );
  AND2_X1 _45529_ (
    .A1(_10850_),
    .A2(_11083_),
    .ZN(_11084_)
  );
  AND2_X1 _45530_ (
    .A1(_10839_),
    .A2(_11084_),
    .ZN(_11085_)
  );
  AND2_X1 _45531_ (
    .A1(_10837_),
    .A2(_11085_),
    .ZN(_11086_)
  );
  INV_X1 _45532_ (
    .A(_11086_),
    .ZN(_11087_)
  );
  AND2_X1 _45533_ (
    .A1(_22031_),
    .A2(_22054_),
    .ZN(_11088_)
  );
  AND2_X1 _45534_ (
    .A1(_22258_),
    .A2(_11088_),
    .ZN(_11089_)
  );
  AND2_X1 _45535_ (
    .A1(_22252_),
    .A2(_11089_),
    .ZN(_11090_)
  );
  INV_X1 _45536_ (
    .A(_11090_),
    .ZN(_11091_)
  );
  AND2_X1 _45537_ (
    .A1(is_beq_bne_blt_bge_bltu_bgeu),
    .A2(_11090_),
    .ZN(_11092_)
  );
  AND2_X1 _45538_ (
    .A1(_11087_),
    .A2(_11092_),
    .ZN(_11093_)
  );
  INV_X1 _45539_ (
    .A(_11093_),
    .ZN(_11094_)
  );
  AND2_X1 _45540_ (
    .A1(_11087_),
    .A2(_11090_),
    .ZN(_11095_)
  );
  INV_X1 _45541_ (
    .A(_11095_),
    .ZN(_11096_)
  );
  AND2_X1 _45542_ (
    .A1(is_beq_bne_blt_bge_bltu_bgeu),
    .A2(resetn),
    .ZN(_11097_)
  );
  AND2_X1 _45543_ (
    .A1(resetn),
    .A2(_11090_),
    .ZN(_11098_)
  );
  AND2_X1 _45544_ (
    .A1(resetn),
    .A2(_11093_),
    .ZN(_11099_)
  );
  INV_X1 _45545_ (
    .A(_11099_),
    .ZN(_11100_)
  );
  AND2_X1 _45546_ (
    .A1(mem_do_prefetch),
    .A2(_21291_),
    .ZN(_11101_)
  );
  AND2_X1 _45547_ (
    .A1(_22271_),
    .A2(_22537_),
    .ZN(_11102_)
  );
  INV_X1 _45548_ (
    .A(_11102_),
    .ZN(_11103_)
  );
  AND2_X1 _45549_ (
    .A1(_02465_),
    .A2(_11091_),
    .ZN(_11104_)
  );
  INV_X1 _45550_ (
    .A(_11104_),
    .ZN(_11105_)
  );
  AND2_X1 _45551_ (
    .A1(_22262_),
    .A2(_11104_),
    .ZN(_11106_)
  );
  AND2_X1 _45552_ (
    .A1(_04960_),
    .A2(_11106_),
    .ZN(_11107_)
  );
  INV_X1 _45553_ (
    .A(_11107_),
    .ZN(_11108_)
  );
  AND2_X1 _45554_ (
    .A1(_22073_),
    .A2(_04958_),
    .ZN(_11109_)
  );
  INV_X1 _45555_ (
    .A(_11109_),
    .ZN(_11110_)
  );
  AND2_X1 _45556_ (
    .A1(_00027_),
    .A2(_22499_),
    .ZN(_11111_)
  );
  INV_X1 _45557_ (
    .A(_11111_),
    .ZN(_11112_)
  );
  AND2_X1 _45558_ (
    .A1(_22271_),
    .A2(_11112_),
    .ZN(_11113_)
  );
  INV_X1 _45559_ (
    .A(_11113_),
    .ZN(_11114_)
  );
  AND2_X1 _45560_ (
    .A1(_22296_),
    .A2(_11091_),
    .ZN(_11115_)
  );
  AND2_X1 _45561_ (
    .A1(_11114_),
    .A2(_11115_),
    .ZN(_11116_)
  );
  AND2_X1 _45562_ (
    .A1(_11110_),
    .A2(_11116_),
    .ZN(_11117_)
  );
  AND2_X1 _45563_ (
    .A1(_11108_),
    .A2(_11117_),
    .ZN(_11118_)
  );
  AND2_X1 _45564_ (
    .A1(_22271_),
    .A2(_22500_),
    .ZN(_11119_)
  );
  INV_X1 _45565_ (
    .A(_11119_),
    .ZN(_11120_)
  );
  AND2_X1 _45566_ (
    .A1(_11103_),
    .A2(_11118_),
    .ZN(_11121_)
  );
  AND2_X1 _45567_ (
    .A1(resetn),
    .A2(_22073_),
    .ZN(_11122_)
  );
  AND2_X1 _45568_ (
    .A1(_05137_),
    .A2(_11122_),
    .ZN(_11123_)
  );
  INV_X1 _45569_ (
    .A(_11123_),
    .ZN(_11124_)
  );
  AND2_X1 _45570_ (
    .A1(_11121_),
    .A2(_11124_),
    .ZN(_11125_)
  );
  INV_X1 _45571_ (
    .A(_11125_),
    .ZN(_11126_)
  );
  AND2_X1 _45572_ (
    .A1(_22283_),
    .A2(_04967_),
    .ZN(_11127_)
  );
  INV_X1 _45573_ (
    .A(_11127_),
    .ZN(_11128_)
  );
  AND2_X1 _45574_ (
    .A1(mem_do_prefetch),
    .A2(_11128_),
    .ZN(_11129_)
  );
  INV_X1 _45575_ (
    .A(_11129_),
    .ZN(_11130_)
  );
  AND2_X1 _45576_ (
    .A1(_21261_),
    .A2(decoder_trigger),
    .ZN(_11131_)
  );
  INV_X1 _45577_ (
    .A(_11131_),
    .ZN(_11132_)
  );
  AND2_X1 _45578_ (
    .A1(_02464_),
    .A2(_11132_),
    .ZN(_11133_)
  );
  INV_X1 _45579_ (
    .A(_11133_),
    .ZN(_11134_)
  );
  AND2_X1 _45580_ (
    .A1(_22067_),
    .A2(_22146_),
    .ZN(_11135_)
  );
  INV_X1 _45581_ (
    .A(_11135_),
    .ZN(_11136_)
  );
  AND2_X1 _45582_ (
    .A1(_11133_),
    .A2(_11136_),
    .ZN(_11137_)
  );
  INV_X1 _45583_ (
    .A(_11137_),
    .ZN(_11138_)
  );
  AND2_X1 _45584_ (
    .A1(is_lb_lh_lw_lbu_lhu),
    .A2(_22271_),
    .ZN(_11139_)
  );
  AND2_X1 _45585_ (
    .A1(_22538_),
    .A2(_11139_),
    .ZN(_11140_)
  );
  INV_X1 _45586_ (
    .A(_11140_),
    .ZN(_11141_)
  );
  AND2_X1 _45587_ (
    .A1(_11130_),
    .A2(_11141_),
    .ZN(_11142_)
  );
  AND2_X1 _45588_ (
    .A1(is_sb_sh_sw),
    .A2(_05841_),
    .ZN(_11143_)
  );
  INV_X1 _45589_ (
    .A(_11143_),
    .ZN(_11144_)
  );
  AND2_X1 _45590_ (
    .A1(_05841_),
    .A2(_11101_),
    .ZN(_11145_)
  );
  INV_X1 _45591_ (
    .A(_11145_),
    .ZN(_11146_)
  );
  AND2_X1 _45592_ (
    .A1(_11144_),
    .A2(_11146_),
    .ZN(_11147_)
  );
  AND2_X1 _45593_ (
    .A1(_11125_),
    .A2(_11138_),
    .ZN(_11148_)
  );
  AND2_X1 _45594_ (
    .A1(_11147_),
    .A2(_11148_),
    .ZN(_11149_)
  );
  AND2_X1 _45595_ (
    .A1(_11142_),
    .A2(_11149_),
    .ZN(_11150_)
  );
  INV_X1 _45596_ (
    .A(_11150_),
    .ZN(_11151_)
  );
  AND2_X1 _45597_ (
    .A1(_21070_),
    .A2(_11126_),
    .ZN(_11152_)
  );
  INV_X1 _45598_ (
    .A(_11152_),
    .ZN(_11153_)
  );
  AND2_X1 _45599_ (
    .A1(_10521_),
    .A2(_11153_),
    .ZN(_11154_)
  );
  AND2_X1 _45600_ (
    .A1(_11151_),
    .A2(_11154_),
    .ZN(_11155_)
  );
  INV_X1 _45601_ (
    .A(_11155_),
    .ZN(_11156_)
  );
  AND2_X1 _45602_ (
    .A1(_11100_),
    .A2(_11156_),
    .ZN(_11157_)
  );
  INV_X1 _45603_ (
    .A(_11157_),
    .ZN(_00339_)
  );
  AND2_X1 _45604_ (
    .A1(_00034_),
    .A2(_22323_),
    .ZN(_11158_)
  );
  INV_X1 _45605_ (
    .A(_11158_),
    .ZN(_11159_)
  );
  AND2_X1 _45606_ (
    .A1(mem_do_rdata),
    .A2(_10521_),
    .ZN(_11160_)
  );
  INV_X1 _45607_ (
    .A(_11160_),
    .ZN(_11161_)
  );
  AND2_X1 _45608_ (
    .A1(resetn),
    .A2(_00034_),
    .ZN(_11162_)
  );
  AND2_X1 _45609_ (
    .A1(_22323_),
    .A2(_11162_),
    .ZN(_11163_)
  );
  INV_X1 _45610_ (
    .A(_11163_),
    .ZN(_11164_)
  );
  AND2_X1 _45611_ (
    .A1(_11161_),
    .A2(_11164_),
    .ZN(_11165_)
  );
  INV_X1 _45612_ (
    .A(_11165_),
    .ZN(_00340_)
  );
  AND2_X1 _45613_ (
    .A1(mem_do_wdata),
    .A2(_10521_),
    .ZN(_11166_)
  );
  INV_X1 _45614_ (
    .A(_11166_),
    .ZN(_11167_)
  );
  AND2_X1 _45615_ (
    .A1(resetn),
    .A2(_00045_),
    .ZN(_11168_)
  );
  AND2_X1 _45616_ (
    .A1(_22320_),
    .A2(_11168_),
    .ZN(_11169_)
  );
  INV_X1 _45617_ (
    .A(_11169_),
    .ZN(_11170_)
  );
  AND2_X1 _45618_ (
    .A1(_11167_),
    .A2(_11170_),
    .ZN(_11171_)
  );
  INV_X1 _45619_ (
    .A(_11171_),
    .ZN(_00341_)
  );
  AND2_X1 _45620_ (
    .A1(_21264_),
    .A2(_21267_),
    .ZN(_11172_)
  );
  INV_X1 _45621_ (
    .A(_11172_),
    .ZN(_11173_)
  );
  AND2_X1 _45622_ (
    .A1(_21263_),
    .A2(_21266_),
    .ZN(_11174_)
  );
  INV_X1 _45623_ (
    .A(_11174_),
    .ZN(_11175_)
  );
  AND2_X1 _45624_ (
    .A1(_21265_),
    .A2(_11174_),
    .ZN(_11176_)
  );
  AND2_X1 _45625_ (
    .A1(_11172_),
    .A2(_11176_),
    .ZN(_11177_)
  );
  AND2_X1 _45626_ (
    .A1(_22556_),
    .A2(_11177_),
    .ZN(_11178_)
  );
  INV_X1 _45627_ (
    .A(_11178_),
    .ZN(_11179_)
  );
  AND2_X1 _45628_ (
    .A1(_21269_),
    .A2(_22530_),
    .ZN(_11180_)
  );
  AND2_X1 _45629_ (
    .A1(_22554_),
    .A2(_11180_),
    .ZN(_11181_)
  );
  INV_X1 _45630_ (
    .A(_11181_),
    .ZN(_11182_)
  );
  AND2_X1 _45631_ (
    .A1(_22326_),
    .A2(_02465_),
    .ZN(_11183_)
  );
  INV_X1 _45632_ (
    .A(_11183_),
    .ZN(_11184_)
  );
  AND2_X1 _45633_ (
    .A1(_11182_),
    .A2(_11184_),
    .ZN(_11185_)
  );
  AND2_X1 _45634_ (
    .A1(_11179_),
    .A2(_11185_),
    .ZN(_11186_)
  );
  AND2_X1 _45635_ (
    .A1(_22332_),
    .A2(_11186_),
    .ZN(_11187_)
  );
  INV_X1 _45636_ (
    .A(_11187_),
    .ZN(_11188_)
  );
  AND2_X1 _45637_ (
    .A1(instr_sh),
    .A2(_22554_),
    .ZN(_11189_)
  );
  INV_X1 _45638_ (
    .A(_11189_),
    .ZN(_11190_)
  );
  AND2_X1 _45639_ (
    .A1(_22556_),
    .A2(_11173_),
    .ZN(_11191_)
  );
  INV_X1 _45640_ (
    .A(_11191_),
    .ZN(_11192_)
  );
  AND2_X1 _45641_ (
    .A1(_11190_),
    .A2(_11192_),
    .ZN(_11193_)
  );
  AND2_X1 _45642_ (
    .A1(_21252_),
    .A2(_11188_),
    .ZN(_11194_)
  );
  INV_X1 _45643_ (
    .A(_11194_),
    .ZN(_11195_)
  );
  AND2_X1 _45644_ (
    .A1(_11187_),
    .A2(_11193_),
    .ZN(_11196_)
  );
  INV_X1 _45645_ (
    .A(_11196_),
    .ZN(_11197_)
  );
  AND2_X1 _45646_ (
    .A1(_11195_),
    .A2(_11197_),
    .ZN(_00342_)
  );
  AND2_X1 _45647_ (
    .A1(_22556_),
    .A2(_11175_),
    .ZN(_11198_)
  );
  INV_X1 _45648_ (
    .A(_11198_),
    .ZN(_11199_)
  );
  AND2_X1 _45649_ (
    .A1(instr_sb),
    .A2(_22554_),
    .ZN(_11200_)
  );
  INV_X1 _45650_ (
    .A(_11200_),
    .ZN(_11201_)
  );
  AND2_X1 _45651_ (
    .A1(_11199_),
    .A2(_11201_),
    .ZN(_11202_)
  );
  AND2_X1 _45652_ (
    .A1(_21253_),
    .A2(_11188_),
    .ZN(_11203_)
  );
  INV_X1 _45653_ (
    .A(_11203_),
    .ZN(_11204_)
  );
  AND2_X1 _45654_ (
    .A1(_11187_),
    .A2(_11202_),
    .ZN(_11205_)
  );
  INV_X1 _45655_ (
    .A(_11205_),
    .ZN(_11206_)
  );
  AND2_X1 _45656_ (
    .A1(_11204_),
    .A2(_11206_),
    .ZN(_00343_)
  );
  AND2_X1 _45657_ (
    .A1(_22272_),
    .A2(_11105_),
    .ZN(_11207_)
  );
  INV_X1 _45658_ (
    .A(_11207_),
    .ZN(_11208_)
  );
  AND2_X1 _45659_ (
    .A1(_22263_),
    .A2(_11104_),
    .ZN(_11209_)
  );
  INV_X1 _45660_ (
    .A(_11209_),
    .ZN(_11210_)
  );
  AND2_X1 _45661_ (
    .A1(_22272_),
    .A2(_11210_),
    .ZN(_11211_)
  );
  INV_X1 _45662_ (
    .A(_11211_),
    .ZN(_11212_)
  );
  AND2_X1 _45663_ (
    .A1(_11120_),
    .A2(_11212_),
    .ZN(_11213_)
  );
  INV_X1 _45664_ (
    .A(_11213_),
    .ZN(_11214_)
  );
  AND2_X1 _45665_ (
    .A1(_04959_),
    .A2(_11214_),
    .ZN(_11215_)
  );
  INV_X1 _45666_ (
    .A(_11215_),
    .ZN(_11216_)
  );
  AND2_X1 _45667_ (
    .A1(_21039_),
    .A2(_11090_),
    .ZN(_11217_)
  );
  INV_X1 _45668_ (
    .A(_11217_),
    .ZN(_11218_)
  );
  AND2_X1 _45669_ (
    .A1(_22263_),
    .A2(_11218_),
    .ZN(_11219_)
  );
  AND2_X1 _45670_ (
    .A1(_11120_),
    .A2(_11219_),
    .ZN(_11220_)
  );
  AND2_X1 _45671_ (
    .A1(_11215_),
    .A2(_11220_),
    .ZN(_11221_)
  );
  AND2_X1 _45672_ (
    .A1(_11096_),
    .A2(_11221_),
    .ZN(_11222_)
  );
  INV_X1 _45673_ (
    .A(_11222_),
    .ZN(_11223_)
  );
  AND2_X1 _45674_ (
    .A1(_21068_),
    .A2(_11216_),
    .ZN(_11224_)
  );
  INV_X1 _45675_ (
    .A(_11224_),
    .ZN(_11225_)
  );
  AND2_X1 _45676_ (
    .A1(resetn),
    .A2(_11225_),
    .ZN(_11226_)
  );
  AND2_X1 _45677_ (
    .A1(_11223_),
    .A2(_11226_),
    .ZN(_00344_)
  );
  AND2_X1 _45678_ (
    .A1(_22072_),
    .A2(_11090_),
    .ZN(_11227_)
  );
  INV_X1 _45679_ (
    .A(_11227_),
    .ZN(_11228_)
  );
  AND2_X1 _45680_ (
    .A1(_11105_),
    .A2(_11228_),
    .ZN(_11229_)
  );
  INV_X1 _45681_ (
    .A(_11229_),
    .ZN(_11230_)
  );
  AND2_X1 _45682_ (
    .A1(latched_stalu),
    .A2(_11230_),
    .ZN(_11231_)
  );
  INV_X1 _45683_ (
    .A(_11231_),
    .ZN(_11232_)
  );
  AND2_X1 _45684_ (
    .A1(_00047_),
    .A2(_11217_),
    .ZN(_11233_)
  );
  INV_X1 _45685_ (
    .A(_11233_),
    .ZN(_11234_)
  );
  AND2_X1 _45686_ (
    .A1(_11232_),
    .A2(_11234_),
    .ZN(_11235_)
  );
  INV_X1 _45687_ (
    .A(_11235_),
    .ZN(_11236_)
  );
  AND2_X1 _45688_ (
    .A1(resetn),
    .A2(_11236_),
    .ZN(_00345_)
  );
  AND2_X1 _45689_ (
    .A1(instr_jalr),
    .A2(_11217_),
    .ZN(_11237_)
  );
  INV_X1 _45690_ (
    .A(_11237_),
    .ZN(_11238_)
  );
  AND2_X1 _45691_ (
    .A1(instr_jal),
    .A2(_02466_),
    .ZN(_11239_)
  );
  INV_X1 _45692_ (
    .A(_11239_),
    .ZN(_11240_)
  );
  AND2_X1 _45693_ (
    .A1(_11238_),
    .A2(_11240_),
    .ZN(_11241_)
  );
  AND2_X1 _45694_ (
    .A1(_11207_),
    .A2(_11241_),
    .ZN(_11242_)
  );
  AND2_X1 _45695_ (
    .A1(_11094_),
    .A2(_11242_),
    .ZN(_11243_)
  );
  INV_X1 _45696_ (
    .A(_11243_),
    .ZN(_11244_)
  );
  AND2_X1 _45697_ (
    .A1(_21066_),
    .A2(_11208_),
    .ZN(_11245_)
  );
  INV_X1 _45698_ (
    .A(_11245_),
    .ZN(_11246_)
  );
  AND2_X1 _45699_ (
    .A1(resetn),
    .A2(_11246_),
    .ZN(_11247_)
  );
  AND2_X1 _45700_ (
    .A1(_11244_),
    .A2(_11247_),
    .ZN(_00346_)
  );
  AND2_X1 _45701_ (
    .A1(_22257_),
    .A2(_02464_),
    .ZN(_11248_)
  );
  INV_X1 _45702_ (
    .A(_11248_),
    .ZN(_11249_)
  );
  AND2_X1 _45703_ (
    .A1(_11159_),
    .A2(_11249_),
    .ZN(_11250_)
  );
  INV_X1 _45704_ (
    .A(_11250_),
    .ZN(_11251_)
  );
  AND2_X1 _45705_ (
    .A1(is_lbu_lhu_lw),
    .A2(_22556_),
    .ZN(_11252_)
  );
  INV_X1 _45706_ (
    .A(_11252_),
    .ZN(_11253_)
  );
  AND2_X1 _45707_ (
    .A1(_21065_),
    .A2(_11250_),
    .ZN(_11254_)
  );
  INV_X1 _45708_ (
    .A(_11254_),
    .ZN(_11255_)
  );
  AND2_X1 _45709_ (
    .A1(_11251_),
    .A2(_11253_),
    .ZN(_11256_)
  );
  INV_X1 _45710_ (
    .A(_11256_),
    .ZN(_11257_)
  );
  AND2_X1 _45711_ (
    .A1(resetn),
    .A2(_11257_),
    .ZN(_11258_)
  );
  AND2_X1 _45712_ (
    .A1(_11255_),
    .A2(_11258_),
    .ZN(_00347_)
  );
  AND2_X1 _45713_ (
    .A1(instr_lh),
    .A2(_22556_),
    .ZN(_11259_)
  );
  INV_X1 _45714_ (
    .A(_11259_),
    .ZN(_11260_)
  );
  AND2_X1 _45715_ (
    .A1(_21064_),
    .A2(_11250_),
    .ZN(_11261_)
  );
  INV_X1 _45716_ (
    .A(_11261_),
    .ZN(_11262_)
  );
  AND2_X1 _45717_ (
    .A1(_11251_),
    .A2(_11260_),
    .ZN(_11263_)
  );
  INV_X1 _45718_ (
    .A(_11263_),
    .ZN(_11264_)
  );
  AND2_X1 _45719_ (
    .A1(resetn),
    .A2(_11264_),
    .ZN(_11265_)
  );
  AND2_X1 _45720_ (
    .A1(_11262_),
    .A2(_11265_),
    .ZN(_00348_)
  );
  AND2_X1 _45721_ (
    .A1(instr_lb),
    .A2(_22556_),
    .ZN(_11266_)
  );
  INV_X1 _45722_ (
    .A(_11266_),
    .ZN(_11267_)
  );
  AND2_X1 _45723_ (
    .A1(_21063_),
    .A2(_11250_),
    .ZN(_11268_)
  );
  INV_X1 _45724_ (
    .A(_11268_),
    .ZN(_11269_)
  );
  AND2_X1 _45725_ (
    .A1(_11251_),
    .A2(_11267_),
    .ZN(_11270_)
  );
  INV_X1 _45726_ (
    .A(_11270_),
    .ZN(_11271_)
  );
  AND2_X1 _45727_ (
    .A1(resetn),
    .A2(_11271_),
    .ZN(_11272_)
  );
  AND2_X1 _45728_ (
    .A1(_11269_),
    .A2(_11272_),
    .ZN(_00349_)
  );
  AND2_X1 _45729_ (
    .A1(resetn),
    .A2(_11218_),
    .ZN(_11273_)
  );
  AND2_X1 _45730_ (
    .A1(_11207_),
    .A2(_11273_),
    .ZN(_11274_)
  );
  INV_X1 _45731_ (
    .A(_11274_),
    .ZN(_11275_)
  );
  AND2_X1 _45732_ (
    .A1(decoded_rd[0]),
    .A2(_02464_),
    .ZN(_11276_)
  );
  AND2_X1 _45733_ (
    .A1(latched_rd[0]),
    .A2(_11275_),
    .ZN(_11277_)
  );
  INV_X1 _45734_ (
    .A(_11277_),
    .ZN(_11278_)
  );
  AND2_X1 _45735_ (
    .A1(_11274_),
    .A2(_11276_),
    .ZN(_11279_)
  );
  INV_X1 _45736_ (
    .A(_11279_),
    .ZN(_11280_)
  );
  AND2_X1 _45737_ (
    .A1(_11278_),
    .A2(_11280_),
    .ZN(_11281_)
  );
  INV_X1 _45738_ (
    .A(_11281_),
    .ZN(_00350_)
  );
  AND2_X1 _45739_ (
    .A1(decoded_rd[1]),
    .A2(_02464_),
    .ZN(_11282_)
  );
  AND2_X1 _45740_ (
    .A1(latched_rd[1]),
    .A2(_11275_),
    .ZN(_11283_)
  );
  INV_X1 _45741_ (
    .A(_11283_),
    .ZN(_11284_)
  );
  AND2_X1 _45742_ (
    .A1(_11274_),
    .A2(_11282_),
    .ZN(_11285_)
  );
  INV_X1 _45743_ (
    .A(_11285_),
    .ZN(_11286_)
  );
  AND2_X1 _45744_ (
    .A1(_11284_),
    .A2(_11286_),
    .ZN(_11287_)
  );
  INV_X1 _45745_ (
    .A(_11287_),
    .ZN(_00351_)
  );
  AND2_X1 _45746_ (
    .A1(decoded_rd[2]),
    .A2(_02464_),
    .ZN(_11288_)
  );
  AND2_X1 _45747_ (
    .A1(latched_rd[2]),
    .A2(_11275_),
    .ZN(_11289_)
  );
  INV_X1 _45748_ (
    .A(_11289_),
    .ZN(_11290_)
  );
  AND2_X1 _45749_ (
    .A1(_11274_),
    .A2(_11288_),
    .ZN(_11291_)
  );
  INV_X1 _45750_ (
    .A(_11291_),
    .ZN(_11292_)
  );
  AND2_X1 _45751_ (
    .A1(_11290_),
    .A2(_11292_),
    .ZN(_11293_)
  );
  INV_X1 _45752_ (
    .A(_11293_),
    .ZN(_00352_)
  );
  AND2_X1 _45753_ (
    .A1(decoded_rd[3]),
    .A2(_02464_),
    .ZN(_11294_)
  );
  AND2_X1 _45754_ (
    .A1(latched_rd[3]),
    .A2(_11275_),
    .ZN(_11295_)
  );
  INV_X1 _45755_ (
    .A(_11295_),
    .ZN(_11296_)
  );
  AND2_X1 _45756_ (
    .A1(_11274_),
    .A2(_11294_),
    .ZN(_11297_)
  );
  INV_X1 _45757_ (
    .A(_11297_),
    .ZN(_11298_)
  );
  AND2_X1 _45758_ (
    .A1(_11296_),
    .A2(_11298_),
    .ZN(_11299_)
  );
  INV_X1 _45759_ (
    .A(_11299_),
    .ZN(_00353_)
  );
  AND2_X1 _45760_ (
    .A1(decoded_rd[4]),
    .A2(_02464_),
    .ZN(_11300_)
  );
  AND2_X1 _45761_ (
    .A1(latched_rd[4]),
    .A2(_11275_),
    .ZN(_11301_)
  );
  INV_X1 _45762_ (
    .A(_11301_),
    .ZN(_11302_)
  );
  AND2_X1 _45763_ (
    .A1(_11274_),
    .A2(_11300_),
    .ZN(_11303_)
  );
  INV_X1 _45764_ (
    .A(_11303_),
    .ZN(_11304_)
  );
  AND2_X1 _45765_ (
    .A1(_11302_),
    .A2(_11304_),
    .ZN(_11305_)
  );
  INV_X1 _45766_ (
    .A(_11305_),
    .ZN(_00354_)
  );
  AND2_X1 _45767_ (
    .A1(mem_do_rinst),
    .A2(_22317_),
    .ZN(_11306_)
  );
  INV_X1 _45768_ (
    .A(_11306_),
    .ZN(_11307_)
  );
  AND2_X1 _45769_ (
    .A1(_21350_),
    .A2(_22308_),
    .ZN(_11308_)
  );
  INV_X1 _45770_ (
    .A(_11308_),
    .ZN(_11309_)
  );
  AND2_X1 _45771_ (
    .A1(_21351_),
    .A2(_22307_),
    .ZN(_11310_)
  );
  INV_X1 _45772_ (
    .A(_11310_),
    .ZN(_11311_)
  );
  AND2_X1 _45773_ (
    .A1(_11309_),
    .A2(_11311_),
    .ZN(_00488_)
  );
  AND2_X1 _45774_ (
    .A1(_21352_),
    .A2(_22308_),
    .ZN(_11312_)
  );
  INV_X1 _45775_ (
    .A(_11312_),
    .ZN(_11313_)
  );
  AND2_X1 _45776_ (
    .A1(_21353_),
    .A2(_22307_),
    .ZN(_11314_)
  );
  INV_X1 _45777_ (
    .A(_11314_),
    .ZN(_11315_)
  );
  AND2_X1 _45778_ (
    .A1(_11313_),
    .A2(_11315_),
    .ZN(_00489_)
  );
  AND2_X1 _45779_ (
    .A1(_00488_),
    .A2(_00489_),
    .ZN(_11316_)
  );
  AND2_X1 _45780_ (
    .A1(_21354_),
    .A2(_22308_),
    .ZN(_11317_)
  );
  INV_X1 _45781_ (
    .A(_11317_),
    .ZN(_11318_)
  );
  AND2_X1 _45782_ (
    .A1(_21355_),
    .A2(_22307_),
    .ZN(_11319_)
  );
  INV_X1 _45783_ (
    .A(_11319_),
    .ZN(_11320_)
  );
  AND2_X1 _45784_ (
    .A1(_11318_),
    .A2(_11320_),
    .ZN(_00490_)
  );
  INV_X1 _45785_ (
    .A(_00490_),
    .ZN(_11321_)
  );
  AND2_X1 _45786_ (
    .A1(_11316_),
    .A2(_00490_),
    .ZN(_11322_)
  );
  AND2_X1 _45787_ (
    .A1(mem_rdata[3]),
    .A2(_22307_),
    .ZN(_11323_)
  );
  INV_X1 _45788_ (
    .A(_11323_),
    .ZN(_11324_)
  );
  AND2_X1 _45789_ (
    .A1(mem_rdata_q[3]),
    .A2(_22308_),
    .ZN(_11325_)
  );
  INV_X1 _45790_ (
    .A(_11325_),
    .ZN(_11326_)
  );
  AND2_X1 _45791_ (
    .A1(_11324_),
    .A2(_11326_),
    .ZN(_11327_)
  );
  INV_X1 _45792_ (
    .A(_11327_),
    .ZN(_00491_)
  );
  AND2_X1 _45793_ (
    .A1(_11322_),
    .A2(_11327_),
    .ZN(_11328_)
  );
  AND2_X1 _45794_ (
    .A1(mem_rdata[6]),
    .A2(_22307_),
    .ZN(_11329_)
  );
  INV_X1 _45795_ (
    .A(_11329_),
    .ZN(_11330_)
  );
  AND2_X1 _45796_ (
    .A1(mem_rdata_q[6]),
    .A2(_22308_),
    .ZN(_11331_)
  );
  INV_X1 _45797_ (
    .A(_11331_),
    .ZN(_11332_)
  );
  AND2_X1 _45798_ (
    .A1(_11330_),
    .A2(_11332_),
    .ZN(_11333_)
  );
  INV_X1 _45799_ (
    .A(_11333_),
    .ZN(_00494_)
  );
  AND2_X1 _45800_ (
    .A1(mem_rdata[4]),
    .A2(_22307_),
    .ZN(_11334_)
  );
  INV_X1 _45801_ (
    .A(_11334_),
    .ZN(_11335_)
  );
  AND2_X1 _45802_ (
    .A1(mem_rdata_q[4]),
    .A2(_22308_),
    .ZN(_11336_)
  );
  INV_X1 _45803_ (
    .A(_11336_),
    .ZN(_11337_)
  );
  AND2_X1 _45804_ (
    .A1(_11335_),
    .A2(_11337_),
    .ZN(_11338_)
  );
  INV_X1 _45805_ (
    .A(_11338_),
    .ZN(_00492_)
  );
  AND2_X1 _45806_ (
    .A1(_11333_),
    .A2(_00492_),
    .ZN(_11339_)
  );
  AND2_X1 _45807_ (
    .A1(mem_rdata[5]),
    .A2(_22307_),
    .ZN(_11340_)
  );
  INV_X1 _45808_ (
    .A(_11340_),
    .ZN(_11341_)
  );
  AND2_X1 _45809_ (
    .A1(mem_rdata_q[5]),
    .A2(_22308_),
    .ZN(_11342_)
  );
  INV_X1 _45810_ (
    .A(_11342_),
    .ZN(_11343_)
  );
  AND2_X1 _45811_ (
    .A1(_11341_),
    .A2(_11343_),
    .ZN(_11344_)
  );
  INV_X1 _45812_ (
    .A(_11344_),
    .ZN(_00493_)
  );
  AND2_X1 _45813_ (
    .A1(_11339_),
    .A2(_00493_),
    .ZN(_11345_)
  );
  AND2_X1 _45814_ (
    .A1(_11328_),
    .A2(_11345_),
    .ZN(_11346_)
  );
  AND2_X1 _45815_ (
    .A1(_11306_),
    .A2(_11346_),
    .ZN(_11347_)
  );
  INV_X1 _45816_ (
    .A(_11347_),
    .ZN(_11348_)
  );
  AND2_X1 _45817_ (
    .A1(instr_lui),
    .A2(_11307_),
    .ZN(_11349_)
  );
  INV_X1 _45818_ (
    .A(_11349_),
    .ZN(_11350_)
  );
  AND2_X1 _45819_ (
    .A1(_11348_),
    .A2(_11350_),
    .ZN(_11351_)
  );
  INV_X1 _45820_ (
    .A(_11351_),
    .ZN(_00355_)
  );
  AND2_X1 _45821_ (
    .A1(_11339_),
    .A2(_11344_),
    .ZN(_11352_)
  );
  AND2_X1 _45822_ (
    .A1(_11328_),
    .A2(_11352_),
    .ZN(_11353_)
  );
  AND2_X1 _45823_ (
    .A1(_11306_),
    .A2(_11353_),
    .ZN(_11354_)
  );
  INV_X1 _45824_ (
    .A(_11354_),
    .ZN(_11355_)
  );
  AND2_X1 _45825_ (
    .A1(instr_auipc),
    .A2(_11307_),
    .ZN(_11356_)
  );
  INV_X1 _45826_ (
    .A(_11356_),
    .ZN(_11357_)
  );
  AND2_X1 _45827_ (
    .A1(_11355_),
    .A2(_11357_),
    .ZN(_11358_)
  );
  INV_X1 _45828_ (
    .A(_11358_),
    .ZN(_00356_)
  );
  AND2_X1 _45829_ (
    .A1(_11338_),
    .A2(_00493_),
    .ZN(_11359_)
  );
  AND2_X1 _45830_ (
    .A1(_00494_),
    .A2(_11359_),
    .ZN(_11360_)
  );
  AND2_X1 _45831_ (
    .A1(_11322_),
    .A2(_00491_),
    .ZN(_11361_)
  );
  AND2_X1 _45832_ (
    .A1(_11360_),
    .A2(_11361_),
    .ZN(_11362_)
  );
  AND2_X1 _45833_ (
    .A1(instr_jal),
    .A2(_11307_),
    .ZN(_11363_)
  );
  INV_X1 _45834_ (
    .A(_11363_),
    .ZN(_11364_)
  );
  AND2_X1 _45835_ (
    .A1(_11306_),
    .A2(_11362_),
    .ZN(_11365_)
  );
  INV_X1 _45836_ (
    .A(_11365_),
    .ZN(_11366_)
  );
  AND2_X1 _45837_ (
    .A1(_11364_),
    .A2(_11366_),
    .ZN(_11367_)
  );
  INV_X1 _45838_ (
    .A(_11367_),
    .ZN(_00357_)
  );
  AND2_X1 _45839_ (
    .A1(resetn),
    .A2(_02901_),
    .ZN(_11368_)
  );
  AND2_X1 _45840_ (
    .A1(instr_beq),
    .A2(_11368_),
    .ZN(_11369_)
  );
  INV_X1 _45841_ (
    .A(_11369_),
    .ZN(_11370_)
  );
  AND2_X1 _45842_ (
    .A1(_21232_),
    .A2(_21233_),
    .ZN(_11371_)
  );
  AND2_X1 _45843_ (
    .A1(_21234_),
    .A2(_11371_),
    .ZN(_11372_)
  );
  INV_X1 _45844_ (
    .A(_11372_),
    .ZN(_11373_)
  );
  AND2_X1 _45845_ (
    .A1(_02900_),
    .A2(_11097_),
    .ZN(_11374_)
  );
  AND2_X1 _45846_ (
    .A1(_11372_),
    .A2(_11374_),
    .ZN(_11375_)
  );
  INV_X1 _45847_ (
    .A(_11375_),
    .ZN(_11376_)
  );
  AND2_X1 _45848_ (
    .A1(_11370_),
    .A2(_11376_),
    .ZN(_11377_)
  );
  INV_X1 _45849_ (
    .A(_11377_),
    .ZN(_00358_)
  );
  AND2_X1 _45850_ (
    .A1(_21233_),
    .A2(_22051_),
    .ZN(_11378_)
  );
  AND2_X1 _45851_ (
    .A1(_21234_),
    .A2(_11378_),
    .ZN(_11379_)
  );
  AND2_X1 _45852_ (
    .A1(_11374_),
    .A2(_11379_),
    .ZN(_11380_)
  );
  INV_X1 _45853_ (
    .A(_11380_),
    .ZN(_11381_)
  );
  AND2_X1 _45854_ (
    .A1(instr_bne),
    .A2(_11368_),
    .ZN(_11382_)
  );
  INV_X1 _45855_ (
    .A(_11382_),
    .ZN(_11383_)
  );
  AND2_X1 _45856_ (
    .A1(_11381_),
    .A2(_11383_),
    .ZN(_11384_)
  );
  INV_X1 _45857_ (
    .A(_11384_),
    .ZN(_00359_)
  );
  AND2_X1 _45858_ (
    .A1(_22050_),
    .A2(_11371_),
    .ZN(_11385_)
  );
  INV_X1 _45859_ (
    .A(_11385_),
    .ZN(_11386_)
  );
  AND2_X1 _45860_ (
    .A1(_11374_),
    .A2(_11385_),
    .ZN(_11387_)
  );
  INV_X1 _45861_ (
    .A(_11387_),
    .ZN(_11388_)
  );
  AND2_X1 _45862_ (
    .A1(instr_blt),
    .A2(_11368_),
    .ZN(_11389_)
  );
  INV_X1 _45863_ (
    .A(_11389_),
    .ZN(_11390_)
  );
  AND2_X1 _45864_ (
    .A1(_11388_),
    .A2(_11390_),
    .ZN(_11391_)
  );
  INV_X1 _45865_ (
    .A(_11391_),
    .ZN(_00360_)
  );
  AND2_X1 _45866_ (
    .A1(_22050_),
    .A2(_11378_),
    .ZN(_11392_)
  );
  INV_X1 _45867_ (
    .A(_11392_),
    .ZN(_11393_)
  );
  AND2_X1 _45868_ (
    .A1(_11374_),
    .A2(_11392_),
    .ZN(_11394_)
  );
  INV_X1 _45869_ (
    .A(_11394_),
    .ZN(_11395_)
  );
  AND2_X1 _45870_ (
    .A1(instr_bge),
    .A2(_11368_),
    .ZN(_11396_)
  );
  INV_X1 _45871_ (
    .A(_11396_),
    .ZN(_11397_)
  );
  AND2_X1 _45872_ (
    .A1(_11395_),
    .A2(_11397_),
    .ZN(_11398_)
  );
  INV_X1 _45873_ (
    .A(_11398_),
    .ZN(_00361_)
  );
  AND2_X1 _45874_ (
    .A1(_22050_),
    .A2(_02904_),
    .ZN(_11399_)
  );
  INV_X1 _45875_ (
    .A(_11399_),
    .ZN(_11400_)
  );
  AND2_X1 _45876_ (
    .A1(_11374_),
    .A2(_11399_),
    .ZN(_11401_)
  );
  INV_X1 _45877_ (
    .A(_11401_),
    .ZN(_11402_)
  );
  AND2_X1 _45878_ (
    .A1(instr_bltu),
    .A2(_11368_),
    .ZN(_11403_)
  );
  INV_X1 _45879_ (
    .A(_11403_),
    .ZN(_11404_)
  );
  AND2_X1 _45880_ (
    .A1(_11402_),
    .A2(_11404_),
    .ZN(_11405_)
  );
  INV_X1 _45881_ (
    .A(_11405_),
    .ZN(_00362_)
  );
  AND2_X1 _45882_ (
    .A1(_22051_),
    .A2(_22052_),
    .ZN(_11406_)
  );
  AND2_X1 _45883_ (
    .A1(_22050_),
    .A2(_11406_),
    .ZN(_11407_)
  );
  INV_X1 _45884_ (
    .A(_11407_),
    .ZN(_11408_)
  );
  AND2_X1 _45885_ (
    .A1(_11374_),
    .A2(_11407_),
    .ZN(_11409_)
  );
  INV_X1 _45886_ (
    .A(_11409_),
    .ZN(_11410_)
  );
  AND2_X1 _45887_ (
    .A1(instr_bgeu),
    .A2(_11368_),
    .ZN(_11411_)
  );
  INV_X1 _45888_ (
    .A(_11411_),
    .ZN(_11412_)
  );
  AND2_X1 _45889_ (
    .A1(_11410_),
    .A2(_11412_),
    .ZN(_11413_)
  );
  INV_X1 _45890_ (
    .A(_11413_),
    .ZN(_00363_)
  );
  AND2_X1 _45891_ (
    .A1(instr_jalr),
    .A2(_11307_),
    .ZN(_11414_)
  );
  INV_X1 _45892_ (
    .A(_11414_),
    .ZN(_11415_)
  );
  AND2_X1 _45893_ (
    .A1(_10421_),
    .A2(_11306_),
    .ZN(_11416_)
  );
  INV_X1 _45894_ (
    .A(_11416_),
    .ZN(_11417_)
  );
  AND2_X1 _45895_ (
    .A1(_10426_),
    .A2(_10431_),
    .ZN(_11418_)
  );
  AND2_X1 _45896_ (
    .A1(_11360_),
    .A2(_11418_),
    .ZN(_11419_)
  );
  AND2_X1 _45897_ (
    .A1(_11328_),
    .A2(_11419_),
    .ZN(_11420_)
  );
  AND2_X1 _45898_ (
    .A1(_11416_),
    .A2(_11420_),
    .ZN(_11421_)
  );
  INV_X1 _45899_ (
    .A(_11421_),
    .ZN(_11422_)
  );
  AND2_X1 _45900_ (
    .A1(_11415_),
    .A2(_11422_),
    .ZN(_11423_)
  );
  INV_X1 _45901_ (
    .A(_11423_),
    .ZN(_00364_)
  );
  AND2_X1 _45902_ (
    .A1(instr_lb),
    .A2(_02901_),
    .ZN(_11424_)
  );
  INV_X1 _45903_ (
    .A(_11424_),
    .ZN(_11425_)
  );
  AND2_X1 _45904_ (
    .A1(is_lb_lh_lw_lbu_lhu),
    .A2(_02900_),
    .ZN(_11426_)
  );
  AND2_X1 _45905_ (
    .A1(_11372_),
    .A2(_11426_),
    .ZN(_11427_)
  );
  INV_X1 _45906_ (
    .A(_11427_),
    .ZN(_11428_)
  );
  AND2_X1 _45907_ (
    .A1(_11425_),
    .A2(_11428_),
    .ZN(_11429_)
  );
  INV_X1 _45908_ (
    .A(_11429_),
    .ZN(_00365_)
  );
  AND2_X1 _45909_ (
    .A1(instr_lh),
    .A2(_02901_),
    .ZN(_11430_)
  );
  INV_X1 _45910_ (
    .A(_11430_),
    .ZN(_11431_)
  );
  AND2_X1 _45911_ (
    .A1(_11379_),
    .A2(_11426_),
    .ZN(_11432_)
  );
  INV_X1 _45912_ (
    .A(_11432_),
    .ZN(_11433_)
  );
  AND2_X1 _45913_ (
    .A1(_11431_),
    .A2(_11433_),
    .ZN(_11434_)
  );
  INV_X1 _45914_ (
    .A(_11434_),
    .ZN(_00366_)
  );
  AND2_X1 _45915_ (
    .A1(instr_lw),
    .A2(_02901_),
    .ZN(_11435_)
  );
  INV_X1 _45916_ (
    .A(_11435_),
    .ZN(_11436_)
  );
  AND2_X1 _45917_ (
    .A1(_02905_),
    .A2(_11426_),
    .ZN(_11437_)
  );
  INV_X1 _45918_ (
    .A(_11437_),
    .ZN(_11438_)
  );
  AND2_X1 _45919_ (
    .A1(_11436_),
    .A2(_11438_),
    .ZN(_11439_)
  );
  INV_X1 _45920_ (
    .A(_11439_),
    .ZN(_00367_)
  );
  AND2_X1 _45921_ (
    .A1(instr_lbu),
    .A2(_02901_),
    .ZN(_11440_)
  );
  INV_X1 _45922_ (
    .A(_11440_),
    .ZN(_11441_)
  );
  AND2_X1 _45923_ (
    .A1(_11385_),
    .A2(_11426_),
    .ZN(_11442_)
  );
  INV_X1 _45924_ (
    .A(_11442_),
    .ZN(_11443_)
  );
  AND2_X1 _45925_ (
    .A1(_11441_),
    .A2(_11443_),
    .ZN(_11444_)
  );
  INV_X1 _45926_ (
    .A(_11444_),
    .ZN(_00368_)
  );
  AND2_X1 _45927_ (
    .A1(instr_lhu),
    .A2(_02901_),
    .ZN(_11445_)
  );
  INV_X1 _45928_ (
    .A(_11445_),
    .ZN(_11446_)
  );
  AND2_X1 _45929_ (
    .A1(_11392_),
    .A2(_11426_),
    .ZN(_11447_)
  );
  INV_X1 _45930_ (
    .A(_11447_),
    .ZN(_11448_)
  );
  AND2_X1 _45931_ (
    .A1(_11446_),
    .A2(_11448_),
    .ZN(_11449_)
  );
  INV_X1 _45932_ (
    .A(_11449_),
    .ZN(_00369_)
  );
  AND2_X1 _45933_ (
    .A1(resetn),
    .A2(_22025_),
    .ZN(_11450_)
  );
  AND2_X1 _45934_ (
    .A1(_22053_),
    .A2(_11450_),
    .ZN(_11451_)
  );
  AND2_X1 _45935_ (
    .A1(_22251_),
    .A2(_11451_),
    .ZN(_11452_)
  );
  AND2_X1 _45936_ (
    .A1(_22268_),
    .A2(_11452_),
    .ZN(_00370_)
  );
  AND2_X1 _45937_ (
    .A1(instr_sh),
    .A2(_02901_),
    .ZN(_11453_)
  );
  INV_X1 _45938_ (
    .A(_11453_),
    .ZN(_11454_)
  );
  AND2_X1 _45939_ (
    .A1(_02907_),
    .A2(_11379_),
    .ZN(_11455_)
  );
  INV_X1 _45940_ (
    .A(_11455_),
    .ZN(_11456_)
  );
  AND2_X1 _45941_ (
    .A1(_11454_),
    .A2(_11456_),
    .ZN(_11457_)
  );
  INV_X1 _45942_ (
    .A(_11457_),
    .ZN(_00371_)
  );
  AND2_X1 _45943_ (
    .A1(instr_addi),
    .A2(_11368_),
    .ZN(_11458_)
  );
  INV_X1 _45944_ (
    .A(_11458_),
    .ZN(_11459_)
  );
  AND2_X1 _45945_ (
    .A1(is_alu_reg_imm),
    .A2(_02900_),
    .ZN(_11460_)
  );
  AND2_X1 _45946_ (
    .A1(resetn),
    .A2(_11460_),
    .ZN(_11461_)
  );
  AND2_X1 _45947_ (
    .A1(_11372_),
    .A2(_11461_),
    .ZN(_11462_)
  );
  INV_X1 _45948_ (
    .A(_11462_),
    .ZN(_11463_)
  );
  AND2_X1 _45949_ (
    .A1(_11459_),
    .A2(_11463_),
    .ZN(_11464_)
  );
  INV_X1 _45950_ (
    .A(_11464_),
    .ZN(_00372_)
  );
  AND2_X1 _45951_ (
    .A1(instr_slti),
    .A2(_11368_),
    .ZN(_11465_)
  );
  INV_X1 _45952_ (
    .A(_11465_),
    .ZN(_11466_)
  );
  AND2_X1 _45953_ (
    .A1(_02905_),
    .A2(_11461_),
    .ZN(_11467_)
  );
  INV_X1 _45954_ (
    .A(_11467_),
    .ZN(_11468_)
  );
  AND2_X1 _45955_ (
    .A1(_11466_),
    .A2(_11468_),
    .ZN(_11469_)
  );
  INV_X1 _45956_ (
    .A(_11469_),
    .ZN(_00373_)
  );
  AND2_X1 _45957_ (
    .A1(_21234_),
    .A2(_11406_),
    .ZN(_11470_)
  );
  INV_X1 _45958_ (
    .A(_11470_),
    .ZN(_11471_)
  );
  AND2_X1 _45959_ (
    .A1(_11461_),
    .A2(_11470_),
    .ZN(_11472_)
  );
  INV_X1 _45960_ (
    .A(_11472_),
    .ZN(_11473_)
  );
  AND2_X1 _45961_ (
    .A1(instr_sltiu),
    .A2(_11368_),
    .ZN(_11474_)
  );
  INV_X1 _45962_ (
    .A(_11474_),
    .ZN(_11475_)
  );
  AND2_X1 _45963_ (
    .A1(_11473_),
    .A2(_11475_),
    .ZN(_11476_)
  );
  INV_X1 _45964_ (
    .A(_11476_),
    .ZN(_00374_)
  );
  AND2_X1 _45965_ (
    .A1(instr_xori),
    .A2(_11368_),
    .ZN(_11477_)
  );
  INV_X1 _45966_ (
    .A(_11477_),
    .ZN(_11478_)
  );
  AND2_X1 _45967_ (
    .A1(_11385_),
    .A2(_11461_),
    .ZN(_11479_)
  );
  INV_X1 _45968_ (
    .A(_11479_),
    .ZN(_11480_)
  );
  AND2_X1 _45969_ (
    .A1(_11478_),
    .A2(_11480_),
    .ZN(_11481_)
  );
  INV_X1 _45970_ (
    .A(_11481_),
    .ZN(_00375_)
  );
  AND2_X1 _45971_ (
    .A1(instr_ori),
    .A2(_11368_),
    .ZN(_11482_)
  );
  INV_X1 _45972_ (
    .A(_11482_),
    .ZN(_11483_)
  );
  AND2_X1 _45973_ (
    .A1(_11399_),
    .A2(_11461_),
    .ZN(_11484_)
  );
  INV_X1 _45974_ (
    .A(_11484_),
    .ZN(_11485_)
  );
  AND2_X1 _45975_ (
    .A1(_11483_),
    .A2(_11485_),
    .ZN(_11486_)
  );
  INV_X1 _45976_ (
    .A(_11486_),
    .ZN(_00376_)
  );
  AND2_X1 _45977_ (
    .A1(instr_andi),
    .A2(_11368_),
    .ZN(_11487_)
  );
  INV_X1 _45978_ (
    .A(_11487_),
    .ZN(_11488_)
  );
  AND2_X1 _45979_ (
    .A1(_11407_),
    .A2(_11461_),
    .ZN(_11489_)
  );
  INV_X1 _45980_ (
    .A(_11489_),
    .ZN(_11490_)
  );
  AND2_X1 _45981_ (
    .A1(_11488_),
    .A2(_11490_),
    .ZN(_11491_)
  );
  INV_X1 _45982_ (
    .A(_11491_),
    .ZN(_00377_)
  );
  AND2_X1 _45983_ (
    .A1(instr_sb),
    .A2(_02901_),
    .ZN(_11492_)
  );
  INV_X1 _45984_ (
    .A(_11492_),
    .ZN(_11493_)
  );
  AND2_X1 _45985_ (
    .A1(_02907_),
    .A2(_11372_),
    .ZN(_11494_)
  );
  INV_X1 _45986_ (
    .A(_11494_),
    .ZN(_11495_)
  );
  AND2_X1 _45987_ (
    .A1(_11493_),
    .A2(_11495_),
    .ZN(_11496_)
  );
  INV_X1 _45988_ (
    .A(_11496_),
    .ZN(_00378_)
  );
  AND2_X1 _45989_ (
    .A1(instr_slli),
    .A2(_02901_),
    .ZN(_11497_)
  );
  INV_X1 _45990_ (
    .A(_11497_),
    .ZN(_11498_)
  );
  AND2_X1 _45991_ (
    .A1(_21245_),
    .A2(_21246_),
    .ZN(_11499_)
  );
  AND2_X1 _45992_ (
    .A1(_21247_),
    .A2(_21248_),
    .ZN(_11500_)
  );
  AND2_X1 _45993_ (
    .A1(_21251_),
    .A2(_11500_),
    .ZN(_11501_)
  );
  AND2_X1 _45994_ (
    .A1(_11499_),
    .A2(_11501_),
    .ZN(_11502_)
  );
  AND2_X1 _45995_ (
    .A1(_21249_),
    .A2(_21250_),
    .ZN(_11503_)
  );
  AND2_X1 _45996_ (
    .A1(_11502_),
    .A2(_11503_),
    .ZN(_11504_)
  );
  INV_X1 _45997_ (
    .A(_11504_),
    .ZN(_11505_)
  );
  AND2_X1 _45998_ (
    .A1(_11379_),
    .A2(_11504_),
    .ZN(_11506_)
  );
  INV_X1 _45999_ (
    .A(_11506_),
    .ZN(_11507_)
  );
  AND2_X1 _46000_ (
    .A1(_11460_),
    .A2(_11506_),
    .ZN(_11508_)
  );
  INV_X1 _46001_ (
    .A(_11508_),
    .ZN(_11509_)
  );
  AND2_X1 _46002_ (
    .A1(_11498_),
    .A2(_11509_),
    .ZN(_11510_)
  );
  INV_X1 _46003_ (
    .A(_11510_),
    .ZN(_00379_)
  );
  AND2_X1 _46004_ (
    .A1(instr_srli),
    .A2(_02901_),
    .ZN(_11511_)
  );
  INV_X1 _46005_ (
    .A(_11511_),
    .ZN(_11512_)
  );
  AND2_X1 _46006_ (
    .A1(is_alu_reg_imm),
    .A2(_11392_),
    .ZN(_11513_)
  );
  AND2_X1 _46007_ (
    .A1(_02900_),
    .A2(_11504_),
    .ZN(_11514_)
  );
  AND2_X1 _46008_ (
    .A1(_11513_),
    .A2(_11514_),
    .ZN(_11515_)
  );
  INV_X1 _46009_ (
    .A(_11515_),
    .ZN(_11516_)
  );
  AND2_X1 _46010_ (
    .A1(_11512_),
    .A2(_11516_),
    .ZN(_11517_)
  );
  INV_X1 _46011_ (
    .A(_11517_),
    .ZN(_00380_)
  );
  AND2_X1 _46012_ (
    .A1(instr_add),
    .A2(_11368_),
    .ZN(_11518_)
  );
  INV_X1 _46013_ (
    .A(_11518_),
    .ZN(_11519_)
  );
  AND2_X1 _46014_ (
    .A1(resetn),
    .A2(is_alu_reg_reg),
    .ZN(_11520_)
  );
  AND2_X1 _46015_ (
    .A1(_11372_),
    .A2(_11520_),
    .ZN(_11521_)
  );
  AND2_X1 _46016_ (
    .A1(_11514_),
    .A2(_11521_),
    .ZN(_11522_)
  );
  INV_X1 _46017_ (
    .A(_11522_),
    .ZN(_11523_)
  );
  AND2_X1 _46018_ (
    .A1(_11519_),
    .A2(_11523_),
    .ZN(_11524_)
  );
  INV_X1 _46019_ (
    .A(_11524_),
    .ZN(_00381_)
  );
  AND2_X1 _46020_ (
    .A1(_21249_),
    .A2(_22040_),
    .ZN(_11525_)
  );
  AND2_X1 _46021_ (
    .A1(_11502_),
    .A2(_11525_),
    .ZN(_11526_)
  );
  INV_X1 _46022_ (
    .A(_11526_),
    .ZN(_11527_)
  );
  AND2_X1 _46023_ (
    .A1(_02900_),
    .A2(_11526_),
    .ZN(_11528_)
  );
  AND2_X1 _46024_ (
    .A1(_11521_),
    .A2(_11528_),
    .ZN(_11529_)
  );
  INV_X1 _46025_ (
    .A(_11529_),
    .ZN(_11530_)
  );
  AND2_X1 _46026_ (
    .A1(instr_sub),
    .A2(_11368_),
    .ZN(_11531_)
  );
  INV_X1 _46027_ (
    .A(_11531_),
    .ZN(_11532_)
  );
  AND2_X1 _46028_ (
    .A1(_11530_),
    .A2(_11532_),
    .ZN(_11533_)
  );
  INV_X1 _46029_ (
    .A(_11533_),
    .ZN(_00382_)
  );
  AND2_X1 _46030_ (
    .A1(instr_sll),
    .A2(_11368_),
    .ZN(_11534_)
  );
  INV_X1 _46031_ (
    .A(_11534_),
    .ZN(_11535_)
  );
  AND2_X1 _46032_ (
    .A1(is_alu_reg_reg),
    .A2(_02900_),
    .ZN(_11536_)
  );
  AND2_X1 _46033_ (
    .A1(_02900_),
    .A2(_11520_),
    .ZN(_11537_)
  );
  AND2_X1 _46034_ (
    .A1(_11506_),
    .A2(_11537_),
    .ZN(_11538_)
  );
  INV_X1 _46035_ (
    .A(_11538_),
    .ZN(_11539_)
  );
  AND2_X1 _46036_ (
    .A1(_11535_),
    .A2(_11539_),
    .ZN(_11540_)
  );
  INV_X1 _46037_ (
    .A(_11540_),
    .ZN(_00383_)
  );
  AND2_X1 _46038_ (
    .A1(instr_slt),
    .A2(_11368_),
    .ZN(_11541_)
  );
  INV_X1 _46039_ (
    .A(_11541_),
    .ZN(_11542_)
  );
  AND2_X1 _46040_ (
    .A1(_11514_),
    .A2(_11520_),
    .ZN(_11543_)
  );
  AND2_X1 _46041_ (
    .A1(_02905_),
    .A2(_11543_),
    .ZN(_11544_)
  );
  INV_X1 _46042_ (
    .A(_11544_),
    .ZN(_11545_)
  );
  AND2_X1 _46043_ (
    .A1(_11542_),
    .A2(_11545_),
    .ZN(_11546_)
  );
  INV_X1 _46044_ (
    .A(_11546_),
    .ZN(_00384_)
  );
  AND2_X1 _46045_ (
    .A1(instr_sltu),
    .A2(_11368_),
    .ZN(_11547_)
  );
  INV_X1 _46046_ (
    .A(_11547_),
    .ZN(_11548_)
  );
  AND2_X1 _46047_ (
    .A1(_11470_),
    .A2(_11543_),
    .ZN(_11549_)
  );
  INV_X1 _46048_ (
    .A(_11549_),
    .ZN(_11550_)
  );
  AND2_X1 _46049_ (
    .A1(_11548_),
    .A2(_11550_),
    .ZN(_11551_)
  );
  INV_X1 _46050_ (
    .A(_11551_),
    .ZN(_00385_)
  );
  AND2_X1 _46051_ (
    .A1(instr_xor),
    .A2(_11368_),
    .ZN(_11552_)
  );
  INV_X1 _46052_ (
    .A(_11552_),
    .ZN(_11553_)
  );
  AND2_X1 _46053_ (
    .A1(_11385_),
    .A2(_11543_),
    .ZN(_11554_)
  );
  INV_X1 _46054_ (
    .A(_11554_),
    .ZN(_11555_)
  );
  AND2_X1 _46055_ (
    .A1(_11553_),
    .A2(_11555_),
    .ZN(_11556_)
  );
  INV_X1 _46056_ (
    .A(_11556_),
    .ZN(_00386_)
  );
  AND2_X1 _46057_ (
    .A1(instr_srl),
    .A2(_11368_),
    .ZN(_11557_)
  );
  INV_X1 _46058_ (
    .A(_11557_),
    .ZN(_11558_)
  );
  AND2_X1 _46059_ (
    .A1(_11392_),
    .A2(_11520_),
    .ZN(_11559_)
  );
  AND2_X1 _46060_ (
    .A1(_11514_),
    .A2(_11559_),
    .ZN(_11560_)
  );
  INV_X1 _46061_ (
    .A(_11560_),
    .ZN(_11561_)
  );
  AND2_X1 _46062_ (
    .A1(_11558_),
    .A2(_11561_),
    .ZN(_11562_)
  );
  INV_X1 _46063_ (
    .A(_11562_),
    .ZN(_00387_)
  );
  AND2_X1 _46064_ (
    .A1(instr_sra),
    .A2(_11368_),
    .ZN(_11563_)
  );
  INV_X1 _46065_ (
    .A(_11563_),
    .ZN(_11564_)
  );
  AND2_X1 _46066_ (
    .A1(_11528_),
    .A2(_11559_),
    .ZN(_11565_)
  );
  INV_X1 _46067_ (
    .A(_11565_),
    .ZN(_11566_)
  );
  AND2_X1 _46068_ (
    .A1(_11564_),
    .A2(_11566_),
    .ZN(_11567_)
  );
  INV_X1 _46069_ (
    .A(_11567_),
    .ZN(_00388_)
  );
  AND2_X1 _46070_ (
    .A1(instr_or),
    .A2(_11368_),
    .ZN(_11568_)
  );
  INV_X1 _46071_ (
    .A(_11568_),
    .ZN(_11569_)
  );
  AND2_X1 _46072_ (
    .A1(_11399_),
    .A2(_11543_),
    .ZN(_11570_)
  );
  INV_X1 _46073_ (
    .A(_11570_),
    .ZN(_11571_)
  );
  AND2_X1 _46074_ (
    .A1(_11569_),
    .A2(_11571_),
    .ZN(_11572_)
  );
  INV_X1 _46075_ (
    .A(_11572_),
    .ZN(_00389_)
  );
  AND2_X1 _46076_ (
    .A1(instr_and),
    .A2(_11368_),
    .ZN(_11573_)
  );
  INV_X1 _46077_ (
    .A(_11573_),
    .ZN(_11574_)
  );
  AND2_X1 _46078_ (
    .A1(_11407_),
    .A2(_11543_),
    .ZN(_11575_)
  );
  INV_X1 _46079_ (
    .A(_11575_),
    .ZN(_11576_)
  );
  AND2_X1 _46080_ (
    .A1(_11574_),
    .A2(_11576_),
    .ZN(_11577_)
  );
  INV_X1 _46081_ (
    .A(_11577_),
    .ZN(_00390_)
  );
  AND2_X1 _46082_ (
    .A1(instr_srai),
    .A2(_02901_),
    .ZN(_11578_)
  );
  INV_X1 _46083_ (
    .A(_11578_),
    .ZN(_11579_)
  );
  AND2_X1 _46084_ (
    .A1(_11513_),
    .A2(_11528_),
    .ZN(_11580_)
  );
  INV_X1 _46085_ (
    .A(_11580_),
    .ZN(_11581_)
  );
  AND2_X1 _46086_ (
    .A1(_11579_),
    .A2(_11581_),
    .ZN(_11582_)
  );
  INV_X1 _46087_ (
    .A(_11582_),
    .ZN(_00391_)
  );
  AND2_X1 _46088_ (
    .A1(instr_rdcycle),
    .A2(_02901_),
    .ZN(_11583_)
  );
  INV_X1 _46089_ (
    .A(_11583_),
    .ZN(_11584_)
  );
  AND2_X1 _46090_ (
    .A1(_21244_),
    .A2(_02900_),
    .ZN(_11585_)
  );
  AND2_X1 _46091_ (
    .A1(_11499_),
    .A2(_11585_),
    .ZN(_11586_)
  );
  AND2_X1 _46092_ (
    .A1(_21247_),
    .A2(_11586_),
    .ZN(_11587_)
  );
  AND2_X1 _46093_ (
    .A1(_21235_),
    .A2(_21236_),
    .ZN(_11588_)
  );
  AND2_X1 _46094_ (
    .A1(_21237_),
    .A2(_21238_),
    .ZN(_11589_)
  );
  AND2_X1 _46095_ (
    .A1(_11588_),
    .A2(_11589_),
    .ZN(_11590_)
  );
  AND2_X1 _46096_ (
    .A1(_22045_),
    .A2(_22046_),
    .ZN(_11591_)
  );
  AND2_X1 _46097_ (
    .A1(_11525_),
    .A2(_11591_),
    .ZN(_11592_)
  );
  AND2_X1 _46098_ (
    .A1(_11590_),
    .A2(_11592_),
    .ZN(_11593_)
  );
  AND2_X1 _46099_ (
    .A1(_22041_),
    .A2(_22042_),
    .ZN(_11594_)
  );
  AND2_X1 _46100_ (
    .A1(_22043_),
    .A2(_22044_),
    .ZN(_11595_)
  );
  AND2_X1 _46101_ (
    .A1(_11594_),
    .A2(_11595_),
    .ZN(_11596_)
  );
  AND2_X1 _46102_ (
    .A1(_21239_),
    .A2(_21248_),
    .ZN(_11597_)
  );
  AND2_X1 _46103_ (
    .A1(_21354_),
    .A2(_21356_),
    .ZN(_11598_)
  );
  AND2_X1 _46104_ (
    .A1(_11597_),
    .A2(_11598_),
    .ZN(_11599_)
  );
  AND2_X1 _46105_ (
    .A1(_11596_),
    .A2(_11599_),
    .ZN(_11600_)
  );
  AND2_X1 _46106_ (
    .A1(_02905_),
    .A2(_11600_),
    .ZN(_11601_)
  );
  AND2_X1 _46107_ (
    .A1(_11593_),
    .A2(_11601_),
    .ZN(_11602_)
  );
  AND2_X1 _46108_ (
    .A1(mem_rdata_q[20]),
    .A2(_00040_),
    .ZN(_11603_)
  );
  INV_X1 _46109_ (
    .A(_11603_),
    .ZN(_11604_)
  );
  AND2_X1 _46110_ (
    .A1(_21242_),
    .A2(_21243_),
    .ZN(_11605_)
  );
  AND2_X1 _46111_ (
    .A1(_21241_),
    .A2(_11604_),
    .ZN(_11606_)
  );
  AND2_X1 _46112_ (
    .A1(_11605_),
    .A2(_11606_),
    .ZN(_11607_)
  );
  AND2_X1 _46113_ (
    .A1(_11602_),
    .A2(_11607_),
    .ZN(_11608_)
  );
  AND2_X1 _46114_ (
    .A1(_11587_),
    .A2(_11608_),
    .ZN(_11609_)
  );
  INV_X1 _46115_ (
    .A(_11609_),
    .ZN(_11610_)
  );
  AND2_X1 _46116_ (
    .A1(_11584_),
    .A2(_11610_),
    .ZN(_11611_)
  );
  INV_X1 _46117_ (
    .A(_11611_),
    .ZN(_00392_)
  );
  AND2_X1 _46118_ (
    .A1(instr_rdcycleh),
    .A2(_02901_),
    .ZN(_11612_)
  );
  INV_X1 _46119_ (
    .A(_11612_),
    .ZN(_11613_)
  );
  AND2_X1 _46120_ (
    .A1(_22039_),
    .A2(_11586_),
    .ZN(_11614_)
  );
  AND2_X1 _46121_ (
    .A1(_11608_),
    .A2(_11614_),
    .ZN(_11615_)
  );
  INV_X1 _46122_ (
    .A(_11615_),
    .ZN(_11616_)
  );
  AND2_X1 _46123_ (
    .A1(_11613_),
    .A2(_11616_),
    .ZN(_11617_)
  );
  INV_X1 _46124_ (
    .A(_11617_),
    .ZN(_00393_)
  );
  AND2_X1 _46125_ (
    .A1(instr_rdinstr),
    .A2(_02901_),
    .ZN(_11618_)
  );
  INV_X1 _46126_ (
    .A(_11618_),
    .ZN(_11619_)
  );
  AND2_X1 _46127_ (
    .A1(_21240_),
    .A2(_22038_),
    .ZN(_11620_)
  );
  AND2_X1 _46128_ (
    .A1(_11605_),
    .A2(_11620_),
    .ZN(_11621_)
  );
  AND2_X1 _46129_ (
    .A1(_11602_),
    .A2(_11621_),
    .ZN(_11622_)
  );
  AND2_X1 _46130_ (
    .A1(_11587_),
    .A2(_11622_),
    .ZN(_11623_)
  );
  INV_X1 _46131_ (
    .A(_11623_),
    .ZN(_11624_)
  );
  AND2_X1 _46132_ (
    .A1(_11619_),
    .A2(_11624_),
    .ZN(_11625_)
  );
  INV_X1 _46133_ (
    .A(_11625_),
    .ZN(_00394_)
  );
  AND2_X1 _46134_ (
    .A1(instr_rdinstrh),
    .A2(_02901_),
    .ZN(_11626_)
  );
  INV_X1 _46135_ (
    .A(_11626_),
    .ZN(_11627_)
  );
  AND2_X1 _46136_ (
    .A1(_11614_),
    .A2(_11622_),
    .ZN(_11628_)
  );
  INV_X1 _46137_ (
    .A(_11628_),
    .ZN(_11629_)
  );
  AND2_X1 _46138_ (
    .A1(_11627_),
    .A2(_11629_),
    .ZN(_11630_)
  );
  INV_X1 _46139_ (
    .A(_11630_),
    .ZN(_00395_)
  );
  AND2_X1 _46140_ (
    .A1(instr_fence),
    .A2(_11368_),
    .ZN(_11631_)
  );
  INV_X1 _46141_ (
    .A(_11631_),
    .ZN(_11632_)
  );
  AND2_X1 _46142_ (
    .A1(resetn),
    .A2(_21357_),
    .ZN(_11633_)
  );
  AND2_X1 _46143_ (
    .A1(_02900_),
    .A2(_11633_),
    .ZN(_11634_)
  );
  AND2_X1 _46144_ (
    .A1(_11591_),
    .A2(_11634_),
    .ZN(_11635_)
  );
  AND2_X1 _46145_ (
    .A1(_21358_),
    .A2(_21359_),
    .ZN(_11636_)
  );
  AND2_X1 _46146_ (
    .A1(_22047_),
    .A2(_22048_),
    .ZN(_11637_)
  );
  AND2_X1 _46147_ (
    .A1(_11636_),
    .A2(_11637_),
    .ZN(_11638_)
  );
  AND2_X1 _46148_ (
    .A1(_11372_),
    .A2(_11638_),
    .ZN(_11639_)
  );
  AND2_X1 _46149_ (
    .A1(_11635_),
    .A2(_11639_),
    .ZN(_11640_)
  );
  INV_X1 _46150_ (
    .A(_11640_),
    .ZN(_11641_)
  );
  AND2_X1 _46151_ (
    .A1(_11632_),
    .A2(_11641_),
    .ZN(_11642_)
  );
  INV_X1 _46152_ (
    .A(_11642_),
    .ZN(_00396_)
  );
  AND2_X1 _46153_ (
    .A1(_21277_),
    .A2(_11307_),
    .ZN(_11643_)
  );
  INV_X1 _46154_ (
    .A(_11643_),
    .ZN(_11644_)
  );
  AND2_X1 _46155_ (
    .A1(_10396_),
    .A2(_11306_),
    .ZN(_11645_)
  );
  INV_X1 _46156_ (
    .A(_11645_),
    .ZN(_11646_)
  );
  AND2_X1 _46157_ (
    .A1(_11644_),
    .A2(_11646_),
    .ZN(_00397_)
  );
  AND2_X1 _46158_ (
    .A1(_21278_),
    .A2(_11307_),
    .ZN(_11647_)
  );
  INV_X1 _46159_ (
    .A(_11647_),
    .ZN(_11648_)
  );
  AND2_X1 _46160_ (
    .A1(_10401_),
    .A2(_11306_),
    .ZN(_11649_)
  );
  INV_X1 _46161_ (
    .A(_11649_),
    .ZN(_11650_)
  );
  AND2_X1 _46162_ (
    .A1(_11648_),
    .A2(_11650_),
    .ZN(_00398_)
  );
  AND2_X1 _46163_ (
    .A1(_21279_),
    .A2(_11307_),
    .ZN(_11651_)
  );
  INV_X1 _46164_ (
    .A(_11651_),
    .ZN(_11652_)
  );
  AND2_X1 _46165_ (
    .A1(_10406_),
    .A2(_11306_),
    .ZN(_11653_)
  );
  INV_X1 _46166_ (
    .A(_11653_),
    .ZN(_11654_)
  );
  AND2_X1 _46167_ (
    .A1(_11652_),
    .A2(_11654_),
    .ZN(_00399_)
  );
  AND2_X1 _46168_ (
    .A1(_21280_),
    .A2(_11307_),
    .ZN(_11655_)
  );
  INV_X1 _46169_ (
    .A(_11655_),
    .ZN(_11656_)
  );
  AND2_X1 _46170_ (
    .A1(_10411_),
    .A2(_11306_),
    .ZN(_11657_)
  );
  INV_X1 _46171_ (
    .A(_11657_),
    .ZN(_11658_)
  );
  AND2_X1 _46172_ (
    .A1(_11656_),
    .A2(_11658_),
    .ZN(_00400_)
  );
  AND2_X1 _46173_ (
    .A1(_21281_),
    .A2(_11307_),
    .ZN(_11659_)
  );
  INV_X1 _46174_ (
    .A(_11659_),
    .ZN(_11660_)
  );
  AND2_X1 _46175_ (
    .A1(_10416_),
    .A2(_11306_),
    .ZN(_11661_)
  );
  INV_X1 _46176_ (
    .A(_11661_),
    .ZN(_11662_)
  );
  AND2_X1 _46177_ (
    .A1(_11660_),
    .A2(_11662_),
    .ZN(_00401_)
  );
  AND2_X1 _46178_ (
    .A1(_21282_),
    .A2(_11307_),
    .ZN(_11663_)
  );
  INV_X1 _46179_ (
    .A(_11663_),
    .ZN(_11664_)
  );
  AND2_X1 _46180_ (
    .A1(_10461_),
    .A2(_11306_),
    .ZN(_11665_)
  );
  INV_X1 _46181_ (
    .A(_11665_),
    .ZN(_11666_)
  );
  AND2_X1 _46182_ (
    .A1(_11664_),
    .A2(_11666_),
    .ZN(_00402_)
  );
  AND2_X1 _46183_ (
    .A1(_21283_),
    .A2(_11307_),
    .ZN(_11667_)
  );
  INV_X1 _46184_ (
    .A(_11667_),
    .ZN(_11668_)
  );
  AND2_X1 _46185_ (
    .A1(_10466_),
    .A2(_11306_),
    .ZN(_11669_)
  );
  INV_X1 _46186_ (
    .A(_11669_),
    .ZN(_11670_)
  );
  AND2_X1 _46187_ (
    .A1(_11668_),
    .A2(_11670_),
    .ZN(_00403_)
  );
  AND2_X1 _46188_ (
    .A1(_21284_),
    .A2(_11307_),
    .ZN(_11671_)
  );
  INV_X1 _46189_ (
    .A(_11671_),
    .ZN(_11672_)
  );
  AND2_X1 _46190_ (
    .A1(_10471_),
    .A2(_11306_),
    .ZN(_11673_)
  );
  INV_X1 _46191_ (
    .A(_11673_),
    .ZN(_11674_)
  );
  AND2_X1 _46192_ (
    .A1(_11672_),
    .A2(_11674_),
    .ZN(_00404_)
  );
  AND2_X1 _46193_ (
    .A1(_21285_),
    .A2(_11307_),
    .ZN(_11675_)
  );
  INV_X1 _46194_ (
    .A(_11675_),
    .ZN(_11676_)
  );
  AND2_X1 _46195_ (
    .A1(_10476_),
    .A2(_11306_),
    .ZN(_11677_)
  );
  INV_X1 _46196_ (
    .A(_11677_),
    .ZN(_11678_)
  );
  AND2_X1 _46197_ (
    .A1(_11676_),
    .A2(_11678_),
    .ZN(_00405_)
  );
  AND2_X1 _46198_ (
    .A1(mem_rdata_q[7]),
    .A2(_02907_),
    .ZN(_11679_)
  );
  INV_X1 _46199_ (
    .A(_11679_),
    .ZN(_11680_)
  );
  AND2_X1 _46200_ (
    .A1(_21262_),
    .A2(_21292_),
    .ZN(_11681_)
  );
  INV_X1 _46201_ (
    .A(_11681_),
    .ZN(_11682_)
  );
  AND2_X1 _46202_ (
    .A1(_21288_),
    .A2(_11681_),
    .ZN(_11683_)
  );
  INV_X1 _46203_ (
    .A(_11683_),
    .ZN(_11684_)
  );
  AND2_X1 _46204_ (
    .A1(mem_rdata_q[20]),
    .A2(_02900_),
    .ZN(_11685_)
  );
  AND2_X1 _46205_ (
    .A1(_11684_),
    .A2(_11685_),
    .ZN(_11686_)
  );
  INV_X1 _46206_ (
    .A(_11686_),
    .ZN(_11687_)
  );
  AND2_X1 _46207_ (
    .A1(decoded_imm[0]),
    .A2(_02901_),
    .ZN(_11688_)
  );
  INV_X1 _46208_ (
    .A(_11688_),
    .ZN(_11689_)
  );
  AND2_X1 _46209_ (
    .A1(_11680_),
    .A2(_11689_),
    .ZN(_11690_)
  );
  AND2_X1 _46210_ (
    .A1(_11687_),
    .A2(_11690_),
    .ZN(_11691_)
  );
  INV_X1 _46211_ (
    .A(_11691_),
    .ZN(_00406_)
  );
  AND2_X1 _46212_ (
    .A1(_21287_),
    .A2(_11307_),
    .ZN(_11692_)
  );
  INV_X1 _46213_ (
    .A(_11692_),
    .ZN(_11693_)
  );
  AND2_X1 _46214_ (
    .A1(_10511_),
    .A2(_11306_),
    .ZN(_11694_)
  );
  INV_X1 _46215_ (
    .A(_11694_),
    .ZN(_11695_)
  );
  AND2_X1 _46216_ (
    .A1(_11693_),
    .A2(_11695_),
    .ZN(_00407_)
  );
  AND2_X1 _46217_ (
    .A1(is_lb_lh_lw_lbu_lhu),
    .A2(_11307_),
    .ZN(_11696_)
  );
  INV_X1 _46218_ (
    .A(_11696_),
    .ZN(_11697_)
  );
  AND2_X1 _46219_ (
    .A1(_11333_),
    .A2(_11338_),
    .ZN(_11698_)
  );
  AND2_X1 _46220_ (
    .A1(_11344_),
    .A2(_11698_),
    .ZN(_11699_)
  );
  AND2_X1 _46221_ (
    .A1(_11316_),
    .A2(_11327_),
    .ZN(_11700_)
  );
  AND2_X1 _46222_ (
    .A1(_11321_),
    .A2(_11700_),
    .ZN(_11701_)
  );
  AND2_X1 _46223_ (
    .A1(_11306_),
    .A2(_11701_),
    .ZN(_11702_)
  );
  AND2_X1 _46224_ (
    .A1(_11699_),
    .A2(_11702_),
    .ZN(_11703_)
  );
  INV_X1 _46225_ (
    .A(_11703_),
    .ZN(_11704_)
  );
  AND2_X1 _46226_ (
    .A1(_11697_),
    .A2(_11704_),
    .ZN(_11705_)
  );
  INV_X1 _46227_ (
    .A(_11705_),
    .ZN(_00408_)
  );
  AND2_X1 _46228_ (
    .A1(is_slli_srli_srai),
    .A2(_02901_),
    .ZN(_11706_)
  );
  INV_X1 _46229_ (
    .A(_11706_),
    .ZN(_11707_)
  );
  AND2_X1 _46230_ (
    .A1(_11505_),
    .A2(_11527_),
    .ZN(_11708_)
  );
  INV_X1 _46231_ (
    .A(_11708_),
    .ZN(_11709_)
  );
  AND2_X1 _46232_ (
    .A1(_11393_),
    .A2(_11507_),
    .ZN(_11710_)
  );
  INV_X1 _46233_ (
    .A(_11710_),
    .ZN(_11711_)
  );
  AND2_X1 _46234_ (
    .A1(_11709_),
    .A2(_11711_),
    .ZN(_11712_)
  );
  AND2_X1 _46235_ (
    .A1(_11460_),
    .A2(_11712_),
    .ZN(_11713_)
  );
  INV_X1 _46236_ (
    .A(_11713_),
    .ZN(_11714_)
  );
  AND2_X1 _46237_ (
    .A1(_11707_),
    .A2(_11714_),
    .ZN(_11715_)
  );
  INV_X1 _46238_ (
    .A(_11715_),
    .ZN(_00409_)
  );
  AND2_X1 _46239_ (
    .A1(is_sb_sh_sw),
    .A2(_11307_),
    .ZN(_11716_)
  );
  INV_X1 _46240_ (
    .A(_11716_),
    .ZN(_11717_)
  );
  AND2_X1 _46241_ (
    .A1(_11333_),
    .A2(_11359_),
    .ZN(_11718_)
  );
  AND2_X1 _46242_ (
    .A1(_11702_),
    .A2(_11718_),
    .ZN(_11719_)
  );
  INV_X1 _46243_ (
    .A(_11719_),
    .ZN(_11720_)
  );
  AND2_X1 _46244_ (
    .A1(_11717_),
    .A2(_11720_),
    .ZN(_11721_)
  );
  INV_X1 _46245_ (
    .A(_11721_),
    .ZN(_00410_)
  );
  AND2_X1 _46246_ (
    .A1(is_sll_srl_sra),
    .A2(_02901_),
    .ZN(_11722_)
  );
  INV_X1 _46247_ (
    .A(_11722_),
    .ZN(_11723_)
  );
  AND2_X1 _46248_ (
    .A1(_11536_),
    .A2(_11712_),
    .ZN(_11724_)
  );
  INV_X1 _46249_ (
    .A(_11724_),
    .ZN(_11725_)
  );
  AND2_X1 _46250_ (
    .A1(_11723_),
    .A2(_11725_),
    .ZN(_11726_)
  );
  INV_X1 _46251_ (
    .A(_11726_),
    .ZN(_00411_)
  );
  AND2_X1 _46252_ (
    .A1(_11097_),
    .A2(_11307_),
    .ZN(_11727_)
  );
  INV_X1 _46253_ (
    .A(_11727_),
    .ZN(_11728_)
  );
  AND2_X1 _46254_ (
    .A1(_11360_),
    .A2(_11702_),
    .ZN(_11729_)
  );
  INV_X1 _46255_ (
    .A(_11729_),
    .ZN(_11730_)
  );
  AND2_X1 _46256_ (
    .A1(_11728_),
    .A2(_11730_),
    .ZN(_11731_)
  );
  INV_X1 _46257_ (
    .A(_11731_),
    .ZN(_00412_)
  );
  AND2_X1 _46258_ (
    .A1(_21056_),
    .A2(_22526_),
    .ZN(_11732_)
  );
  AND2_X1 _46259_ (
    .A1(_22525_),
    .A2(_11732_),
    .ZN(_11733_)
  );
  INV_X1 _46260_ (
    .A(_11733_),
    .ZN(_11734_)
  );
  AND2_X1 _46261_ (
    .A1(_02901_),
    .A2(_11734_),
    .ZN(_00413_)
  );
  AND2_X1 _46262_ (
    .A1(_11352_),
    .A2(_11702_),
    .ZN(_11735_)
  );
  INV_X1 _46263_ (
    .A(_11735_),
    .ZN(_11736_)
  );
  AND2_X1 _46264_ (
    .A1(is_alu_reg_imm),
    .A2(_11307_),
    .ZN(_11737_)
  );
  INV_X1 _46265_ (
    .A(_11737_),
    .ZN(_11738_)
  );
  AND2_X1 _46266_ (
    .A1(_11736_),
    .A2(_11738_),
    .ZN(_11739_)
  );
  INV_X1 _46267_ (
    .A(_11739_),
    .ZN(_00414_)
  );
  AND2_X1 _46268_ (
    .A1(_11400_),
    .A2(_11408_),
    .ZN(_11740_)
  );
  AND2_X1 _46269_ (
    .A1(_11471_),
    .A2(_11740_),
    .ZN(_11741_)
  );
  AND2_X1 _46270_ (
    .A1(_21262_),
    .A2(_02906_),
    .ZN(_11742_)
  );
  AND2_X1 _46271_ (
    .A1(_11373_),
    .A2(_11386_),
    .ZN(_11743_)
  );
  AND2_X1 _46272_ (
    .A1(_11742_),
    .A2(_11743_),
    .ZN(_11744_)
  );
  AND2_X1 _46273_ (
    .A1(_11741_),
    .A2(_11744_),
    .ZN(_11745_)
  );
  INV_X1 _46274_ (
    .A(_11745_),
    .ZN(_11746_)
  );
  AND2_X1 _46275_ (
    .A1(is_jalr_addi_slti_sltiu_xori_ori_andi),
    .A2(_02901_),
    .ZN(_11747_)
  );
  INV_X1 _46276_ (
    .A(_11747_),
    .ZN(_11748_)
  );
  AND2_X1 _46277_ (
    .A1(_02900_),
    .A2(_11682_),
    .ZN(_11749_)
  );
  AND2_X1 _46278_ (
    .A1(_11746_),
    .A2(_11749_),
    .ZN(_11750_)
  );
  INV_X1 _46279_ (
    .A(_11750_),
    .ZN(_11751_)
  );
  AND2_X1 _46280_ (
    .A1(_11748_),
    .A2(_11751_),
    .ZN(_11752_)
  );
  INV_X1 _46281_ (
    .A(_11752_),
    .ZN(_00415_)
  );
  AND2_X1 _46282_ (
    .A1(_21039_),
    .A2(_22506_),
    .ZN(_11753_)
  );
  INV_X1 _46283_ (
    .A(_11753_),
    .ZN(_11754_)
  );
  AND2_X1 _46284_ (
    .A1(_11368_),
    .A2(_11754_),
    .ZN(_00416_)
  );
  AND2_X1 _46285_ (
    .A1(is_alu_reg_reg),
    .A2(_11307_),
    .ZN(_11755_)
  );
  INV_X1 _46286_ (
    .A(_11755_),
    .ZN(_11756_)
  );
  AND2_X1 _46287_ (
    .A1(_11345_),
    .A2(_11702_),
    .ZN(_11757_)
  );
  INV_X1 _46288_ (
    .A(_11757_),
    .ZN(_11758_)
  );
  AND2_X1 _46289_ (
    .A1(_11756_),
    .A2(_11758_),
    .ZN(_11759_)
  );
  INV_X1 _46290_ (
    .A(_11759_),
    .ZN(_00417_)
  );
  AND2_X1 _46291_ (
    .A1(_21070_),
    .A2(_21071_),
    .ZN(_11760_)
  );
  INV_X1 _46292_ (
    .A(_11760_),
    .ZN(_11761_)
  );
  AND2_X1 _46293_ (
    .A1(_21069_),
    .A2(_11760_),
    .ZN(_11762_)
  );
  INV_X1 _46294_ (
    .A(_11762_),
    .ZN(_11763_)
  );
  AND2_X1 _46295_ (
    .A1(_22299_),
    .A2(_11760_),
    .ZN(_11764_)
  );
  INV_X1 _46296_ (
    .A(_11764_),
    .ZN(_11765_)
  );
  AND2_X1 _46297_ (
    .A1(resetn),
    .A2(_22305_),
    .ZN(_11766_)
  );
  AND2_X1 _46298_ (
    .A1(resetn),
    .A2(_22076_),
    .ZN(_11767_)
  );
  AND2_X1 _46299_ (
    .A1(_22305_),
    .A2(_11767_),
    .ZN(_11768_)
  );
  AND2_X1 _46300_ (
    .A1(_22305_),
    .A2(_11763_),
    .ZN(_11769_)
  );
  AND2_X1 _46301_ (
    .A1(_11765_),
    .A2(_11768_),
    .ZN(_11770_)
  );
  INV_X1 _46302_ (
    .A(_11770_),
    .ZN(_11771_)
  );
  AND2_X1 _46303_ (
    .A1(mem_instr),
    .A2(_11771_),
    .ZN(_11772_)
  );
  INV_X1 _46304_ (
    .A(_11772_),
    .ZN(_11773_)
  );
  AND2_X1 _46305_ (
    .A1(_21038_),
    .A2(_11767_),
    .ZN(_11774_)
  );
  AND2_X1 _46306_ (
    .A1(_11761_),
    .A2(_11768_),
    .ZN(_11775_)
  );
  AND2_X1 _46307_ (
    .A1(_21038_),
    .A2(_11775_),
    .ZN(_11776_)
  );
  INV_X1 _46308_ (
    .A(_11776_),
    .ZN(_11777_)
  );
  AND2_X1 _46309_ (
    .A1(_11773_),
    .A2(_11777_),
    .ZN(_11778_)
  );
  INV_X1 _46310_ (
    .A(_11778_),
    .ZN(_00418_)
  );
  AND2_X1 _46311_ (
    .A1(_11764_),
    .A2(_11768_),
    .ZN(_11779_)
  );
  INV_X1 _46312_ (
    .A(_11779_),
    .ZN(_11780_)
  );
  AND2_X1 _46313_ (
    .A1(resetn),
    .A2(trap),
    .ZN(_11781_)
  );
  AND2_X1 _46314_ (
    .A1(_22075_),
    .A2(_11781_),
    .ZN(_11782_)
  );
  INV_X1 _46315_ (
    .A(_11782_),
    .ZN(_11783_)
  );
  AND2_X1 _46316_ (
    .A1(_21348_),
    .A2(_22062_),
    .ZN(_11784_)
  );
  INV_X1 _46317_ (
    .A(_11784_),
    .ZN(_11785_)
  );
  AND2_X1 _46318_ (
    .A1(_21349_),
    .A2(_22061_),
    .ZN(_11786_)
  );
  INV_X1 _46319_ (
    .A(_11786_),
    .ZN(_11787_)
  );
  AND2_X1 _46320_ (
    .A1(_11785_),
    .A2(_11787_),
    .ZN(_11788_)
  );
  INV_X1 _46321_ (
    .A(_11788_),
    .ZN(_11789_)
  );
  AND2_X1 _46322_ (
    .A1(_22306_),
    .A2(_11767_),
    .ZN(_11790_)
  );
  AND2_X1 _46323_ (
    .A1(_11788_),
    .A2(_11790_),
    .ZN(_11791_)
  );
  INV_X1 _46324_ (
    .A(_11791_),
    .ZN(_11792_)
  );
  AND2_X1 _46325_ (
    .A1(_11780_),
    .A2(_11783_),
    .ZN(_11793_)
  );
  AND2_X1 _46326_ (
    .A1(_11792_),
    .A2(_11793_),
    .ZN(_11794_)
  );
  AND2_X1 _46327_ (
    .A1(_22308_),
    .A2(_11789_),
    .ZN(_11795_)
  );
  INV_X1 _46328_ (
    .A(_11795_),
    .ZN(_11796_)
  );
  AND2_X1 _46329_ (
    .A1(_11767_),
    .A2(_11795_),
    .ZN(_11797_)
  );
  INV_X1 _46330_ (
    .A(_11797_),
    .ZN(_11798_)
  );
  AND2_X1 _46331_ (
    .A1(_11794_),
    .A2(_11798_),
    .ZN(_11799_)
  );
  INV_X1 _46332_ (
    .A(_11799_),
    .ZN(_11800_)
  );
  AND2_X1 _46333_ (
    .A1(mem_valid),
    .A2(_11800_),
    .ZN(_11801_)
  );
  INV_X1 _46334_ (
    .A(_11801_),
    .ZN(_11802_)
  );
  AND2_X1 _46335_ (
    .A1(_11771_),
    .A2(_11802_),
    .ZN(_11803_)
  );
  INV_X1 _46336_ (
    .A(_11803_),
    .ZN(_00419_)
  );
  AND2_X1 _46337_ (
    .A1(reg_out[2]),
    .A2(_02913_),
    .ZN(_11804_)
  );
  INV_X1 _46338_ (
    .A(_11804_),
    .ZN(_11805_)
  );
  AND2_X1 _46339_ (
    .A1(_02933_),
    .A2(_11805_),
    .ZN(_11806_)
  );
  INV_X1 _46340_ (
    .A(_11806_),
    .ZN(_11807_)
  );
  AND2_X1 _46341_ (
    .A1(_11761_),
    .A2(_11807_),
    .ZN(_11808_)
  );
  INV_X1 _46342_ (
    .A(_11808_),
    .ZN(_11809_)
  );
  AND2_X1 _46343_ (
    .A1(reg_op1[2]),
    .A2(_11760_),
    .ZN(_11810_)
  );
  INV_X1 _46344_ (
    .A(_11810_),
    .ZN(_11811_)
  );
  AND2_X1 _46345_ (
    .A1(_11809_),
    .A2(_11811_),
    .ZN(_11812_)
  );
  INV_X1 _46346_ (
    .A(_11812_),
    .ZN(mem_la_addr[2])
  );
  AND2_X1 _46347_ (
    .A1(_21294_),
    .A2(_11771_),
    .ZN(_11813_)
  );
  INV_X1 _46348_ (
    .A(_11813_),
    .ZN(_11814_)
  );
  AND2_X1 _46349_ (
    .A1(_11770_),
    .A2(_11812_),
    .ZN(_11815_)
  );
  INV_X1 _46350_ (
    .A(_11815_),
    .ZN(_11816_)
  );
  AND2_X1 _46351_ (
    .A1(_11814_),
    .A2(_11816_),
    .ZN(_00420_)
  );
  AND2_X1 _46352_ (
    .A1(reg_out[3]),
    .A2(_02913_),
    .ZN(_11817_)
  );
  INV_X1 _46353_ (
    .A(_11817_),
    .ZN(_11818_)
  );
  AND2_X1 _46354_ (
    .A1(_02949_),
    .A2(_11818_),
    .ZN(_11819_)
  );
  INV_X1 _46355_ (
    .A(_11819_),
    .ZN(_11820_)
  );
  AND2_X1 _46356_ (
    .A1(_11761_),
    .A2(_11820_),
    .ZN(_11821_)
  );
  INV_X1 _46357_ (
    .A(_11821_),
    .ZN(_11822_)
  );
  AND2_X1 _46358_ (
    .A1(reg_op1[3]),
    .A2(_11760_),
    .ZN(_11823_)
  );
  INV_X1 _46359_ (
    .A(_11823_),
    .ZN(_11824_)
  );
  AND2_X1 _46360_ (
    .A1(_11822_),
    .A2(_11824_),
    .ZN(_11825_)
  );
  INV_X1 _46361_ (
    .A(_11825_),
    .ZN(mem_la_addr[3])
  );
  AND2_X1 _46362_ (
    .A1(_21295_),
    .A2(_11771_),
    .ZN(_11826_)
  );
  INV_X1 _46363_ (
    .A(_11826_),
    .ZN(_11827_)
  );
  AND2_X1 _46364_ (
    .A1(_11770_),
    .A2(_11825_),
    .ZN(_11828_)
  );
  INV_X1 _46365_ (
    .A(_11828_),
    .ZN(_11829_)
  );
  AND2_X1 _46366_ (
    .A1(_11827_),
    .A2(_11829_),
    .ZN(_00421_)
  );
  AND2_X1 _46367_ (
    .A1(reg_out[4]),
    .A2(_02913_),
    .ZN(_11830_)
  );
  INV_X1 _46368_ (
    .A(_11830_),
    .ZN(_11831_)
  );
  AND2_X1 _46369_ (
    .A1(_02965_),
    .A2(_11831_),
    .ZN(_11832_)
  );
  INV_X1 _46370_ (
    .A(_11832_),
    .ZN(_11833_)
  );
  AND2_X1 _46371_ (
    .A1(_11761_),
    .A2(_11833_),
    .ZN(_11834_)
  );
  INV_X1 _46372_ (
    .A(_11834_),
    .ZN(_11835_)
  );
  AND2_X1 _46373_ (
    .A1(reg_op1[4]),
    .A2(_11760_),
    .ZN(_11836_)
  );
  INV_X1 _46374_ (
    .A(_11836_),
    .ZN(_11837_)
  );
  AND2_X1 _46375_ (
    .A1(_11835_),
    .A2(_11837_),
    .ZN(_11838_)
  );
  INV_X1 _46376_ (
    .A(_11838_),
    .ZN(mem_la_addr[4])
  );
  AND2_X1 _46377_ (
    .A1(_21296_),
    .A2(_11771_),
    .ZN(_11839_)
  );
  INV_X1 _46378_ (
    .A(_11839_),
    .ZN(_11840_)
  );
  AND2_X1 _46379_ (
    .A1(_11770_),
    .A2(_11838_),
    .ZN(_11841_)
  );
  INV_X1 _46380_ (
    .A(_11841_),
    .ZN(_11842_)
  );
  AND2_X1 _46381_ (
    .A1(_11840_),
    .A2(_11842_),
    .ZN(_00422_)
  );
  AND2_X1 _46382_ (
    .A1(reg_out[5]),
    .A2(_02913_),
    .ZN(_11843_)
  );
  INV_X1 _46383_ (
    .A(_11843_),
    .ZN(_11844_)
  );
  AND2_X1 _46384_ (
    .A1(_02981_),
    .A2(_11844_),
    .ZN(_11845_)
  );
  INV_X1 _46385_ (
    .A(_11845_),
    .ZN(_11846_)
  );
  AND2_X1 _46386_ (
    .A1(_11761_),
    .A2(_11846_),
    .ZN(_11847_)
  );
  INV_X1 _46387_ (
    .A(_11847_),
    .ZN(_11848_)
  );
  AND2_X1 _46388_ (
    .A1(reg_op1[5]),
    .A2(_11760_),
    .ZN(_11849_)
  );
  INV_X1 _46389_ (
    .A(_11849_),
    .ZN(_11850_)
  );
  AND2_X1 _46390_ (
    .A1(_11848_),
    .A2(_11850_),
    .ZN(_11851_)
  );
  INV_X1 _46391_ (
    .A(_11851_),
    .ZN(mem_la_addr[5])
  );
  AND2_X1 _46392_ (
    .A1(_21297_),
    .A2(_11771_),
    .ZN(_11852_)
  );
  INV_X1 _46393_ (
    .A(_11852_),
    .ZN(_11853_)
  );
  AND2_X1 _46394_ (
    .A1(_11770_),
    .A2(_11851_),
    .ZN(_11854_)
  );
  INV_X1 _46395_ (
    .A(_11854_),
    .ZN(_11855_)
  );
  AND2_X1 _46396_ (
    .A1(_11853_),
    .A2(_11855_),
    .ZN(_00423_)
  );
  AND2_X1 _46397_ (
    .A1(reg_out[6]),
    .A2(_02913_),
    .ZN(_11856_)
  );
  INV_X1 _46398_ (
    .A(_11856_),
    .ZN(_11857_)
  );
  AND2_X1 _46399_ (
    .A1(_02997_),
    .A2(_11857_),
    .ZN(_11858_)
  );
  INV_X1 _46400_ (
    .A(_11858_),
    .ZN(_11859_)
  );
  AND2_X1 _46401_ (
    .A1(_11761_),
    .A2(_11859_),
    .ZN(_11860_)
  );
  INV_X1 _46402_ (
    .A(_11860_),
    .ZN(_11861_)
  );
  AND2_X1 _46403_ (
    .A1(reg_op1[6]),
    .A2(_11760_),
    .ZN(_11862_)
  );
  INV_X1 _46404_ (
    .A(_11862_),
    .ZN(_11863_)
  );
  AND2_X1 _46405_ (
    .A1(_11861_),
    .A2(_11863_),
    .ZN(_11864_)
  );
  INV_X1 _46406_ (
    .A(_11864_),
    .ZN(mem_la_addr[6])
  );
  AND2_X1 _46407_ (
    .A1(_21298_),
    .A2(_11771_),
    .ZN(_11865_)
  );
  INV_X1 _46408_ (
    .A(_11865_),
    .ZN(_11866_)
  );
  AND2_X1 _46409_ (
    .A1(_11770_),
    .A2(_11864_),
    .ZN(_11867_)
  );
  INV_X1 _46410_ (
    .A(_11867_),
    .ZN(_11868_)
  );
  AND2_X1 _46411_ (
    .A1(_11866_),
    .A2(_11868_),
    .ZN(_00424_)
  );
  AND2_X1 _46412_ (
    .A1(reg_out[7]),
    .A2(_02913_),
    .ZN(_11869_)
  );
  INV_X1 _46413_ (
    .A(_11869_),
    .ZN(_11870_)
  );
  AND2_X1 _46414_ (
    .A1(_03013_),
    .A2(_11870_),
    .ZN(_11871_)
  );
  INV_X1 _46415_ (
    .A(_11871_),
    .ZN(_11872_)
  );
  AND2_X1 _46416_ (
    .A1(_11761_),
    .A2(_11872_),
    .ZN(_11873_)
  );
  INV_X1 _46417_ (
    .A(_11873_),
    .ZN(_11874_)
  );
  AND2_X1 _46418_ (
    .A1(reg_op1[7]),
    .A2(_11760_),
    .ZN(_11875_)
  );
  INV_X1 _46419_ (
    .A(_11875_),
    .ZN(_11876_)
  );
  AND2_X1 _46420_ (
    .A1(_11874_),
    .A2(_11876_),
    .ZN(_11877_)
  );
  INV_X1 _46421_ (
    .A(_11877_),
    .ZN(mem_la_addr[7])
  );
  AND2_X1 _46422_ (
    .A1(_21299_),
    .A2(_11771_),
    .ZN(_11878_)
  );
  INV_X1 _46423_ (
    .A(_11878_),
    .ZN(_11879_)
  );
  AND2_X1 _46424_ (
    .A1(_11770_),
    .A2(_11877_),
    .ZN(_11880_)
  );
  INV_X1 _46425_ (
    .A(_11880_),
    .ZN(_11881_)
  );
  AND2_X1 _46426_ (
    .A1(_11879_),
    .A2(_11881_),
    .ZN(_00425_)
  );
  AND2_X1 _46427_ (
    .A1(reg_out[8]),
    .A2(_02913_),
    .ZN(_11882_)
  );
  INV_X1 _46428_ (
    .A(_11882_),
    .ZN(_11883_)
  );
  AND2_X1 _46429_ (
    .A1(_03029_),
    .A2(_11883_),
    .ZN(_11884_)
  );
  INV_X1 _46430_ (
    .A(_11884_),
    .ZN(_11885_)
  );
  AND2_X1 _46431_ (
    .A1(_11761_),
    .A2(_11885_),
    .ZN(_11886_)
  );
  INV_X1 _46432_ (
    .A(_11886_),
    .ZN(_11887_)
  );
  AND2_X1 _46433_ (
    .A1(reg_op1[8]),
    .A2(_11760_),
    .ZN(_11888_)
  );
  INV_X1 _46434_ (
    .A(_11888_),
    .ZN(_11889_)
  );
  AND2_X1 _46435_ (
    .A1(_11887_),
    .A2(_11889_),
    .ZN(_11890_)
  );
  INV_X1 _46436_ (
    .A(_11890_),
    .ZN(mem_la_addr[8])
  );
  AND2_X1 _46437_ (
    .A1(_21300_),
    .A2(_11771_),
    .ZN(_11891_)
  );
  INV_X1 _46438_ (
    .A(_11891_),
    .ZN(_11892_)
  );
  AND2_X1 _46439_ (
    .A1(_11770_),
    .A2(_11890_),
    .ZN(_11893_)
  );
  INV_X1 _46440_ (
    .A(_11893_),
    .ZN(_11894_)
  );
  AND2_X1 _46441_ (
    .A1(_11892_),
    .A2(_11894_),
    .ZN(_00426_)
  );
  AND2_X1 _46442_ (
    .A1(reg_out[9]),
    .A2(_02913_),
    .ZN(_11895_)
  );
  INV_X1 _46443_ (
    .A(_11895_),
    .ZN(_11896_)
  );
  AND2_X1 _46444_ (
    .A1(_03045_),
    .A2(_11896_),
    .ZN(_11897_)
  );
  INV_X1 _46445_ (
    .A(_11897_),
    .ZN(_11898_)
  );
  AND2_X1 _46446_ (
    .A1(_11761_),
    .A2(_11898_),
    .ZN(_11899_)
  );
  INV_X1 _46447_ (
    .A(_11899_),
    .ZN(_11900_)
  );
  AND2_X1 _46448_ (
    .A1(reg_op1[9]),
    .A2(_11760_),
    .ZN(_11901_)
  );
  INV_X1 _46449_ (
    .A(_11901_),
    .ZN(_11902_)
  );
  AND2_X1 _46450_ (
    .A1(_11900_),
    .A2(_11902_),
    .ZN(_11903_)
  );
  INV_X1 _46451_ (
    .A(_11903_),
    .ZN(mem_la_addr[9])
  );
  AND2_X1 _46452_ (
    .A1(_21301_),
    .A2(_11771_),
    .ZN(_11904_)
  );
  INV_X1 _46453_ (
    .A(_11904_),
    .ZN(_11905_)
  );
  AND2_X1 _46454_ (
    .A1(_11770_),
    .A2(_11903_),
    .ZN(_11906_)
  );
  INV_X1 _46455_ (
    .A(_11906_),
    .ZN(_11907_)
  );
  AND2_X1 _46456_ (
    .A1(_11905_),
    .A2(_11907_),
    .ZN(_00427_)
  );
  AND2_X1 _46457_ (
    .A1(reg_out[10]),
    .A2(_02913_),
    .ZN(_11908_)
  );
  INV_X1 _46458_ (
    .A(_11908_),
    .ZN(_11909_)
  );
  AND2_X1 _46459_ (
    .A1(_03061_),
    .A2(_11909_),
    .ZN(_11910_)
  );
  INV_X1 _46460_ (
    .A(_11910_),
    .ZN(_11911_)
  );
  AND2_X1 _46461_ (
    .A1(_11761_),
    .A2(_11911_),
    .ZN(_11912_)
  );
  INV_X1 _46462_ (
    .A(_11912_),
    .ZN(_11913_)
  );
  AND2_X1 _46463_ (
    .A1(reg_op1[10]),
    .A2(_11760_),
    .ZN(_11914_)
  );
  INV_X1 _46464_ (
    .A(_11914_),
    .ZN(_11915_)
  );
  AND2_X1 _46465_ (
    .A1(_11913_),
    .A2(_11915_),
    .ZN(_11916_)
  );
  INV_X1 _46466_ (
    .A(_11916_),
    .ZN(mem_la_addr[10])
  );
  AND2_X1 _46467_ (
    .A1(_21302_),
    .A2(_11771_),
    .ZN(_11917_)
  );
  INV_X1 _46468_ (
    .A(_11917_),
    .ZN(_11918_)
  );
  AND2_X1 _46469_ (
    .A1(_11770_),
    .A2(_11916_),
    .ZN(_11919_)
  );
  INV_X1 _46470_ (
    .A(_11919_),
    .ZN(_11920_)
  );
  AND2_X1 _46471_ (
    .A1(_11918_),
    .A2(_11920_),
    .ZN(_00428_)
  );
  AND2_X1 _46472_ (
    .A1(reg_out[11]),
    .A2(_02913_),
    .ZN(_11921_)
  );
  INV_X1 _46473_ (
    .A(_11921_),
    .ZN(_11922_)
  );
  AND2_X1 _46474_ (
    .A1(_03077_),
    .A2(_11922_),
    .ZN(_11923_)
  );
  INV_X1 _46475_ (
    .A(_11923_),
    .ZN(_11924_)
  );
  AND2_X1 _46476_ (
    .A1(_11761_),
    .A2(_11924_),
    .ZN(_11925_)
  );
  INV_X1 _46477_ (
    .A(_11925_),
    .ZN(_11926_)
  );
  AND2_X1 _46478_ (
    .A1(reg_op1[11]),
    .A2(_11760_),
    .ZN(_11927_)
  );
  INV_X1 _46479_ (
    .A(_11927_),
    .ZN(_11928_)
  );
  AND2_X1 _46480_ (
    .A1(_11926_),
    .A2(_11928_),
    .ZN(_11929_)
  );
  INV_X1 _46481_ (
    .A(_11929_),
    .ZN(mem_la_addr[11])
  );
  AND2_X1 _46482_ (
    .A1(_21303_),
    .A2(_11771_),
    .ZN(_11930_)
  );
  INV_X1 _46483_ (
    .A(_11930_),
    .ZN(_11931_)
  );
  AND2_X1 _46484_ (
    .A1(_11770_),
    .A2(_11929_),
    .ZN(_11932_)
  );
  INV_X1 _46485_ (
    .A(_11932_),
    .ZN(_11933_)
  );
  AND2_X1 _46486_ (
    .A1(_11931_),
    .A2(_11933_),
    .ZN(_00429_)
  );
  AND2_X1 _46487_ (
    .A1(reg_out[12]),
    .A2(_02913_),
    .ZN(_11934_)
  );
  INV_X1 _46488_ (
    .A(_11934_),
    .ZN(_11935_)
  );
  AND2_X1 _46489_ (
    .A1(_03093_),
    .A2(_11935_),
    .ZN(_11936_)
  );
  INV_X1 _46490_ (
    .A(_11936_),
    .ZN(_11937_)
  );
  AND2_X1 _46491_ (
    .A1(_11761_),
    .A2(_11937_),
    .ZN(_11938_)
  );
  INV_X1 _46492_ (
    .A(_11938_),
    .ZN(_11939_)
  );
  AND2_X1 _46493_ (
    .A1(reg_op1[12]),
    .A2(_11760_),
    .ZN(_11940_)
  );
  INV_X1 _46494_ (
    .A(_11940_),
    .ZN(_11941_)
  );
  AND2_X1 _46495_ (
    .A1(_11939_),
    .A2(_11941_),
    .ZN(_11942_)
  );
  INV_X1 _46496_ (
    .A(_11942_),
    .ZN(mem_la_addr[12])
  );
  AND2_X1 _46497_ (
    .A1(_21304_),
    .A2(_11771_),
    .ZN(_11943_)
  );
  INV_X1 _46498_ (
    .A(_11943_),
    .ZN(_11944_)
  );
  AND2_X1 _46499_ (
    .A1(_11770_),
    .A2(_11942_),
    .ZN(_11945_)
  );
  INV_X1 _46500_ (
    .A(_11945_),
    .ZN(_11946_)
  );
  AND2_X1 _46501_ (
    .A1(_11944_),
    .A2(_11946_),
    .ZN(_00430_)
  );
  AND2_X1 _46502_ (
    .A1(reg_out[13]),
    .A2(_02913_),
    .ZN(_11947_)
  );
  INV_X1 _46503_ (
    .A(_11947_),
    .ZN(_11948_)
  );
  AND2_X1 _46504_ (
    .A1(_03109_),
    .A2(_11948_),
    .ZN(_11949_)
  );
  INV_X1 _46505_ (
    .A(_11949_),
    .ZN(_11950_)
  );
  AND2_X1 _46506_ (
    .A1(_11761_),
    .A2(_11950_),
    .ZN(_11951_)
  );
  INV_X1 _46507_ (
    .A(_11951_),
    .ZN(_11952_)
  );
  AND2_X1 _46508_ (
    .A1(reg_op1[13]),
    .A2(_11760_),
    .ZN(_11953_)
  );
  INV_X1 _46509_ (
    .A(_11953_),
    .ZN(_11954_)
  );
  AND2_X1 _46510_ (
    .A1(_11952_),
    .A2(_11954_),
    .ZN(_11955_)
  );
  INV_X1 _46511_ (
    .A(_11955_),
    .ZN(mem_la_addr[13])
  );
  AND2_X1 _46512_ (
    .A1(_21305_),
    .A2(_11771_),
    .ZN(_11956_)
  );
  INV_X1 _46513_ (
    .A(_11956_),
    .ZN(_11957_)
  );
  AND2_X1 _46514_ (
    .A1(_11770_),
    .A2(_11955_),
    .ZN(_11958_)
  );
  INV_X1 _46515_ (
    .A(_11958_),
    .ZN(_11959_)
  );
  AND2_X1 _46516_ (
    .A1(_11957_),
    .A2(_11959_),
    .ZN(_00431_)
  );
  AND2_X1 _46517_ (
    .A1(reg_out[14]),
    .A2(_02913_),
    .ZN(_11960_)
  );
  INV_X1 _46518_ (
    .A(_11960_),
    .ZN(_11961_)
  );
  AND2_X1 _46519_ (
    .A1(_03125_),
    .A2(_11961_),
    .ZN(_11962_)
  );
  INV_X1 _46520_ (
    .A(_11962_),
    .ZN(_11963_)
  );
  AND2_X1 _46521_ (
    .A1(_11761_),
    .A2(_11963_),
    .ZN(_11964_)
  );
  INV_X1 _46522_ (
    .A(_11964_),
    .ZN(_11965_)
  );
  AND2_X1 _46523_ (
    .A1(reg_op1[14]),
    .A2(_11760_),
    .ZN(_11966_)
  );
  INV_X1 _46524_ (
    .A(_11966_),
    .ZN(_11967_)
  );
  AND2_X1 _46525_ (
    .A1(_11965_),
    .A2(_11967_),
    .ZN(_11968_)
  );
  INV_X1 _46526_ (
    .A(_11968_),
    .ZN(mem_la_addr[14])
  );
  AND2_X1 _46527_ (
    .A1(_21306_),
    .A2(_11771_),
    .ZN(_11969_)
  );
  INV_X1 _46528_ (
    .A(_11969_),
    .ZN(_11970_)
  );
  AND2_X1 _46529_ (
    .A1(_11770_),
    .A2(_11968_),
    .ZN(_11971_)
  );
  INV_X1 _46530_ (
    .A(_11971_),
    .ZN(_11972_)
  );
  AND2_X1 _46531_ (
    .A1(_11970_),
    .A2(_11972_),
    .ZN(_00432_)
  );
  AND2_X1 _46532_ (
    .A1(reg_out[15]),
    .A2(_02913_),
    .ZN(_11973_)
  );
  INV_X1 _46533_ (
    .A(_11973_),
    .ZN(_11974_)
  );
  AND2_X1 _46534_ (
    .A1(_03141_),
    .A2(_11974_),
    .ZN(_11975_)
  );
  INV_X1 _46535_ (
    .A(_11975_),
    .ZN(_11976_)
  );
  AND2_X1 _46536_ (
    .A1(_11761_),
    .A2(_11976_),
    .ZN(_11977_)
  );
  INV_X1 _46537_ (
    .A(_11977_),
    .ZN(_11978_)
  );
  AND2_X1 _46538_ (
    .A1(reg_op1[15]),
    .A2(_11760_),
    .ZN(_11979_)
  );
  INV_X1 _46539_ (
    .A(_11979_),
    .ZN(_11980_)
  );
  AND2_X1 _46540_ (
    .A1(_11978_),
    .A2(_11980_),
    .ZN(_11981_)
  );
  INV_X1 _46541_ (
    .A(_11981_),
    .ZN(mem_la_addr[15])
  );
  AND2_X1 _46542_ (
    .A1(_21307_),
    .A2(_11771_),
    .ZN(_11982_)
  );
  INV_X1 _46543_ (
    .A(_11982_),
    .ZN(_11983_)
  );
  AND2_X1 _46544_ (
    .A1(_11770_),
    .A2(_11981_),
    .ZN(_11984_)
  );
  INV_X1 _46545_ (
    .A(_11984_),
    .ZN(_11985_)
  );
  AND2_X1 _46546_ (
    .A1(_11983_),
    .A2(_11985_),
    .ZN(_00433_)
  );
  AND2_X1 _46547_ (
    .A1(reg_out[16]),
    .A2(_02913_),
    .ZN(_11986_)
  );
  INV_X1 _46548_ (
    .A(_11986_),
    .ZN(_11987_)
  );
  AND2_X1 _46549_ (
    .A1(_03157_),
    .A2(_11987_),
    .ZN(_11988_)
  );
  INV_X1 _46550_ (
    .A(_11988_),
    .ZN(_11989_)
  );
  AND2_X1 _46551_ (
    .A1(_11761_),
    .A2(_11989_),
    .ZN(_11990_)
  );
  INV_X1 _46552_ (
    .A(_11990_),
    .ZN(_11991_)
  );
  AND2_X1 _46553_ (
    .A1(reg_op1[16]),
    .A2(_11760_),
    .ZN(_11992_)
  );
  INV_X1 _46554_ (
    .A(_11992_),
    .ZN(_11993_)
  );
  AND2_X1 _46555_ (
    .A1(_11991_),
    .A2(_11993_),
    .ZN(_11994_)
  );
  INV_X1 _46556_ (
    .A(_11994_),
    .ZN(mem_la_addr[16])
  );
  AND2_X1 _46557_ (
    .A1(_21308_),
    .A2(_11771_),
    .ZN(_11995_)
  );
  INV_X1 _46558_ (
    .A(_11995_),
    .ZN(_11996_)
  );
  AND2_X1 _46559_ (
    .A1(_11770_),
    .A2(_11994_),
    .ZN(_11997_)
  );
  INV_X1 _46560_ (
    .A(_11997_),
    .ZN(_11998_)
  );
  AND2_X1 _46561_ (
    .A1(_11996_),
    .A2(_11998_),
    .ZN(_00434_)
  );
  AND2_X1 _46562_ (
    .A1(reg_out[17]),
    .A2(_02913_),
    .ZN(_11999_)
  );
  INV_X1 _46563_ (
    .A(_11999_),
    .ZN(_12000_)
  );
  AND2_X1 _46564_ (
    .A1(_03173_),
    .A2(_12000_),
    .ZN(_12001_)
  );
  INV_X1 _46565_ (
    .A(_12001_),
    .ZN(_12002_)
  );
  AND2_X1 _46566_ (
    .A1(_11761_),
    .A2(_12002_),
    .ZN(_12003_)
  );
  INV_X1 _46567_ (
    .A(_12003_),
    .ZN(_12004_)
  );
  AND2_X1 _46568_ (
    .A1(reg_op1[17]),
    .A2(_11760_),
    .ZN(_12005_)
  );
  INV_X1 _46569_ (
    .A(_12005_),
    .ZN(_12006_)
  );
  AND2_X1 _46570_ (
    .A1(_12004_),
    .A2(_12006_),
    .ZN(_12007_)
  );
  INV_X1 _46571_ (
    .A(_12007_),
    .ZN(mem_la_addr[17])
  );
  AND2_X1 _46572_ (
    .A1(_21309_),
    .A2(_11771_),
    .ZN(_12008_)
  );
  INV_X1 _46573_ (
    .A(_12008_),
    .ZN(_12009_)
  );
  AND2_X1 _46574_ (
    .A1(_11770_),
    .A2(_12007_),
    .ZN(_12010_)
  );
  INV_X1 _46575_ (
    .A(_12010_),
    .ZN(_12011_)
  );
  AND2_X1 _46576_ (
    .A1(_12009_),
    .A2(_12011_),
    .ZN(_00435_)
  );
  AND2_X1 _46577_ (
    .A1(reg_out[18]),
    .A2(_02913_),
    .ZN(_12012_)
  );
  INV_X1 _46578_ (
    .A(_12012_),
    .ZN(_12013_)
  );
  AND2_X1 _46579_ (
    .A1(_03189_),
    .A2(_12013_),
    .ZN(_12014_)
  );
  INV_X1 _46580_ (
    .A(_12014_),
    .ZN(_12015_)
  );
  AND2_X1 _46581_ (
    .A1(_11761_),
    .A2(_12015_),
    .ZN(_12016_)
  );
  INV_X1 _46582_ (
    .A(_12016_),
    .ZN(_12017_)
  );
  AND2_X1 _46583_ (
    .A1(reg_op1[18]),
    .A2(_11760_),
    .ZN(_12018_)
  );
  INV_X1 _46584_ (
    .A(_12018_),
    .ZN(_12019_)
  );
  AND2_X1 _46585_ (
    .A1(_12017_),
    .A2(_12019_),
    .ZN(_12020_)
  );
  INV_X1 _46586_ (
    .A(_12020_),
    .ZN(mem_la_addr[18])
  );
  AND2_X1 _46587_ (
    .A1(_21310_),
    .A2(_11771_),
    .ZN(_12021_)
  );
  INV_X1 _46588_ (
    .A(_12021_),
    .ZN(_12022_)
  );
  AND2_X1 _46589_ (
    .A1(_11770_),
    .A2(_12020_),
    .ZN(_12023_)
  );
  INV_X1 _46590_ (
    .A(_12023_),
    .ZN(_12024_)
  );
  AND2_X1 _46591_ (
    .A1(_12022_),
    .A2(_12024_),
    .ZN(_00436_)
  );
  AND2_X1 _46592_ (
    .A1(reg_out[19]),
    .A2(_02913_),
    .ZN(_12025_)
  );
  INV_X1 _46593_ (
    .A(_12025_),
    .ZN(_12026_)
  );
  AND2_X1 _46594_ (
    .A1(_03205_),
    .A2(_12026_),
    .ZN(_12027_)
  );
  INV_X1 _46595_ (
    .A(_12027_),
    .ZN(_12028_)
  );
  AND2_X1 _46596_ (
    .A1(_11761_),
    .A2(_12028_),
    .ZN(_12029_)
  );
  INV_X1 _46597_ (
    .A(_12029_),
    .ZN(_12030_)
  );
  AND2_X1 _46598_ (
    .A1(reg_op1[19]),
    .A2(_11760_),
    .ZN(_12031_)
  );
  INV_X1 _46599_ (
    .A(_12031_),
    .ZN(_12032_)
  );
  AND2_X1 _46600_ (
    .A1(_12030_),
    .A2(_12032_),
    .ZN(_12033_)
  );
  INV_X1 _46601_ (
    .A(_12033_),
    .ZN(mem_la_addr[19])
  );
  AND2_X1 _46602_ (
    .A1(_21311_),
    .A2(_11771_),
    .ZN(_12034_)
  );
  INV_X1 _46603_ (
    .A(_12034_),
    .ZN(_12035_)
  );
  AND2_X1 _46604_ (
    .A1(_11770_),
    .A2(_12033_),
    .ZN(_12036_)
  );
  INV_X1 _46605_ (
    .A(_12036_),
    .ZN(_12037_)
  );
  AND2_X1 _46606_ (
    .A1(_12035_),
    .A2(_12037_),
    .ZN(_00437_)
  );
  AND2_X1 _46607_ (
    .A1(reg_out[20]),
    .A2(_02913_),
    .ZN(_12038_)
  );
  INV_X1 _46608_ (
    .A(_12038_),
    .ZN(_12039_)
  );
  AND2_X1 _46609_ (
    .A1(_03221_),
    .A2(_12039_),
    .ZN(_12040_)
  );
  INV_X1 _46610_ (
    .A(_12040_),
    .ZN(_12041_)
  );
  AND2_X1 _46611_ (
    .A1(_11761_),
    .A2(_12041_),
    .ZN(_12042_)
  );
  INV_X1 _46612_ (
    .A(_12042_),
    .ZN(_12043_)
  );
  AND2_X1 _46613_ (
    .A1(reg_op1[20]),
    .A2(_11760_),
    .ZN(_12044_)
  );
  INV_X1 _46614_ (
    .A(_12044_),
    .ZN(_12045_)
  );
  AND2_X1 _46615_ (
    .A1(_12043_),
    .A2(_12045_),
    .ZN(_12046_)
  );
  INV_X1 _46616_ (
    .A(_12046_),
    .ZN(mem_la_addr[20])
  );
  AND2_X1 _46617_ (
    .A1(_21312_),
    .A2(_11771_),
    .ZN(_12047_)
  );
  INV_X1 _46618_ (
    .A(_12047_),
    .ZN(_12048_)
  );
  AND2_X1 _46619_ (
    .A1(_11770_),
    .A2(_12046_),
    .ZN(_12049_)
  );
  INV_X1 _46620_ (
    .A(_12049_),
    .ZN(_12050_)
  );
  AND2_X1 _46621_ (
    .A1(_12048_),
    .A2(_12050_),
    .ZN(_00438_)
  );
  AND2_X1 _46622_ (
    .A1(reg_out[21]),
    .A2(_02913_),
    .ZN(_12051_)
  );
  INV_X1 _46623_ (
    .A(_12051_),
    .ZN(_12052_)
  );
  AND2_X1 _46624_ (
    .A1(_03237_),
    .A2(_12052_),
    .ZN(_12053_)
  );
  INV_X1 _46625_ (
    .A(_12053_),
    .ZN(_12054_)
  );
  AND2_X1 _46626_ (
    .A1(_11761_),
    .A2(_12054_),
    .ZN(_12055_)
  );
  INV_X1 _46627_ (
    .A(_12055_),
    .ZN(_12056_)
  );
  AND2_X1 _46628_ (
    .A1(reg_op1[21]),
    .A2(_11760_),
    .ZN(_12057_)
  );
  INV_X1 _46629_ (
    .A(_12057_),
    .ZN(_12058_)
  );
  AND2_X1 _46630_ (
    .A1(_12056_),
    .A2(_12058_),
    .ZN(_12059_)
  );
  INV_X1 _46631_ (
    .A(_12059_),
    .ZN(mem_la_addr[21])
  );
  AND2_X1 _46632_ (
    .A1(_21313_),
    .A2(_11771_),
    .ZN(_12060_)
  );
  INV_X1 _46633_ (
    .A(_12060_),
    .ZN(_12061_)
  );
  AND2_X1 _46634_ (
    .A1(_11770_),
    .A2(_12059_),
    .ZN(_12062_)
  );
  INV_X1 _46635_ (
    .A(_12062_),
    .ZN(_12063_)
  );
  AND2_X1 _46636_ (
    .A1(_12061_),
    .A2(_12063_),
    .ZN(_00439_)
  );
  AND2_X1 _46637_ (
    .A1(reg_out[22]),
    .A2(_02913_),
    .ZN(_12064_)
  );
  INV_X1 _46638_ (
    .A(_12064_),
    .ZN(_12065_)
  );
  AND2_X1 _46639_ (
    .A1(_03253_),
    .A2(_12065_),
    .ZN(_12066_)
  );
  INV_X1 _46640_ (
    .A(_12066_),
    .ZN(_12067_)
  );
  AND2_X1 _46641_ (
    .A1(_11761_),
    .A2(_12067_),
    .ZN(_12068_)
  );
  INV_X1 _46642_ (
    .A(_12068_),
    .ZN(_12069_)
  );
  AND2_X1 _46643_ (
    .A1(reg_op1[22]),
    .A2(_11760_),
    .ZN(_12070_)
  );
  INV_X1 _46644_ (
    .A(_12070_),
    .ZN(_12071_)
  );
  AND2_X1 _46645_ (
    .A1(_12069_),
    .A2(_12071_),
    .ZN(_12072_)
  );
  INV_X1 _46646_ (
    .A(_12072_),
    .ZN(mem_la_addr[22])
  );
  AND2_X1 _46647_ (
    .A1(_21314_),
    .A2(_11771_),
    .ZN(_12073_)
  );
  INV_X1 _46648_ (
    .A(_12073_),
    .ZN(_12074_)
  );
  AND2_X1 _46649_ (
    .A1(_11770_),
    .A2(_12072_),
    .ZN(_12075_)
  );
  INV_X1 _46650_ (
    .A(_12075_),
    .ZN(_12076_)
  );
  AND2_X1 _46651_ (
    .A1(_12074_),
    .A2(_12076_),
    .ZN(_00440_)
  );
  AND2_X1 _46652_ (
    .A1(reg_out[23]),
    .A2(_02913_),
    .ZN(_12077_)
  );
  INV_X1 _46653_ (
    .A(_12077_),
    .ZN(_12078_)
  );
  AND2_X1 _46654_ (
    .A1(_03269_),
    .A2(_12078_),
    .ZN(_12079_)
  );
  INV_X1 _46655_ (
    .A(_12079_),
    .ZN(_12080_)
  );
  AND2_X1 _46656_ (
    .A1(_11761_),
    .A2(_12080_),
    .ZN(_12081_)
  );
  INV_X1 _46657_ (
    .A(_12081_),
    .ZN(_12082_)
  );
  AND2_X1 _46658_ (
    .A1(reg_op1[23]),
    .A2(_11760_),
    .ZN(_12083_)
  );
  INV_X1 _46659_ (
    .A(_12083_),
    .ZN(_12084_)
  );
  AND2_X1 _46660_ (
    .A1(_12082_),
    .A2(_12084_),
    .ZN(_12085_)
  );
  INV_X1 _46661_ (
    .A(_12085_),
    .ZN(mem_la_addr[23])
  );
  AND2_X1 _46662_ (
    .A1(_21315_),
    .A2(_11771_),
    .ZN(_12086_)
  );
  INV_X1 _46663_ (
    .A(_12086_),
    .ZN(_12087_)
  );
  AND2_X1 _46664_ (
    .A1(_11770_),
    .A2(_12085_),
    .ZN(_12088_)
  );
  INV_X1 _46665_ (
    .A(_12088_),
    .ZN(_12089_)
  );
  AND2_X1 _46666_ (
    .A1(_12087_),
    .A2(_12089_),
    .ZN(_00441_)
  );
  AND2_X1 _46667_ (
    .A1(reg_out[24]),
    .A2(_02913_),
    .ZN(_12090_)
  );
  INV_X1 _46668_ (
    .A(_12090_),
    .ZN(_12091_)
  );
  AND2_X1 _46669_ (
    .A1(_03285_),
    .A2(_12091_),
    .ZN(_12092_)
  );
  INV_X1 _46670_ (
    .A(_12092_),
    .ZN(_12093_)
  );
  AND2_X1 _46671_ (
    .A1(_11761_),
    .A2(_12093_),
    .ZN(_12094_)
  );
  INV_X1 _46672_ (
    .A(_12094_),
    .ZN(_12095_)
  );
  AND2_X1 _46673_ (
    .A1(reg_op1[24]),
    .A2(_11760_),
    .ZN(_12096_)
  );
  INV_X1 _46674_ (
    .A(_12096_),
    .ZN(_12097_)
  );
  AND2_X1 _46675_ (
    .A1(_12095_),
    .A2(_12097_),
    .ZN(_12098_)
  );
  INV_X1 _46676_ (
    .A(_12098_),
    .ZN(mem_la_addr[24])
  );
  AND2_X1 _46677_ (
    .A1(_21316_),
    .A2(_11771_),
    .ZN(_12099_)
  );
  INV_X1 _46678_ (
    .A(_12099_),
    .ZN(_12100_)
  );
  AND2_X1 _46679_ (
    .A1(_11770_),
    .A2(_12098_),
    .ZN(_12101_)
  );
  INV_X1 _46680_ (
    .A(_12101_),
    .ZN(_12102_)
  );
  AND2_X1 _46681_ (
    .A1(_12100_),
    .A2(_12102_),
    .ZN(_00442_)
  );
  AND2_X1 _46682_ (
    .A1(reg_out[25]),
    .A2(_02913_),
    .ZN(_12103_)
  );
  INV_X1 _46683_ (
    .A(_12103_),
    .ZN(_12104_)
  );
  AND2_X1 _46684_ (
    .A1(_03301_),
    .A2(_12104_),
    .ZN(_12105_)
  );
  INV_X1 _46685_ (
    .A(_12105_),
    .ZN(_12106_)
  );
  AND2_X1 _46686_ (
    .A1(_11761_),
    .A2(_12106_),
    .ZN(_12107_)
  );
  INV_X1 _46687_ (
    .A(_12107_),
    .ZN(_12108_)
  );
  AND2_X1 _46688_ (
    .A1(reg_op1[25]),
    .A2(_11760_),
    .ZN(_12109_)
  );
  INV_X1 _46689_ (
    .A(_12109_),
    .ZN(_12110_)
  );
  AND2_X1 _46690_ (
    .A1(_12108_),
    .A2(_12110_),
    .ZN(_12111_)
  );
  INV_X1 _46691_ (
    .A(_12111_),
    .ZN(mem_la_addr[25])
  );
  AND2_X1 _46692_ (
    .A1(_21317_),
    .A2(_11771_),
    .ZN(_12112_)
  );
  INV_X1 _46693_ (
    .A(_12112_),
    .ZN(_12113_)
  );
  AND2_X1 _46694_ (
    .A1(_11770_),
    .A2(_12111_),
    .ZN(_12114_)
  );
  INV_X1 _46695_ (
    .A(_12114_),
    .ZN(_12115_)
  );
  AND2_X1 _46696_ (
    .A1(_12113_),
    .A2(_12115_),
    .ZN(_00443_)
  );
  AND2_X1 _46697_ (
    .A1(reg_out[26]),
    .A2(_02913_),
    .ZN(_12116_)
  );
  INV_X1 _46698_ (
    .A(_12116_),
    .ZN(_12117_)
  );
  AND2_X1 _46699_ (
    .A1(_03317_),
    .A2(_12117_),
    .ZN(_12118_)
  );
  INV_X1 _46700_ (
    .A(_12118_),
    .ZN(_12119_)
  );
  AND2_X1 _46701_ (
    .A1(_11761_),
    .A2(_12119_),
    .ZN(_12120_)
  );
  INV_X1 _46702_ (
    .A(_12120_),
    .ZN(_12121_)
  );
  AND2_X1 _46703_ (
    .A1(reg_op1[26]),
    .A2(_11760_),
    .ZN(_12122_)
  );
  INV_X1 _46704_ (
    .A(_12122_),
    .ZN(_12123_)
  );
  AND2_X1 _46705_ (
    .A1(_12121_),
    .A2(_12123_),
    .ZN(_12124_)
  );
  INV_X1 _46706_ (
    .A(_12124_),
    .ZN(mem_la_addr[26])
  );
  AND2_X1 _46707_ (
    .A1(_21318_),
    .A2(_11771_),
    .ZN(_12125_)
  );
  INV_X1 _46708_ (
    .A(_12125_),
    .ZN(_12126_)
  );
  AND2_X1 _46709_ (
    .A1(_11770_),
    .A2(_12124_),
    .ZN(_12127_)
  );
  INV_X1 _46710_ (
    .A(_12127_),
    .ZN(_12128_)
  );
  AND2_X1 _46711_ (
    .A1(_12126_),
    .A2(_12128_),
    .ZN(_00444_)
  );
  AND2_X1 _46712_ (
    .A1(reg_out[27]),
    .A2(_02913_),
    .ZN(_12129_)
  );
  INV_X1 _46713_ (
    .A(_12129_),
    .ZN(_12130_)
  );
  AND2_X1 _46714_ (
    .A1(_03333_),
    .A2(_12130_),
    .ZN(_12131_)
  );
  INV_X1 _46715_ (
    .A(_12131_),
    .ZN(_12132_)
  );
  AND2_X1 _46716_ (
    .A1(_11761_),
    .A2(_12132_),
    .ZN(_12133_)
  );
  INV_X1 _46717_ (
    .A(_12133_),
    .ZN(_12134_)
  );
  AND2_X1 _46718_ (
    .A1(reg_op1[27]),
    .A2(_11760_),
    .ZN(_12135_)
  );
  INV_X1 _46719_ (
    .A(_12135_),
    .ZN(_12136_)
  );
  AND2_X1 _46720_ (
    .A1(_12134_),
    .A2(_12136_),
    .ZN(_12137_)
  );
  INV_X1 _46721_ (
    .A(_12137_),
    .ZN(mem_la_addr[27])
  );
  AND2_X1 _46722_ (
    .A1(_21319_),
    .A2(_11771_),
    .ZN(_12138_)
  );
  INV_X1 _46723_ (
    .A(_12138_),
    .ZN(_12139_)
  );
  AND2_X1 _46724_ (
    .A1(_11770_),
    .A2(_12137_),
    .ZN(_12140_)
  );
  INV_X1 _46725_ (
    .A(_12140_),
    .ZN(_12141_)
  );
  AND2_X1 _46726_ (
    .A1(_12139_),
    .A2(_12141_),
    .ZN(_00445_)
  );
  AND2_X1 _46727_ (
    .A1(reg_out[28]),
    .A2(_02913_),
    .ZN(_12142_)
  );
  INV_X1 _46728_ (
    .A(_12142_),
    .ZN(_12143_)
  );
  AND2_X1 _46729_ (
    .A1(_03349_),
    .A2(_12143_),
    .ZN(_12144_)
  );
  INV_X1 _46730_ (
    .A(_12144_),
    .ZN(_12145_)
  );
  AND2_X1 _46731_ (
    .A1(_11761_),
    .A2(_12145_),
    .ZN(_12146_)
  );
  INV_X1 _46732_ (
    .A(_12146_),
    .ZN(_12147_)
  );
  AND2_X1 _46733_ (
    .A1(reg_op1[28]),
    .A2(_11760_),
    .ZN(_12148_)
  );
  INV_X1 _46734_ (
    .A(_12148_),
    .ZN(_12149_)
  );
  AND2_X1 _46735_ (
    .A1(_12147_),
    .A2(_12149_),
    .ZN(_12150_)
  );
  INV_X1 _46736_ (
    .A(_12150_),
    .ZN(mem_la_addr[28])
  );
  AND2_X1 _46737_ (
    .A1(_21320_),
    .A2(_11771_),
    .ZN(_12151_)
  );
  INV_X1 _46738_ (
    .A(_12151_),
    .ZN(_12152_)
  );
  AND2_X1 _46739_ (
    .A1(_11770_),
    .A2(_12150_),
    .ZN(_12153_)
  );
  INV_X1 _46740_ (
    .A(_12153_),
    .ZN(_12154_)
  );
  AND2_X1 _46741_ (
    .A1(_12152_),
    .A2(_12154_),
    .ZN(_00446_)
  );
  AND2_X1 _46742_ (
    .A1(reg_out[29]),
    .A2(_02913_),
    .ZN(_12155_)
  );
  INV_X1 _46743_ (
    .A(_12155_),
    .ZN(_12156_)
  );
  AND2_X1 _46744_ (
    .A1(_03365_),
    .A2(_12156_),
    .ZN(_12157_)
  );
  INV_X1 _46745_ (
    .A(_12157_),
    .ZN(_12158_)
  );
  AND2_X1 _46746_ (
    .A1(_11761_),
    .A2(_12158_),
    .ZN(_12159_)
  );
  INV_X1 _46747_ (
    .A(_12159_),
    .ZN(_12160_)
  );
  AND2_X1 _46748_ (
    .A1(reg_op1[29]),
    .A2(_11760_),
    .ZN(_12161_)
  );
  INV_X1 _46749_ (
    .A(_12161_),
    .ZN(_12162_)
  );
  AND2_X1 _46750_ (
    .A1(_12160_),
    .A2(_12162_),
    .ZN(_12163_)
  );
  INV_X1 _46751_ (
    .A(_12163_),
    .ZN(mem_la_addr[29])
  );
  AND2_X1 _46752_ (
    .A1(_21321_),
    .A2(_11771_),
    .ZN(_12164_)
  );
  INV_X1 _46753_ (
    .A(_12164_),
    .ZN(_12165_)
  );
  AND2_X1 _46754_ (
    .A1(_11770_),
    .A2(_12163_),
    .ZN(_12166_)
  );
  INV_X1 _46755_ (
    .A(_12166_),
    .ZN(_12167_)
  );
  AND2_X1 _46756_ (
    .A1(_12165_),
    .A2(_12167_),
    .ZN(_00447_)
  );
  AND2_X1 _46757_ (
    .A1(reg_out[30]),
    .A2(_02913_),
    .ZN(_12168_)
  );
  INV_X1 _46758_ (
    .A(_12168_),
    .ZN(_12169_)
  );
  AND2_X1 _46759_ (
    .A1(_03381_),
    .A2(_12169_),
    .ZN(_12170_)
  );
  INV_X1 _46760_ (
    .A(_12170_),
    .ZN(_12171_)
  );
  AND2_X1 _46761_ (
    .A1(_11761_),
    .A2(_12171_),
    .ZN(_12172_)
  );
  INV_X1 _46762_ (
    .A(_12172_),
    .ZN(_12173_)
  );
  AND2_X1 _46763_ (
    .A1(reg_op1[30]),
    .A2(_11760_),
    .ZN(_12174_)
  );
  INV_X1 _46764_ (
    .A(_12174_),
    .ZN(_12175_)
  );
  AND2_X1 _46765_ (
    .A1(_12173_),
    .A2(_12175_),
    .ZN(_12176_)
  );
  INV_X1 _46766_ (
    .A(_12176_),
    .ZN(mem_la_addr[30])
  );
  AND2_X1 _46767_ (
    .A1(_21322_),
    .A2(_11771_),
    .ZN(_12177_)
  );
  INV_X1 _46768_ (
    .A(_12177_),
    .ZN(_12178_)
  );
  AND2_X1 _46769_ (
    .A1(_11770_),
    .A2(_12176_),
    .ZN(_12179_)
  );
  INV_X1 _46770_ (
    .A(_12179_),
    .ZN(_12180_)
  );
  AND2_X1 _46771_ (
    .A1(_12178_),
    .A2(_12180_),
    .ZN(_00448_)
  );
  AND2_X1 _46772_ (
    .A1(reg_out[31]),
    .A2(_02913_),
    .ZN(_12181_)
  );
  INV_X1 _46773_ (
    .A(_12181_),
    .ZN(_12182_)
  );
  AND2_X1 _46774_ (
    .A1(_03397_),
    .A2(_12182_),
    .ZN(_12183_)
  );
  INV_X1 _46775_ (
    .A(_12183_),
    .ZN(_12184_)
  );
  AND2_X1 _46776_ (
    .A1(_11761_),
    .A2(_12184_),
    .ZN(_12185_)
  );
  INV_X1 _46777_ (
    .A(_12185_),
    .ZN(_12186_)
  );
  AND2_X1 _46778_ (
    .A1(reg_op1[31]),
    .A2(_11760_),
    .ZN(_12187_)
  );
  INV_X1 _46779_ (
    .A(_12187_),
    .ZN(_12188_)
  );
  AND2_X1 _46780_ (
    .A1(_12186_),
    .A2(_12188_),
    .ZN(_12189_)
  );
  INV_X1 _46781_ (
    .A(_12189_),
    .ZN(mem_la_addr[31])
  );
  AND2_X1 _46782_ (
    .A1(_21323_),
    .A2(_11771_),
    .ZN(_12190_)
  );
  INV_X1 _46783_ (
    .A(_12190_),
    .ZN(_12191_)
  );
  AND2_X1 _46784_ (
    .A1(_11770_),
    .A2(_12189_),
    .ZN(_12192_)
  );
  INV_X1 _46785_ (
    .A(_12192_),
    .ZN(_12193_)
  );
  AND2_X1 _46786_ (
    .A1(_12191_),
    .A2(_12193_),
    .ZN(_00449_)
  );
  AND2_X1 _46787_ (
    .A1(_21252_),
    .A2(_21253_),
    .ZN(_12194_)
  );
  INV_X1 _46788_ (
    .A(_12194_),
    .ZN(_12195_)
  );
  AND2_X1 _46789_ (
    .A1(_21252_),
    .A2(_22066_),
    .ZN(_12196_)
  );
  INV_X1 _46790_ (
    .A(_12196_),
    .ZN(_12197_)
  );
  AND2_X1 _46791_ (
    .A1(_21253_),
    .A2(_22065_),
    .ZN(_12198_)
  );
  INV_X1 _46792_ (
    .A(_12198_),
    .ZN(_12199_)
  );
  AND2_X1 _46793_ (
    .A1(_12197_),
    .A2(_12199_),
    .ZN(_12200_)
  );
  INV_X1 _46794_ (
    .A(_12200_),
    .ZN(_12201_)
  );
  AND2_X1 _46795_ (
    .A1(_12195_),
    .A2(_12200_),
    .ZN(_12202_)
  );
  INV_X1 _46796_ (
    .A(_12202_),
    .ZN(_12203_)
  );
  AND2_X1 _46797_ (
    .A1(reg_op2[0]),
    .A2(_12203_),
    .ZN(mem_la_wdata[0])
  );
  AND2_X1 _46798_ (
    .A1(mem_do_wdata),
    .A2(_11768_),
    .ZN(_12204_)
  );
  INV_X1 _46799_ (
    .A(_12204_),
    .ZN(_12205_)
  );
  AND2_X1 _46800_ (
    .A1(mem_la_wdata[0]),
    .A2(_12204_),
    .ZN(_12206_)
  );
  INV_X1 _46801_ (
    .A(_12206_),
    .ZN(_12207_)
  );
  AND2_X1 _46802_ (
    .A1(mem_wdata[0]),
    .A2(_12205_),
    .ZN(_12208_)
  );
  INV_X1 _46803_ (
    .A(_12208_),
    .ZN(_12209_)
  );
  AND2_X1 _46804_ (
    .A1(_12207_),
    .A2(_12209_),
    .ZN(_12210_)
  );
  INV_X1 _46805_ (
    .A(_12210_),
    .ZN(_00450_)
  );
  AND2_X1 _46806_ (
    .A1(reg_op2[1]),
    .A2(_12203_),
    .ZN(mem_la_wdata[1])
  );
  AND2_X1 _46807_ (
    .A1(_12204_),
    .A2(mem_la_wdata[1]),
    .ZN(_12211_)
  );
  INV_X1 _46808_ (
    .A(_12211_),
    .ZN(_12212_)
  );
  AND2_X1 _46809_ (
    .A1(mem_wdata[1]),
    .A2(_12205_),
    .ZN(_12213_)
  );
  INV_X1 _46810_ (
    .A(_12213_),
    .ZN(_12214_)
  );
  AND2_X1 _46811_ (
    .A1(_12212_),
    .A2(_12214_),
    .ZN(_12215_)
  );
  INV_X1 _46812_ (
    .A(_12215_),
    .ZN(_00451_)
  );
  AND2_X1 _46813_ (
    .A1(reg_op2[2]),
    .A2(_12203_),
    .ZN(mem_la_wdata[2])
  );
  AND2_X1 _46814_ (
    .A1(_12204_),
    .A2(mem_la_wdata[2]),
    .ZN(_12216_)
  );
  INV_X1 _46815_ (
    .A(_12216_),
    .ZN(_12217_)
  );
  AND2_X1 _46816_ (
    .A1(mem_wdata[2]),
    .A2(_12205_),
    .ZN(_12218_)
  );
  INV_X1 _46817_ (
    .A(_12218_),
    .ZN(_12219_)
  );
  AND2_X1 _46818_ (
    .A1(_12217_),
    .A2(_12219_),
    .ZN(_12220_)
  );
  INV_X1 _46819_ (
    .A(_12220_),
    .ZN(_00452_)
  );
  AND2_X1 _46820_ (
    .A1(reg_op2[3]),
    .A2(_12203_),
    .ZN(mem_la_wdata[3])
  );
  AND2_X1 _46821_ (
    .A1(mem_wdata[3]),
    .A2(_12205_),
    .ZN(_12221_)
  );
  INV_X1 _46822_ (
    .A(_12221_),
    .ZN(_12222_)
  );
  AND2_X1 _46823_ (
    .A1(_12204_),
    .A2(mem_la_wdata[3]),
    .ZN(_12223_)
  );
  INV_X1 _46824_ (
    .A(_12223_),
    .ZN(_12224_)
  );
  AND2_X1 _46825_ (
    .A1(_12222_),
    .A2(_12224_),
    .ZN(_12225_)
  );
  INV_X1 _46826_ (
    .A(_12225_),
    .ZN(_00453_)
  );
  AND2_X1 _46827_ (
    .A1(reg_op2[4]),
    .A2(_12203_),
    .ZN(mem_la_wdata[4])
  );
  AND2_X1 _46828_ (
    .A1(mem_wdata[4]),
    .A2(_12205_),
    .ZN(_12226_)
  );
  INV_X1 _46829_ (
    .A(_12226_),
    .ZN(_12227_)
  );
  AND2_X1 _46830_ (
    .A1(_12204_),
    .A2(mem_la_wdata[4]),
    .ZN(_12228_)
  );
  INV_X1 _46831_ (
    .A(_12228_),
    .ZN(_12229_)
  );
  AND2_X1 _46832_ (
    .A1(_12227_),
    .A2(_12229_),
    .ZN(_12230_)
  );
  INV_X1 _46833_ (
    .A(_12230_),
    .ZN(_00454_)
  );
  AND2_X1 _46834_ (
    .A1(reg_op2[5]),
    .A2(_12203_),
    .ZN(mem_la_wdata[5])
  );
  AND2_X1 _46835_ (
    .A1(_12204_),
    .A2(mem_la_wdata[5]),
    .ZN(_12231_)
  );
  INV_X1 _46836_ (
    .A(_12231_),
    .ZN(_12232_)
  );
  AND2_X1 _46837_ (
    .A1(mem_wdata[5]),
    .A2(_12205_),
    .ZN(_12233_)
  );
  INV_X1 _46838_ (
    .A(_12233_),
    .ZN(_12234_)
  );
  AND2_X1 _46839_ (
    .A1(_12232_),
    .A2(_12234_),
    .ZN(_12235_)
  );
  INV_X1 _46840_ (
    .A(_12235_),
    .ZN(_00455_)
  );
  AND2_X1 _46841_ (
    .A1(reg_op2[6]),
    .A2(_12203_),
    .ZN(mem_la_wdata[6])
  );
  AND2_X1 _46842_ (
    .A1(mem_wdata[6]),
    .A2(_12205_),
    .ZN(_12236_)
  );
  INV_X1 _46843_ (
    .A(_12236_),
    .ZN(_12237_)
  );
  AND2_X1 _46844_ (
    .A1(_12204_),
    .A2(mem_la_wdata[6]),
    .ZN(_12238_)
  );
  INV_X1 _46845_ (
    .A(_12238_),
    .ZN(_12239_)
  );
  AND2_X1 _46846_ (
    .A1(_12237_),
    .A2(_12239_),
    .ZN(_12240_)
  );
  INV_X1 _46847_ (
    .A(_12240_),
    .ZN(_00456_)
  );
  AND2_X1 _46848_ (
    .A1(reg_op2[7]),
    .A2(_12203_),
    .ZN(mem_la_wdata[7])
  );
  AND2_X1 _46849_ (
    .A1(mem_wdata[7]),
    .A2(_12205_),
    .ZN(_12241_)
  );
  INV_X1 _46850_ (
    .A(_12241_),
    .ZN(_12242_)
  );
  AND2_X1 _46851_ (
    .A1(_12204_),
    .A2(mem_la_wdata[7]),
    .ZN(_12243_)
  );
  INV_X1 _46852_ (
    .A(_12243_),
    .ZN(_12244_)
  );
  AND2_X1 _46853_ (
    .A1(_12242_),
    .A2(_12244_),
    .ZN(_12245_)
  );
  INV_X1 _46854_ (
    .A(_12245_),
    .ZN(_00457_)
  );
  AND2_X1 _46855_ (
    .A1(reg_op2[0]),
    .A2(_12196_),
    .ZN(_12246_)
  );
  INV_X1 _46856_ (
    .A(_12246_),
    .ZN(_12247_)
  );
  AND2_X1 _46857_ (
    .A1(reg_op2[8]),
    .A2(_12198_),
    .ZN(_12248_)
  );
  INV_X1 _46858_ (
    .A(_12248_),
    .ZN(_12249_)
  );
  AND2_X1 _46859_ (
    .A1(_12247_),
    .A2(_12249_),
    .ZN(_12250_)
  );
  AND2_X1 _46860_ (
    .A1(reg_op2[8]),
    .A2(_12194_),
    .ZN(_12251_)
  );
  INV_X1 _46861_ (
    .A(_12251_),
    .ZN(_12252_)
  );
  AND2_X1 _46862_ (
    .A1(_12250_),
    .A2(_12252_),
    .ZN(_12253_)
  );
  INV_X1 _46863_ (
    .A(_12253_),
    .ZN(mem_la_wdata[8])
  );
  AND2_X1 _46864_ (
    .A1(_12204_),
    .A2(_12253_),
    .ZN(_12254_)
  );
  INV_X1 _46865_ (
    .A(_12254_),
    .ZN(_12255_)
  );
  AND2_X1 _46866_ (
    .A1(_21324_),
    .A2(_12205_),
    .ZN(_12256_)
  );
  INV_X1 _46867_ (
    .A(_12256_),
    .ZN(_12257_)
  );
  AND2_X1 _46868_ (
    .A1(_12255_),
    .A2(_12257_),
    .ZN(_00458_)
  );
  AND2_X1 _46869_ (
    .A1(reg_op2[1]),
    .A2(_12196_),
    .ZN(_12258_)
  );
  INV_X1 _46870_ (
    .A(_12258_),
    .ZN(_12259_)
  );
  AND2_X1 _46871_ (
    .A1(reg_op2[9]),
    .A2(_12198_),
    .ZN(_12260_)
  );
  INV_X1 _46872_ (
    .A(_12260_),
    .ZN(_12261_)
  );
  AND2_X1 _46873_ (
    .A1(_12259_),
    .A2(_12261_),
    .ZN(_12262_)
  );
  AND2_X1 _46874_ (
    .A1(reg_op2[9]),
    .A2(_12194_),
    .ZN(_12263_)
  );
  INV_X1 _46875_ (
    .A(_12263_),
    .ZN(_12264_)
  );
  AND2_X1 _46876_ (
    .A1(_12262_),
    .A2(_12264_),
    .ZN(_12265_)
  );
  INV_X1 _46877_ (
    .A(_12265_),
    .ZN(mem_la_wdata[9])
  );
  AND2_X1 _46878_ (
    .A1(_12204_),
    .A2(_12265_),
    .ZN(_12266_)
  );
  INV_X1 _46879_ (
    .A(_12266_),
    .ZN(_12267_)
  );
  AND2_X1 _46880_ (
    .A1(_21325_),
    .A2(_12205_),
    .ZN(_12268_)
  );
  INV_X1 _46881_ (
    .A(_12268_),
    .ZN(_12269_)
  );
  AND2_X1 _46882_ (
    .A1(_12267_),
    .A2(_12269_),
    .ZN(_00459_)
  );
  AND2_X1 _46883_ (
    .A1(reg_op2[2]),
    .A2(_12196_),
    .ZN(_12270_)
  );
  INV_X1 _46884_ (
    .A(_12270_),
    .ZN(_12271_)
  );
  AND2_X1 _46885_ (
    .A1(reg_op2[10]),
    .A2(_12198_),
    .ZN(_12272_)
  );
  INV_X1 _46886_ (
    .A(_12272_),
    .ZN(_12273_)
  );
  AND2_X1 _46887_ (
    .A1(_12271_),
    .A2(_12273_),
    .ZN(_12274_)
  );
  AND2_X1 _46888_ (
    .A1(reg_op2[10]),
    .A2(_12194_),
    .ZN(_12275_)
  );
  INV_X1 _46889_ (
    .A(_12275_),
    .ZN(_12276_)
  );
  AND2_X1 _46890_ (
    .A1(_12274_),
    .A2(_12276_),
    .ZN(_12277_)
  );
  INV_X1 _46891_ (
    .A(_12277_),
    .ZN(mem_la_wdata[10])
  );
  AND2_X1 _46892_ (
    .A1(_12204_),
    .A2(_12277_),
    .ZN(_12278_)
  );
  INV_X1 _46893_ (
    .A(_12278_),
    .ZN(_12279_)
  );
  AND2_X1 _46894_ (
    .A1(_21326_),
    .A2(_12205_),
    .ZN(_12280_)
  );
  INV_X1 _46895_ (
    .A(_12280_),
    .ZN(_12281_)
  );
  AND2_X1 _46896_ (
    .A1(_12279_),
    .A2(_12281_),
    .ZN(_00460_)
  );
  AND2_X1 _46897_ (
    .A1(reg_op2[3]),
    .A2(_12196_),
    .ZN(_12282_)
  );
  INV_X1 _46898_ (
    .A(_12282_),
    .ZN(_12283_)
  );
  AND2_X1 _46899_ (
    .A1(reg_op2[11]),
    .A2(_12198_),
    .ZN(_12284_)
  );
  INV_X1 _46900_ (
    .A(_12284_),
    .ZN(_12285_)
  );
  AND2_X1 _46901_ (
    .A1(_12283_),
    .A2(_12285_),
    .ZN(_12286_)
  );
  AND2_X1 _46902_ (
    .A1(reg_op2[11]),
    .A2(_12194_),
    .ZN(_12287_)
  );
  INV_X1 _46903_ (
    .A(_12287_),
    .ZN(_12288_)
  );
  AND2_X1 _46904_ (
    .A1(_12286_),
    .A2(_12288_),
    .ZN(_12289_)
  );
  INV_X1 _46905_ (
    .A(_12289_),
    .ZN(mem_la_wdata[11])
  );
  AND2_X1 _46906_ (
    .A1(_12204_),
    .A2(_12289_),
    .ZN(_12290_)
  );
  INV_X1 _46907_ (
    .A(_12290_),
    .ZN(_12291_)
  );
  AND2_X1 _46908_ (
    .A1(_21327_),
    .A2(_12205_),
    .ZN(_12292_)
  );
  INV_X1 _46909_ (
    .A(_12292_),
    .ZN(_12293_)
  );
  AND2_X1 _46910_ (
    .A1(_12291_),
    .A2(_12293_),
    .ZN(_00461_)
  );
  AND2_X1 _46911_ (
    .A1(reg_op2[4]),
    .A2(_12196_),
    .ZN(_12294_)
  );
  INV_X1 _46912_ (
    .A(_12294_),
    .ZN(_12295_)
  );
  AND2_X1 _46913_ (
    .A1(reg_op2[12]),
    .A2(_12198_),
    .ZN(_12296_)
  );
  INV_X1 _46914_ (
    .A(_12296_),
    .ZN(_12297_)
  );
  AND2_X1 _46915_ (
    .A1(_12295_),
    .A2(_12297_),
    .ZN(_12298_)
  );
  AND2_X1 _46916_ (
    .A1(reg_op2[12]),
    .A2(_12194_),
    .ZN(_12299_)
  );
  INV_X1 _46917_ (
    .A(_12299_),
    .ZN(_12300_)
  );
  AND2_X1 _46918_ (
    .A1(_12298_),
    .A2(_12300_),
    .ZN(_12301_)
  );
  INV_X1 _46919_ (
    .A(_12301_),
    .ZN(mem_la_wdata[12])
  );
  AND2_X1 _46920_ (
    .A1(_12204_),
    .A2(_12301_),
    .ZN(_12302_)
  );
  INV_X1 _46921_ (
    .A(_12302_),
    .ZN(_12303_)
  );
  AND2_X1 _46922_ (
    .A1(_21328_),
    .A2(_12205_),
    .ZN(_12304_)
  );
  INV_X1 _46923_ (
    .A(_12304_),
    .ZN(_12305_)
  );
  AND2_X1 _46924_ (
    .A1(_12303_),
    .A2(_12305_),
    .ZN(_00462_)
  );
  AND2_X1 _46925_ (
    .A1(reg_op2[5]),
    .A2(_12196_),
    .ZN(_12306_)
  );
  INV_X1 _46926_ (
    .A(_12306_),
    .ZN(_12307_)
  );
  AND2_X1 _46927_ (
    .A1(reg_op2[13]),
    .A2(_12198_),
    .ZN(_12308_)
  );
  INV_X1 _46928_ (
    .A(_12308_),
    .ZN(_12309_)
  );
  AND2_X1 _46929_ (
    .A1(_12307_),
    .A2(_12309_),
    .ZN(_12310_)
  );
  AND2_X1 _46930_ (
    .A1(reg_op2[13]),
    .A2(_12194_),
    .ZN(_12311_)
  );
  INV_X1 _46931_ (
    .A(_12311_),
    .ZN(_12312_)
  );
  AND2_X1 _46932_ (
    .A1(_12310_),
    .A2(_12312_),
    .ZN(_12313_)
  );
  INV_X1 _46933_ (
    .A(_12313_),
    .ZN(mem_la_wdata[13])
  );
  AND2_X1 _46934_ (
    .A1(_12204_),
    .A2(_12313_),
    .ZN(_12314_)
  );
  INV_X1 _46935_ (
    .A(_12314_),
    .ZN(_12315_)
  );
  AND2_X1 _46936_ (
    .A1(_21329_),
    .A2(_12205_),
    .ZN(_12316_)
  );
  INV_X1 _46937_ (
    .A(_12316_),
    .ZN(_12317_)
  );
  AND2_X1 _46938_ (
    .A1(_12315_),
    .A2(_12317_),
    .ZN(_00463_)
  );
  AND2_X1 _46939_ (
    .A1(reg_op2[6]),
    .A2(_12196_),
    .ZN(_12318_)
  );
  INV_X1 _46940_ (
    .A(_12318_),
    .ZN(_12319_)
  );
  AND2_X1 _46941_ (
    .A1(reg_op2[14]),
    .A2(_12198_),
    .ZN(_12320_)
  );
  INV_X1 _46942_ (
    .A(_12320_),
    .ZN(_12321_)
  );
  AND2_X1 _46943_ (
    .A1(_12319_),
    .A2(_12321_),
    .ZN(_12322_)
  );
  AND2_X1 _46944_ (
    .A1(reg_op2[14]),
    .A2(_12194_),
    .ZN(_12323_)
  );
  INV_X1 _46945_ (
    .A(_12323_),
    .ZN(_12324_)
  );
  AND2_X1 _46946_ (
    .A1(_12322_),
    .A2(_12324_),
    .ZN(_12325_)
  );
  INV_X1 _46947_ (
    .A(_12325_),
    .ZN(mem_la_wdata[14])
  );
  AND2_X1 _46948_ (
    .A1(_12204_),
    .A2(_12325_),
    .ZN(_12326_)
  );
  INV_X1 _46949_ (
    .A(_12326_),
    .ZN(_12327_)
  );
  AND2_X1 _46950_ (
    .A1(_21330_),
    .A2(_12205_),
    .ZN(_12328_)
  );
  INV_X1 _46951_ (
    .A(_12328_),
    .ZN(_12329_)
  );
  AND2_X1 _46952_ (
    .A1(_12327_),
    .A2(_12329_),
    .ZN(_00464_)
  );
  AND2_X1 _46953_ (
    .A1(reg_op2[7]),
    .A2(_12196_),
    .ZN(_12330_)
  );
  INV_X1 _46954_ (
    .A(_12330_),
    .ZN(_12331_)
  );
  AND2_X1 _46955_ (
    .A1(reg_op2[15]),
    .A2(_12198_),
    .ZN(_12332_)
  );
  INV_X1 _46956_ (
    .A(_12332_),
    .ZN(_12333_)
  );
  AND2_X1 _46957_ (
    .A1(_12331_),
    .A2(_12333_),
    .ZN(_12334_)
  );
  AND2_X1 _46958_ (
    .A1(reg_op2[15]),
    .A2(_12194_),
    .ZN(_12335_)
  );
  INV_X1 _46959_ (
    .A(_12335_),
    .ZN(_12336_)
  );
  AND2_X1 _46960_ (
    .A1(_12334_),
    .A2(_12336_),
    .ZN(_12337_)
  );
  INV_X1 _46961_ (
    .A(_12337_),
    .ZN(mem_la_wdata[15])
  );
  AND2_X1 _46962_ (
    .A1(_12204_),
    .A2(_12337_),
    .ZN(_12338_)
  );
  INV_X1 _46963_ (
    .A(_12338_),
    .ZN(_12339_)
  );
  AND2_X1 _46964_ (
    .A1(_21331_),
    .A2(_12205_),
    .ZN(_12340_)
  );
  INV_X1 _46965_ (
    .A(_12340_),
    .ZN(_12341_)
  );
  AND2_X1 _46966_ (
    .A1(_12339_),
    .A2(_12341_),
    .ZN(_00465_)
  );
  AND2_X1 _46967_ (
    .A1(reg_op2[16]),
    .A2(_12194_),
    .ZN(_12342_)
  );
  INV_X1 _46968_ (
    .A(_12342_),
    .ZN(_12343_)
  );
  AND2_X1 _46969_ (
    .A1(reg_op2[0]),
    .A2(_12201_),
    .ZN(_12344_)
  );
  INV_X1 _46970_ (
    .A(_12344_),
    .ZN(_12345_)
  );
  AND2_X1 _46971_ (
    .A1(_12343_),
    .A2(_12345_),
    .ZN(_12346_)
  );
  INV_X1 _46972_ (
    .A(_12346_),
    .ZN(mem_la_wdata[16])
  );
  AND2_X1 _46973_ (
    .A1(_12204_),
    .A2(_12346_),
    .ZN(_12347_)
  );
  INV_X1 _46974_ (
    .A(_12347_),
    .ZN(_12348_)
  );
  AND2_X1 _46975_ (
    .A1(_21332_),
    .A2(_12205_),
    .ZN(_12349_)
  );
  INV_X1 _46976_ (
    .A(_12349_),
    .ZN(_12350_)
  );
  AND2_X1 _46977_ (
    .A1(_12348_),
    .A2(_12350_),
    .ZN(_00466_)
  );
  AND2_X1 _46978_ (
    .A1(reg_op2[17]),
    .A2(_12194_),
    .ZN(_12351_)
  );
  INV_X1 _46979_ (
    .A(_12351_),
    .ZN(_12352_)
  );
  AND2_X1 _46980_ (
    .A1(reg_op2[1]),
    .A2(_12201_),
    .ZN(_12353_)
  );
  INV_X1 _46981_ (
    .A(_12353_),
    .ZN(_12354_)
  );
  AND2_X1 _46982_ (
    .A1(_12352_),
    .A2(_12354_),
    .ZN(_12355_)
  );
  INV_X1 _46983_ (
    .A(_12355_),
    .ZN(mem_la_wdata[17])
  );
  AND2_X1 _46984_ (
    .A1(_12204_),
    .A2(_12355_),
    .ZN(_12356_)
  );
  INV_X1 _46985_ (
    .A(_12356_),
    .ZN(_12357_)
  );
  AND2_X1 _46986_ (
    .A1(_21333_),
    .A2(_12205_),
    .ZN(_12358_)
  );
  INV_X1 _46987_ (
    .A(_12358_),
    .ZN(_12359_)
  );
  AND2_X1 _46988_ (
    .A1(_12357_),
    .A2(_12359_),
    .ZN(_00467_)
  );
  AND2_X1 _46989_ (
    .A1(reg_op2[18]),
    .A2(_12194_),
    .ZN(_12360_)
  );
  INV_X1 _46990_ (
    .A(_12360_),
    .ZN(_12361_)
  );
  AND2_X1 _46991_ (
    .A1(reg_op2[2]),
    .A2(_12201_),
    .ZN(_12362_)
  );
  INV_X1 _46992_ (
    .A(_12362_),
    .ZN(_12363_)
  );
  AND2_X1 _46993_ (
    .A1(_12361_),
    .A2(_12363_),
    .ZN(_12364_)
  );
  INV_X1 _46994_ (
    .A(_12364_),
    .ZN(mem_la_wdata[18])
  );
  AND2_X1 _46995_ (
    .A1(_12204_),
    .A2(_12364_),
    .ZN(_12365_)
  );
  INV_X1 _46996_ (
    .A(_12365_),
    .ZN(_12366_)
  );
  AND2_X1 _46997_ (
    .A1(_21334_),
    .A2(_12205_),
    .ZN(_12367_)
  );
  INV_X1 _46998_ (
    .A(_12367_),
    .ZN(_12368_)
  );
  AND2_X1 _46999_ (
    .A1(_12366_),
    .A2(_12368_),
    .ZN(_00468_)
  );
  AND2_X1 _47000_ (
    .A1(reg_op2[19]),
    .A2(_12194_),
    .ZN(_12369_)
  );
  INV_X1 _47001_ (
    .A(_12369_),
    .ZN(_12370_)
  );
  AND2_X1 _47002_ (
    .A1(reg_op2[3]),
    .A2(_12201_),
    .ZN(_12371_)
  );
  INV_X1 _47003_ (
    .A(_12371_),
    .ZN(_12372_)
  );
  AND2_X1 _47004_ (
    .A1(_12370_),
    .A2(_12372_),
    .ZN(_12373_)
  );
  INV_X1 _47005_ (
    .A(_12373_),
    .ZN(mem_la_wdata[19])
  );
  AND2_X1 _47006_ (
    .A1(_12204_),
    .A2(_12373_),
    .ZN(_12374_)
  );
  INV_X1 _47007_ (
    .A(_12374_),
    .ZN(_12375_)
  );
  AND2_X1 _47008_ (
    .A1(_21335_),
    .A2(_12205_),
    .ZN(_12376_)
  );
  INV_X1 _47009_ (
    .A(_12376_),
    .ZN(_12377_)
  );
  AND2_X1 _47010_ (
    .A1(_12375_),
    .A2(_12377_),
    .ZN(_00469_)
  );
  AND2_X1 _47011_ (
    .A1(reg_op2[20]),
    .A2(_12194_),
    .ZN(_12378_)
  );
  INV_X1 _47012_ (
    .A(_12378_),
    .ZN(_12379_)
  );
  AND2_X1 _47013_ (
    .A1(reg_op2[4]),
    .A2(_12201_),
    .ZN(_12380_)
  );
  INV_X1 _47014_ (
    .A(_12380_),
    .ZN(_12381_)
  );
  AND2_X1 _47015_ (
    .A1(_12379_),
    .A2(_12381_),
    .ZN(_12382_)
  );
  INV_X1 _47016_ (
    .A(_12382_),
    .ZN(mem_la_wdata[20])
  );
  AND2_X1 _47017_ (
    .A1(_12204_),
    .A2(_12382_),
    .ZN(_12383_)
  );
  INV_X1 _47018_ (
    .A(_12383_),
    .ZN(_12384_)
  );
  AND2_X1 _47019_ (
    .A1(_21336_),
    .A2(_12205_),
    .ZN(_12385_)
  );
  INV_X1 _47020_ (
    .A(_12385_),
    .ZN(_12386_)
  );
  AND2_X1 _47021_ (
    .A1(_12384_),
    .A2(_12386_),
    .ZN(_00470_)
  );
  AND2_X1 _47022_ (
    .A1(reg_op2[21]),
    .A2(_12194_),
    .ZN(_12387_)
  );
  INV_X1 _47023_ (
    .A(_12387_),
    .ZN(_12388_)
  );
  AND2_X1 _47024_ (
    .A1(reg_op2[5]),
    .A2(_12201_),
    .ZN(_12389_)
  );
  INV_X1 _47025_ (
    .A(_12389_),
    .ZN(_12390_)
  );
  AND2_X1 _47026_ (
    .A1(_12388_),
    .A2(_12390_),
    .ZN(_12391_)
  );
  INV_X1 _47027_ (
    .A(_12391_),
    .ZN(mem_la_wdata[21])
  );
  AND2_X1 _47028_ (
    .A1(_12204_),
    .A2(_12391_),
    .ZN(_12392_)
  );
  INV_X1 _47029_ (
    .A(_12392_),
    .ZN(_12393_)
  );
  AND2_X1 _47030_ (
    .A1(_21337_),
    .A2(_12205_),
    .ZN(_12394_)
  );
  INV_X1 _47031_ (
    .A(_12394_),
    .ZN(_12395_)
  );
  AND2_X1 _47032_ (
    .A1(_12393_),
    .A2(_12395_),
    .ZN(_00471_)
  );
  AND2_X1 _47033_ (
    .A1(reg_op2[22]),
    .A2(_12194_),
    .ZN(_12396_)
  );
  INV_X1 _47034_ (
    .A(_12396_),
    .ZN(_12397_)
  );
  AND2_X1 _47035_ (
    .A1(reg_op2[6]),
    .A2(_12201_),
    .ZN(_12398_)
  );
  INV_X1 _47036_ (
    .A(_12398_),
    .ZN(_12399_)
  );
  AND2_X1 _47037_ (
    .A1(_12397_),
    .A2(_12399_),
    .ZN(_12400_)
  );
  INV_X1 _47038_ (
    .A(_12400_),
    .ZN(mem_la_wdata[22])
  );
  AND2_X1 _47039_ (
    .A1(_12204_),
    .A2(_12400_),
    .ZN(_12401_)
  );
  INV_X1 _47040_ (
    .A(_12401_),
    .ZN(_12402_)
  );
  AND2_X1 _47041_ (
    .A1(_21338_),
    .A2(_12205_),
    .ZN(_12403_)
  );
  INV_X1 _47042_ (
    .A(_12403_),
    .ZN(_12404_)
  );
  AND2_X1 _47043_ (
    .A1(_12402_),
    .A2(_12404_),
    .ZN(_00472_)
  );
  AND2_X1 _47044_ (
    .A1(reg_op2[23]),
    .A2(_12194_),
    .ZN(_12405_)
  );
  INV_X1 _47045_ (
    .A(_12405_),
    .ZN(_12406_)
  );
  AND2_X1 _47046_ (
    .A1(reg_op2[7]),
    .A2(_12201_),
    .ZN(_12407_)
  );
  INV_X1 _47047_ (
    .A(_12407_),
    .ZN(_12408_)
  );
  AND2_X1 _47048_ (
    .A1(_12406_),
    .A2(_12408_),
    .ZN(_12409_)
  );
  INV_X1 _47049_ (
    .A(_12409_),
    .ZN(mem_la_wdata[23])
  );
  AND2_X1 _47050_ (
    .A1(_12204_),
    .A2(_12409_),
    .ZN(_12410_)
  );
  INV_X1 _47051_ (
    .A(_12410_),
    .ZN(_12411_)
  );
  AND2_X1 _47052_ (
    .A1(_21339_),
    .A2(_12205_),
    .ZN(_12412_)
  );
  INV_X1 _47053_ (
    .A(_12412_),
    .ZN(_12413_)
  );
  AND2_X1 _47054_ (
    .A1(_12411_),
    .A2(_12413_),
    .ZN(_00473_)
  );
  AND2_X1 _47055_ (
    .A1(reg_op2[24]),
    .A2(_12194_),
    .ZN(_12414_)
  );
  INV_X1 _47056_ (
    .A(_12414_),
    .ZN(_12415_)
  );
  AND2_X1 _47057_ (
    .A1(_12250_),
    .A2(_12415_),
    .ZN(_12416_)
  );
  INV_X1 _47058_ (
    .A(_12416_),
    .ZN(mem_la_wdata[24])
  );
  AND2_X1 _47059_ (
    .A1(_12204_),
    .A2(_12416_),
    .ZN(_12417_)
  );
  INV_X1 _47060_ (
    .A(_12417_),
    .ZN(_12418_)
  );
  AND2_X1 _47061_ (
    .A1(_21340_),
    .A2(_12205_),
    .ZN(_12419_)
  );
  INV_X1 _47062_ (
    .A(_12419_),
    .ZN(_12420_)
  );
  AND2_X1 _47063_ (
    .A1(_12418_),
    .A2(_12420_),
    .ZN(_00474_)
  );
  AND2_X1 _47064_ (
    .A1(reg_op2[25]),
    .A2(_12194_),
    .ZN(_12421_)
  );
  INV_X1 _47065_ (
    .A(_12421_),
    .ZN(_12422_)
  );
  AND2_X1 _47066_ (
    .A1(_12262_),
    .A2(_12422_),
    .ZN(_12423_)
  );
  INV_X1 _47067_ (
    .A(_12423_),
    .ZN(mem_la_wdata[25])
  );
  AND2_X1 _47068_ (
    .A1(_12204_),
    .A2(_12423_),
    .ZN(_12424_)
  );
  INV_X1 _47069_ (
    .A(_12424_),
    .ZN(_12425_)
  );
  AND2_X1 _47070_ (
    .A1(_21341_),
    .A2(_12205_),
    .ZN(_12426_)
  );
  INV_X1 _47071_ (
    .A(_12426_),
    .ZN(_12427_)
  );
  AND2_X1 _47072_ (
    .A1(_12425_),
    .A2(_12427_),
    .ZN(_00475_)
  );
  AND2_X1 _47073_ (
    .A1(reg_op2[26]),
    .A2(_12194_),
    .ZN(_12428_)
  );
  INV_X1 _47074_ (
    .A(_12428_),
    .ZN(_12429_)
  );
  AND2_X1 _47075_ (
    .A1(_12274_),
    .A2(_12429_),
    .ZN(_12430_)
  );
  INV_X1 _47076_ (
    .A(_12430_),
    .ZN(mem_la_wdata[26])
  );
  AND2_X1 _47077_ (
    .A1(_12204_),
    .A2(_12430_),
    .ZN(_12431_)
  );
  INV_X1 _47078_ (
    .A(_12431_),
    .ZN(_12432_)
  );
  AND2_X1 _47079_ (
    .A1(_21342_),
    .A2(_12205_),
    .ZN(_12433_)
  );
  INV_X1 _47080_ (
    .A(_12433_),
    .ZN(_12434_)
  );
  AND2_X1 _47081_ (
    .A1(_12432_),
    .A2(_12434_),
    .ZN(_00476_)
  );
  AND2_X1 _47082_ (
    .A1(reg_op2[27]),
    .A2(_12194_),
    .ZN(_12435_)
  );
  INV_X1 _47083_ (
    .A(_12435_),
    .ZN(_12436_)
  );
  AND2_X1 _47084_ (
    .A1(_12286_),
    .A2(_12436_),
    .ZN(_12437_)
  );
  INV_X1 _47085_ (
    .A(_12437_),
    .ZN(mem_la_wdata[27])
  );
  AND2_X1 _47086_ (
    .A1(_12204_),
    .A2(_12437_),
    .ZN(_12438_)
  );
  INV_X1 _47087_ (
    .A(_12438_),
    .ZN(_12439_)
  );
  AND2_X1 _47088_ (
    .A1(_21343_),
    .A2(_12205_),
    .ZN(_12440_)
  );
  INV_X1 _47089_ (
    .A(_12440_),
    .ZN(_12441_)
  );
  AND2_X1 _47090_ (
    .A1(_12439_),
    .A2(_12441_),
    .ZN(_00477_)
  );
  AND2_X1 _47091_ (
    .A1(reg_op2[28]),
    .A2(_12194_),
    .ZN(_12442_)
  );
  INV_X1 _47092_ (
    .A(_12442_),
    .ZN(_12443_)
  );
  AND2_X1 _47093_ (
    .A1(_12298_),
    .A2(_12443_),
    .ZN(_12444_)
  );
  INV_X1 _47094_ (
    .A(_12444_),
    .ZN(mem_la_wdata[28])
  );
  AND2_X1 _47095_ (
    .A1(_12204_),
    .A2(_12444_),
    .ZN(_12445_)
  );
  INV_X1 _47096_ (
    .A(_12445_),
    .ZN(_12446_)
  );
  AND2_X1 _47097_ (
    .A1(_21344_),
    .A2(_12205_),
    .ZN(_12447_)
  );
  INV_X1 _47098_ (
    .A(_12447_),
    .ZN(_12448_)
  );
  AND2_X1 _47099_ (
    .A1(_12446_),
    .A2(_12448_),
    .ZN(_00478_)
  );
  AND2_X1 _47100_ (
    .A1(reg_op2[29]),
    .A2(_12194_),
    .ZN(_12449_)
  );
  INV_X1 _47101_ (
    .A(_12449_),
    .ZN(_12450_)
  );
  AND2_X1 _47102_ (
    .A1(_12310_),
    .A2(_12450_),
    .ZN(_12451_)
  );
  INV_X1 _47103_ (
    .A(_12451_),
    .ZN(mem_la_wdata[29])
  );
  AND2_X1 _47104_ (
    .A1(_12204_),
    .A2(_12451_),
    .ZN(_12452_)
  );
  INV_X1 _47105_ (
    .A(_12452_),
    .ZN(_12453_)
  );
  AND2_X1 _47106_ (
    .A1(_21345_),
    .A2(_12205_),
    .ZN(_12454_)
  );
  INV_X1 _47107_ (
    .A(_12454_),
    .ZN(_12455_)
  );
  AND2_X1 _47108_ (
    .A1(_12453_),
    .A2(_12455_),
    .ZN(_00479_)
  );
  AND2_X1 _47109_ (
    .A1(reg_op2[30]),
    .A2(_12194_),
    .ZN(_12456_)
  );
  INV_X1 _47110_ (
    .A(_12456_),
    .ZN(_12457_)
  );
  AND2_X1 _47111_ (
    .A1(_12322_),
    .A2(_12457_),
    .ZN(_12458_)
  );
  INV_X1 _47112_ (
    .A(_12458_),
    .ZN(mem_la_wdata[30])
  );
  AND2_X1 _47113_ (
    .A1(_12204_),
    .A2(_12458_),
    .ZN(_12459_)
  );
  INV_X1 _47114_ (
    .A(_12459_),
    .ZN(_12460_)
  );
  AND2_X1 _47115_ (
    .A1(_21346_),
    .A2(_12205_),
    .ZN(_12461_)
  );
  INV_X1 _47116_ (
    .A(_12461_),
    .ZN(_12462_)
  );
  AND2_X1 _47117_ (
    .A1(_12460_),
    .A2(_12462_),
    .ZN(_00480_)
  );
  AND2_X1 _47118_ (
    .A1(reg_op2[31]),
    .A2(_12194_),
    .ZN(_12463_)
  );
  INV_X1 _47119_ (
    .A(_12463_),
    .ZN(_12464_)
  );
  AND2_X1 _47120_ (
    .A1(_12334_),
    .A2(_12464_),
    .ZN(_12465_)
  );
  INV_X1 _47121_ (
    .A(_12465_),
    .ZN(mem_la_wdata[31])
  );
  AND2_X1 _47122_ (
    .A1(_12204_),
    .A2(_12465_),
    .ZN(_12466_)
  );
  INV_X1 _47123_ (
    .A(_12466_),
    .ZN(_12467_)
  );
  AND2_X1 _47124_ (
    .A1(_21347_),
    .A2(_12205_),
    .ZN(_12468_)
  );
  INV_X1 _47125_ (
    .A(_12468_),
    .ZN(_12469_)
  );
  AND2_X1 _47126_ (
    .A1(_12467_),
    .A2(_12469_),
    .ZN(_00481_)
  );
  AND2_X1 _47127_ (
    .A1(mem_wstrb[0]),
    .A2(_11771_),
    .ZN(_12470_)
  );
  INV_X1 _47128_ (
    .A(_12470_),
    .ZN(_12471_)
  );
  AND2_X1 _47129_ (
    .A1(_29146_[1]),
    .A2(_12198_),
    .ZN(_12472_)
  );
  INV_X1 _47130_ (
    .A(_12472_),
    .ZN(_12473_)
  );
  AND2_X1 _47131_ (
    .A1(_12195_),
    .A2(_12473_),
    .ZN(_12474_)
  );
  INV_X1 _47132_ (
    .A(_12474_),
    .ZN(_12475_)
  );
  AND2_X1 _47133_ (
    .A1(_22024_),
    .A2(_12196_),
    .ZN(_12476_)
  );
  AND2_X1 _47134_ (
    .A1(_00044_),
    .A2(_12476_),
    .ZN(_12477_)
  );
  INV_X1 _47135_ (
    .A(_12477_),
    .ZN(_12478_)
  );
  AND2_X1 _47136_ (
    .A1(_12474_),
    .A2(_12478_),
    .ZN(_12479_)
  );
  INV_X1 _47137_ (
    .A(_12479_),
    .ZN(mem_la_wstrb[0])
  );
  AND2_X1 _47138_ (
    .A1(_11762_),
    .A2(_12204_),
    .ZN(_12480_)
  );
  AND2_X1 _47139_ (
    .A1(mem_la_wstrb[0]),
    .A2(_12480_),
    .ZN(_12481_)
  );
  INV_X1 _47140_ (
    .A(_12481_),
    .ZN(_12482_)
  );
  AND2_X1 _47141_ (
    .A1(mem_do_wdata),
    .A2(_11766_),
    .ZN(mem_la_write)
  );
  AND2_X1 _47142_ (
    .A1(_12471_),
    .A2(_12482_),
    .ZN(_12483_)
  );
  INV_X1 _47143_ (
    .A(_12483_),
    .ZN(_00482_)
  );
  AND2_X1 _47144_ (
    .A1(mem_wstrb[1]),
    .A2(_11771_),
    .ZN(_12484_)
  );
  INV_X1 _47145_ (
    .A(_12484_),
    .ZN(_12485_)
  );
  AND2_X1 _47146_ (
    .A1(reg_op1[0]),
    .A2(_12476_),
    .ZN(_12486_)
  );
  INV_X1 _47147_ (
    .A(_12486_),
    .ZN(_12487_)
  );
  AND2_X1 _47148_ (
    .A1(_12474_),
    .A2(_12487_),
    .ZN(_12488_)
  );
  INV_X1 _47149_ (
    .A(_12488_),
    .ZN(mem_la_wstrb[1])
  );
  AND2_X1 _47150_ (
    .A1(_12480_),
    .A2(mem_la_wstrb[1]),
    .ZN(_12489_)
  );
  INV_X1 _47151_ (
    .A(_12489_),
    .ZN(_12490_)
  );
  AND2_X1 _47152_ (
    .A1(_12485_),
    .A2(_12490_),
    .ZN(_12491_)
  );
  INV_X1 _47153_ (
    .A(_12491_),
    .ZN(_00483_)
  );
  AND2_X1 _47154_ (
    .A1(mem_wstrb[2]),
    .A2(_11771_),
    .ZN(_12492_)
  );
  INV_X1 _47155_ (
    .A(_12492_),
    .ZN(_12493_)
  );
  AND2_X1 _47156_ (
    .A1(reg_op1[1]),
    .A2(_12198_),
    .ZN(_12494_)
  );
  INV_X1 _47157_ (
    .A(_12494_),
    .ZN(_12495_)
  );
  AND2_X1 _47158_ (
    .A1(_12195_),
    .A2(_12495_),
    .ZN(_12496_)
  );
  AND2_X1 _47159_ (
    .A1(reg_op1[1]),
    .A2(_12196_),
    .ZN(_12497_)
  );
  AND2_X1 _47160_ (
    .A1(_00044_),
    .A2(_12497_),
    .ZN(_12498_)
  );
  INV_X1 _47161_ (
    .A(_12498_),
    .ZN(_12499_)
  );
  AND2_X1 _47162_ (
    .A1(_12496_),
    .A2(_12499_),
    .ZN(_12500_)
  );
  INV_X1 _47163_ (
    .A(_12500_),
    .ZN(mem_la_wstrb[2])
  );
  AND2_X1 _47164_ (
    .A1(_12480_),
    .A2(mem_la_wstrb[2]),
    .ZN(_12501_)
  );
  INV_X1 _47165_ (
    .A(_12501_),
    .ZN(_12502_)
  );
  AND2_X1 _47166_ (
    .A1(_12493_),
    .A2(_12502_),
    .ZN(_12503_)
  );
  INV_X1 _47167_ (
    .A(_12503_),
    .ZN(_00484_)
  );
  AND2_X1 _47168_ (
    .A1(mem_wstrb[3]),
    .A2(_11771_),
    .ZN(_12504_)
  );
  INV_X1 _47169_ (
    .A(_12504_),
    .ZN(_12505_)
  );
  AND2_X1 _47170_ (
    .A1(reg_op1[0]),
    .A2(_12497_),
    .ZN(_12506_)
  );
  INV_X1 _47171_ (
    .A(_12506_),
    .ZN(_12507_)
  );
  AND2_X1 _47172_ (
    .A1(_12496_),
    .A2(_12507_),
    .ZN(_12508_)
  );
  INV_X1 _47173_ (
    .A(_12508_),
    .ZN(mem_la_wstrb[3])
  );
  AND2_X1 _47174_ (
    .A1(_12480_),
    .A2(mem_la_wstrb[3]),
    .ZN(_12509_)
  );
  INV_X1 _47175_ (
    .A(_12509_),
    .ZN(_12510_)
  );
  AND2_X1 _47176_ (
    .A1(_12505_),
    .A2(_12510_),
    .ZN(_12511_)
  );
  INV_X1 _47177_ (
    .A(_12511_),
    .ZN(_00485_)
  );
  AND2_X1 _47178_ (
    .A1(_22061_),
    .A2(_22062_),
    .ZN(_12512_)
  );
  INV_X1 _47179_ (
    .A(_12512_),
    .ZN(_12513_)
  );
  AND2_X1 _47180_ (
    .A1(_21070_),
    .A2(_12512_),
    .ZN(_12514_)
  );
  INV_X1 _47181_ (
    .A(_12514_),
    .ZN(_12515_)
  );
  AND2_X1 _47182_ (
    .A1(_22076_),
    .A2(_12515_),
    .ZN(_12516_)
  );
  AND2_X1 _47183_ (
    .A1(_11796_),
    .A2(_12516_),
    .ZN(_12517_)
  );
  INV_X1 _47184_ (
    .A(_12517_),
    .ZN(_12518_)
  );
  AND2_X1 _47185_ (
    .A1(resetn),
    .A2(_12518_),
    .ZN(_12519_)
  );
  INV_X1 _47186_ (
    .A(_12519_),
    .ZN(_12520_)
  );
  AND2_X1 _47187_ (
    .A1(_11791_),
    .A2(_12513_),
    .ZN(_12521_)
  );
  INV_X1 _47188_ (
    .A(_12521_),
    .ZN(_12522_)
  );
  AND2_X1 _47189_ (
    .A1(_11780_),
    .A2(_12522_),
    .ZN(_12523_)
  );
  AND2_X1 _47190_ (
    .A1(_12520_),
    .A2(_12523_),
    .ZN(_12524_)
  );
  INV_X1 _47191_ (
    .A(_12524_),
    .ZN(_12525_)
  );
  AND2_X1 _47192_ (
    .A1(_22307_),
    .A2(_22310_),
    .ZN(_12526_)
  );
  AND2_X1 _47193_ (
    .A1(_11767_),
    .A2(_11786_),
    .ZN(_12527_)
  );
  AND2_X1 _47194_ (
    .A1(_12526_),
    .A2(_12527_),
    .ZN(_12528_)
  );
  INV_X1 _47195_ (
    .A(_12528_),
    .ZN(_12529_)
  );
  AND2_X1 _47196_ (
    .A1(_11769_),
    .A2(_11774_),
    .ZN(_12530_)
  );
  INV_X1 _47197_ (
    .A(_12530_),
    .ZN(_12531_)
  );
  AND2_X1 _47198_ (
    .A1(_12529_),
    .A2(_12531_),
    .ZN(_12532_)
  );
  AND2_X1 _47199_ (
    .A1(_21348_),
    .A2(_12525_),
    .ZN(_12533_)
  );
  INV_X1 _47200_ (
    .A(_12533_),
    .ZN(_12534_)
  );
  AND2_X1 _47201_ (
    .A1(_12524_),
    .A2(_12532_),
    .ZN(_12535_)
  );
  INV_X1 _47202_ (
    .A(_12535_),
    .ZN(_12536_)
  );
  AND2_X1 _47203_ (
    .A1(_12534_),
    .A2(_12536_),
    .ZN(_00486_)
  );
  AND2_X1 _47204_ (
    .A1(_12205_),
    .A2(_12529_),
    .ZN(_12537_)
  );
  AND2_X1 _47205_ (
    .A1(_21349_),
    .A2(_12525_),
    .ZN(_12538_)
  );
  INV_X1 _47206_ (
    .A(_12538_),
    .ZN(_12539_)
  );
  AND2_X1 _47207_ (
    .A1(_12524_),
    .A2(_12537_),
    .ZN(_12540_)
  );
  INV_X1 _47208_ (
    .A(_12540_),
    .ZN(_12541_)
  );
  AND2_X1 _47209_ (
    .A1(_12539_),
    .A2(_12541_),
    .ZN(_00487_)
  );
  AND2_X1 _47210_ (
    .A1(latched_store),
    .A2(_00030_),
    .ZN(_12542_)
  );
  INV_X1 _47211_ (
    .A(_12542_),
    .ZN(_12543_)
  );
  AND2_X1 _47212_ (
    .A1(_21066_),
    .A2(_12543_),
    .ZN(_12544_)
  );
  INV_X1 _47213_ (
    .A(_12544_),
    .ZN(_12545_)
  );
  AND2_X1 _47214_ (
    .A1(_02911_),
    .A2(_12545_),
    .ZN(_12546_)
  );
  AND2_X1 _47215_ (
    .A1(latched_rd[3]),
    .A2(_12546_),
    .ZN(_12547_)
  );
  INV_X1 _47216_ (
    .A(_12547_),
    .ZN(_12548_)
  );
  AND2_X1 _47217_ (
    .A1(_21254_),
    .A2(_21255_),
    .ZN(_12549_)
  );
  INV_X1 _47218_ (
    .A(_12549_),
    .ZN(_12550_)
  );
  AND2_X1 _47219_ (
    .A1(_21256_),
    .A2(_21258_),
    .ZN(_12551_)
  );
  AND2_X1 _47220_ (
    .A1(_12549_),
    .A2(_12551_),
    .ZN(_12552_)
  );
  AND2_X1 _47221_ (
    .A1(_21257_),
    .A2(_12552_),
    .ZN(_12553_)
  );
  INV_X1 _47222_ (
    .A(_12553_),
    .ZN(_12554_)
  );
  AND2_X1 _47223_ (
    .A1(_12546_),
    .A2(_12554_),
    .ZN(_12555_)
  );
  AND2_X1 _47224_ (
    .A1(latched_rd[0]),
    .A2(_12555_),
    .ZN(_12556_)
  );
  AND2_X1 _47225_ (
    .A1(_21255_),
    .A2(_12556_),
    .ZN(_12557_)
  );
  AND2_X1 _47226_ (
    .A1(_12547_),
    .A2(_12551_),
    .ZN(_12558_)
  );
  AND2_X1 _47227_ (
    .A1(_12557_),
    .A2(_12558_),
    .ZN(_12559_)
  );
  INV_X1 _47228_ (
    .A(_12559_),
    .ZN(_12560_)
  );
  AND2_X1 _47229_ (
    .A1(_03402_),
    .A2(_12542_),
    .ZN(_12561_)
  );
  INV_X1 _47230_ (
    .A(_12561_),
    .ZN(_12562_)
  );
  AND2_X1 _47231_ (
    .A1(reg_pc[3]),
    .A2(reg_pc[2]),
    .ZN(_12563_)
  );
  INV_X1 _47232_ (
    .A(_12563_),
    .ZN(_12564_)
  );
  AND2_X1 _47233_ (
    .A1(reg_pc[4]),
    .A2(_12563_),
    .ZN(_12565_)
  );
  INV_X1 _47234_ (
    .A(_12565_),
    .ZN(_12566_)
  );
  AND2_X1 _47235_ (
    .A1(reg_pc[5]),
    .A2(_12565_),
    .ZN(_12567_)
  );
  INV_X1 _47236_ (
    .A(_12567_),
    .ZN(_12568_)
  );
  AND2_X1 _47237_ (
    .A1(reg_pc[6]),
    .A2(_12567_),
    .ZN(_12569_)
  );
  INV_X1 _47238_ (
    .A(_12569_),
    .ZN(_12570_)
  );
  AND2_X1 _47239_ (
    .A1(reg_pc[7]),
    .A2(_12569_),
    .ZN(_12571_)
  );
  INV_X1 _47240_ (
    .A(_12571_),
    .ZN(_12572_)
  );
  AND2_X1 _47241_ (
    .A1(reg_pc[8]),
    .A2(_12571_),
    .ZN(_12573_)
  );
  INV_X1 _47242_ (
    .A(_12573_),
    .ZN(_12574_)
  );
  AND2_X1 _47243_ (
    .A1(reg_pc[9]),
    .A2(_12573_),
    .ZN(_12575_)
  );
  INV_X1 _47244_ (
    .A(_12575_),
    .ZN(_12576_)
  );
  AND2_X1 _47245_ (
    .A1(reg_pc[10]),
    .A2(_12575_),
    .ZN(_12577_)
  );
  INV_X1 _47246_ (
    .A(_12577_),
    .ZN(_12578_)
  );
  AND2_X1 _47247_ (
    .A1(reg_pc[11]),
    .A2(_12577_),
    .ZN(_12579_)
  );
  INV_X1 _47248_ (
    .A(_12579_),
    .ZN(_12580_)
  );
  AND2_X1 _47249_ (
    .A1(reg_pc[12]),
    .A2(_12579_),
    .ZN(_12581_)
  );
  INV_X1 _47250_ (
    .A(_12581_),
    .ZN(_12582_)
  );
  AND2_X1 _47251_ (
    .A1(reg_pc[13]),
    .A2(_12581_),
    .ZN(_12583_)
  );
  INV_X1 _47252_ (
    .A(_12583_),
    .ZN(_12584_)
  );
  AND2_X1 _47253_ (
    .A1(reg_pc[14]),
    .A2(_12583_),
    .ZN(_12585_)
  );
  INV_X1 _47254_ (
    .A(_12585_),
    .ZN(_12586_)
  );
  AND2_X1 _47255_ (
    .A1(reg_pc[15]),
    .A2(_12585_),
    .ZN(_12587_)
  );
  INV_X1 _47256_ (
    .A(_12587_),
    .ZN(_12588_)
  );
  AND2_X1 _47257_ (
    .A1(reg_pc[16]),
    .A2(_12587_),
    .ZN(_12589_)
  );
  INV_X1 _47258_ (
    .A(_12589_),
    .ZN(_12590_)
  );
  AND2_X1 _47259_ (
    .A1(reg_pc[17]),
    .A2(_12589_),
    .ZN(_12591_)
  );
  INV_X1 _47260_ (
    .A(_12591_),
    .ZN(_12592_)
  );
  AND2_X1 _47261_ (
    .A1(reg_pc[18]),
    .A2(_12591_),
    .ZN(_12593_)
  );
  INV_X1 _47262_ (
    .A(_12593_),
    .ZN(_12594_)
  );
  AND2_X1 _47263_ (
    .A1(reg_pc[19]),
    .A2(_12593_),
    .ZN(_12595_)
  );
  INV_X1 _47264_ (
    .A(_12595_),
    .ZN(_12596_)
  );
  AND2_X1 _47265_ (
    .A1(reg_pc[20]),
    .A2(_12595_),
    .ZN(_12597_)
  );
  INV_X1 _47266_ (
    .A(_12597_),
    .ZN(_12598_)
  );
  AND2_X1 _47267_ (
    .A1(reg_pc[21]),
    .A2(_12597_),
    .ZN(_12599_)
  );
  INV_X1 _47268_ (
    .A(_12599_),
    .ZN(_12600_)
  );
  AND2_X1 _47269_ (
    .A1(reg_pc[22]),
    .A2(_12599_),
    .ZN(_12601_)
  );
  INV_X1 _47270_ (
    .A(_12601_),
    .ZN(_12602_)
  );
  AND2_X1 _47271_ (
    .A1(reg_pc[23]),
    .A2(_12601_),
    .ZN(_12603_)
  );
  INV_X1 _47272_ (
    .A(_12603_),
    .ZN(_12604_)
  );
  AND2_X1 _47273_ (
    .A1(reg_pc[24]),
    .A2(_12603_),
    .ZN(_12605_)
  );
  INV_X1 _47274_ (
    .A(_12605_),
    .ZN(_12606_)
  );
  AND2_X1 _47275_ (
    .A1(reg_pc[25]),
    .A2(_12605_),
    .ZN(_12607_)
  );
  INV_X1 _47276_ (
    .A(_12607_),
    .ZN(_12608_)
  );
  AND2_X1 _47277_ (
    .A1(reg_pc[26]),
    .A2(_12607_),
    .ZN(_12609_)
  );
  INV_X1 _47278_ (
    .A(_12609_),
    .ZN(_12610_)
  );
  AND2_X1 _47279_ (
    .A1(reg_pc[27]),
    .A2(_12609_),
    .ZN(_12611_)
  );
  INV_X1 _47280_ (
    .A(_12611_),
    .ZN(_12612_)
  );
  AND2_X1 _47281_ (
    .A1(reg_pc[28]),
    .A2(_12611_),
    .ZN(_12613_)
  );
  INV_X1 _47282_ (
    .A(_12613_),
    .ZN(_12614_)
  );
  AND2_X1 _47283_ (
    .A1(reg_pc[29]),
    .A2(_12613_),
    .ZN(_12615_)
  );
  INV_X1 _47284_ (
    .A(_12615_),
    .ZN(_12616_)
  );
  AND2_X1 _47285_ (
    .A1(reg_pc[30]),
    .A2(_12615_),
    .ZN(_12617_)
  );
  INV_X1 _47286_ (
    .A(_12617_),
    .ZN(_12618_)
  );
  AND2_X1 _47287_ (
    .A1(reg_pc[31]),
    .A2(_12617_),
    .ZN(_12619_)
  );
  INV_X1 _47288_ (
    .A(_12619_),
    .ZN(_12620_)
  );
  AND2_X1 _47289_ (
    .A1(_21073_),
    .A2(_12618_),
    .ZN(_12621_)
  );
  INV_X1 _47290_ (
    .A(_12621_),
    .ZN(_12622_)
  );
  AND2_X1 _47291_ (
    .A1(latched_branch),
    .A2(_12620_),
    .ZN(_12623_)
  );
  AND2_X1 _47292_ (
    .A1(_12622_),
    .A2(_12623_),
    .ZN(_12624_)
  );
  INV_X1 _47293_ (
    .A(_12624_),
    .ZN(_12625_)
  );
  AND2_X1 _47294_ (
    .A1(_12562_),
    .A2(_12625_),
    .ZN(_12626_)
  );
  INV_X1 _47295_ (
    .A(_12626_),
    .ZN(_12627_)
  );
  AND2_X1 _47296_ (
    .A1(_12555_),
    .A2(_12627_),
    .ZN(_12628_)
  );
  AND2_X1 _47297_ (
    .A1(_12559_),
    .A2(_12628_),
    .ZN(_12629_)
  );
  INV_X1 _47298_ (
    .A(_12629_),
    .ZN(_12630_)
  );
  AND2_X1 _47299_ (
    .A1(\cpuregs[9] [31]),
    .A2(_12560_),
    .ZN(_12631_)
  );
  INV_X1 _47300_ (
    .A(_12631_),
    .ZN(_12632_)
  );
  AND2_X1 _47301_ (
    .A1(_12630_),
    .A2(_12632_),
    .ZN(_12633_)
  );
  INV_X1 _47302_ (
    .A(_12633_),
    .ZN(_00495_)
  );
  AND2_X1 _47303_ (
    .A1(_12547_),
    .A2(_12552_),
    .ZN(_12634_)
  );
  INV_X1 _47304_ (
    .A(_12634_),
    .ZN(_12635_)
  );
  AND2_X1 _47305_ (
    .A1(_12546_),
    .A2(_12550_),
    .ZN(_12636_)
  );
  INV_X1 _47306_ (
    .A(_12636_),
    .ZN(_12637_)
  );
  AND2_X1 _47307_ (
    .A1(\cpuregs[8] [31]),
    .A2(_12635_),
    .ZN(_12638_)
  );
  INV_X1 _47308_ (
    .A(_12638_),
    .ZN(_12639_)
  );
  AND2_X1 _47309_ (
    .A1(_12628_),
    .A2(_12634_),
    .ZN(_12640_)
  );
  INV_X1 _47310_ (
    .A(_12640_),
    .ZN(_12641_)
  );
  AND2_X1 _47311_ (
    .A1(_12639_),
    .A2(_12641_),
    .ZN(_12642_)
  );
  INV_X1 _47312_ (
    .A(_12642_),
    .ZN(_00496_)
  );
  AND2_X1 _47313_ (
    .A1(latched_rd[1]),
    .A2(_12556_),
    .ZN(_12643_)
  );
  AND2_X1 _47314_ (
    .A1(latched_rd[2]),
    .A2(_12546_),
    .ZN(_12644_)
  );
  INV_X1 _47315_ (
    .A(_12644_),
    .ZN(_12645_)
  );
  AND2_X1 _47316_ (
    .A1(latched_rd[4]),
    .A2(_12546_),
    .ZN(_12646_)
  );
  INV_X1 _47317_ (
    .A(_12646_),
    .ZN(_12647_)
  );
  AND2_X1 _47318_ (
    .A1(_12548_),
    .A2(_12647_),
    .ZN(_12648_)
  );
  AND2_X1 _47319_ (
    .A1(_12644_),
    .A2(_12648_),
    .ZN(_12649_)
  );
  AND2_X1 _47320_ (
    .A1(_12643_),
    .A2(_12649_),
    .ZN(_12650_)
  );
  INV_X1 _47321_ (
    .A(_12650_),
    .ZN(_12651_)
  );
  AND2_X1 _47322_ (
    .A1(_12628_),
    .A2(_12650_),
    .ZN(_12652_)
  );
  INV_X1 _47323_ (
    .A(_12652_),
    .ZN(_12653_)
  );
  AND2_X1 _47324_ (
    .A1(\cpuregs[7] [31]),
    .A2(_12651_),
    .ZN(_12654_)
  );
  INV_X1 _47325_ (
    .A(_12654_),
    .ZN(_12655_)
  );
  AND2_X1 _47326_ (
    .A1(_12653_),
    .A2(_12655_),
    .ZN(_12656_)
  );
  INV_X1 _47327_ (
    .A(_12656_),
    .ZN(_00497_)
  );
  AND2_X1 _47328_ (
    .A1(_21254_),
    .A2(latched_rd[1]),
    .ZN(_12657_)
  );
  AND2_X1 _47329_ (
    .A1(_12649_),
    .A2(_12657_),
    .ZN(_12658_)
  );
  INV_X1 _47330_ (
    .A(_12658_),
    .ZN(_12659_)
  );
  AND2_X1 _47331_ (
    .A1(_12628_),
    .A2(_12658_),
    .ZN(_12660_)
  );
  INV_X1 _47332_ (
    .A(_12660_),
    .ZN(_12661_)
  );
  AND2_X1 _47333_ (
    .A1(\cpuregs[6] [31]),
    .A2(_12659_),
    .ZN(_12662_)
  );
  INV_X1 _47334_ (
    .A(_12662_),
    .ZN(_12663_)
  );
  AND2_X1 _47335_ (
    .A1(_12661_),
    .A2(_12663_),
    .ZN(_12664_)
  );
  INV_X1 _47336_ (
    .A(_12664_),
    .ZN(_00498_)
  );
  AND2_X1 _47337_ (
    .A1(_12557_),
    .A2(_12649_),
    .ZN(_12665_)
  );
  INV_X1 _47338_ (
    .A(_12665_),
    .ZN(_12666_)
  );
  AND2_X1 _47339_ (
    .A1(_12628_),
    .A2(_12665_),
    .ZN(_12667_)
  );
  INV_X1 _47340_ (
    .A(_12667_),
    .ZN(_12668_)
  );
  AND2_X1 _47341_ (
    .A1(\cpuregs[5] [31]),
    .A2(_12666_),
    .ZN(_12669_)
  );
  INV_X1 _47342_ (
    .A(_12669_),
    .ZN(_12670_)
  );
  AND2_X1 _47343_ (
    .A1(_12668_),
    .A2(_12670_),
    .ZN(_12671_)
  );
  INV_X1 _47344_ (
    .A(_12671_),
    .ZN(_00499_)
  );
  AND2_X1 _47345_ (
    .A1(_12549_),
    .A2(_12649_),
    .ZN(_12672_)
  );
  INV_X1 _47346_ (
    .A(_12672_),
    .ZN(_12673_)
  );
  AND2_X1 _47347_ (
    .A1(_12628_),
    .A2(_12672_),
    .ZN(_12674_)
  );
  INV_X1 _47348_ (
    .A(_12674_),
    .ZN(_12675_)
  );
  AND2_X1 _47349_ (
    .A1(\cpuregs[4] [31]),
    .A2(_12673_),
    .ZN(_12676_)
  );
  INV_X1 _47350_ (
    .A(_12676_),
    .ZN(_12677_)
  );
  AND2_X1 _47351_ (
    .A1(_12675_),
    .A2(_12677_),
    .ZN(_12678_)
  );
  INV_X1 _47352_ (
    .A(_12678_),
    .ZN(_00500_)
  );
  AND2_X1 _47353_ (
    .A1(_12645_),
    .A2(_12648_),
    .ZN(_12679_)
  );
  AND2_X1 _47354_ (
    .A1(_12643_),
    .A2(_12679_),
    .ZN(_12680_)
  );
  INV_X1 _47355_ (
    .A(_12680_),
    .ZN(_12681_)
  );
  AND2_X1 _47356_ (
    .A1(_12628_),
    .A2(_12680_),
    .ZN(_12682_)
  );
  INV_X1 _47357_ (
    .A(_12682_),
    .ZN(_12683_)
  );
  AND2_X1 _47358_ (
    .A1(\cpuregs[3] [31]),
    .A2(_12681_),
    .ZN(_12684_)
  );
  INV_X1 _47359_ (
    .A(_12684_),
    .ZN(_12685_)
  );
  AND2_X1 _47360_ (
    .A1(_12683_),
    .A2(_12685_),
    .ZN(_12686_)
  );
  INV_X1 _47361_ (
    .A(_12686_),
    .ZN(_00501_)
  );
  AND2_X1 _47362_ (
    .A1(latched_rd[4]),
    .A2(_12547_),
    .ZN(_12687_)
  );
  AND2_X1 _47363_ (
    .A1(latched_rd[2]),
    .A2(_12687_),
    .ZN(_12688_)
  );
  AND2_X1 _47364_ (
    .A1(_12643_),
    .A2(_12688_),
    .ZN(_12689_)
  );
  INV_X1 _47365_ (
    .A(_12689_),
    .ZN(_12690_)
  );
  AND2_X1 _47366_ (
    .A1(_12628_),
    .A2(_12689_),
    .ZN(_12691_)
  );
  INV_X1 _47367_ (
    .A(_12691_),
    .ZN(_12692_)
  );
  AND2_X1 _47368_ (
    .A1(\cpuregs[31] [31]),
    .A2(_12690_),
    .ZN(_12693_)
  );
  INV_X1 _47369_ (
    .A(_12693_),
    .ZN(_12694_)
  );
  AND2_X1 _47370_ (
    .A1(_12692_),
    .A2(_12694_),
    .ZN(_12695_)
  );
  INV_X1 _47371_ (
    .A(_12695_),
    .ZN(_00502_)
  );
  AND2_X1 _47372_ (
    .A1(_12657_),
    .A2(_12688_),
    .ZN(_12696_)
  );
  INV_X1 _47373_ (
    .A(_12696_),
    .ZN(_12697_)
  );
  AND2_X1 _47374_ (
    .A1(_12628_),
    .A2(_12696_),
    .ZN(_12698_)
  );
  INV_X1 _47375_ (
    .A(_12698_),
    .ZN(_12699_)
  );
  AND2_X1 _47376_ (
    .A1(\cpuregs[30] [31]),
    .A2(_12697_),
    .ZN(_12700_)
  );
  INV_X1 _47377_ (
    .A(_12700_),
    .ZN(_12701_)
  );
  AND2_X1 _47378_ (
    .A1(_12699_),
    .A2(_12701_),
    .ZN(_12702_)
  );
  INV_X1 _47379_ (
    .A(_12702_),
    .ZN(_00503_)
  );
  AND2_X1 _47380_ (
    .A1(_12546_),
    .A2(_12657_),
    .ZN(_12703_)
  );
  AND2_X1 _47381_ (
    .A1(_12679_),
    .A2(_12703_),
    .ZN(_12704_)
  );
  INV_X1 _47382_ (
    .A(_12704_),
    .ZN(_12705_)
  );
  AND2_X1 _47383_ (
    .A1(_12626_),
    .A2(_12704_),
    .ZN(_12706_)
  );
  INV_X1 _47384_ (
    .A(_12706_),
    .ZN(_12707_)
  );
  AND2_X1 _47385_ (
    .A1(_21361_),
    .A2(_12705_),
    .ZN(_12708_)
  );
  INV_X1 _47386_ (
    .A(_12708_),
    .ZN(_12709_)
  );
  AND2_X1 _47387_ (
    .A1(_12707_),
    .A2(_12709_),
    .ZN(_00504_)
  );
  AND2_X1 _47388_ (
    .A1(_12557_),
    .A2(_12688_),
    .ZN(_12710_)
  );
  INV_X1 _47389_ (
    .A(_12710_),
    .ZN(_12711_)
  );
  AND2_X1 _47390_ (
    .A1(_12628_),
    .A2(_12710_),
    .ZN(_12712_)
  );
  INV_X1 _47391_ (
    .A(_12712_),
    .ZN(_12713_)
  );
  AND2_X1 _47392_ (
    .A1(\cpuregs[29] [31]),
    .A2(_12711_),
    .ZN(_12714_)
  );
  INV_X1 _47393_ (
    .A(_12714_),
    .ZN(_12715_)
  );
  AND2_X1 _47394_ (
    .A1(_12713_),
    .A2(_12715_),
    .ZN(_12716_)
  );
  INV_X1 _47395_ (
    .A(_12716_),
    .ZN(_00505_)
  );
  AND2_X1 _47396_ (
    .A1(_12549_),
    .A2(_12688_),
    .ZN(_12717_)
  );
  INV_X1 _47397_ (
    .A(_12717_),
    .ZN(_12718_)
  );
  AND2_X1 _47398_ (
    .A1(_12628_),
    .A2(_12717_),
    .ZN(_12719_)
  );
  INV_X1 _47399_ (
    .A(_12719_),
    .ZN(_12720_)
  );
  AND2_X1 _47400_ (
    .A1(\cpuregs[28] [31]),
    .A2(_12718_),
    .ZN(_12721_)
  );
  INV_X1 _47401_ (
    .A(_12721_),
    .ZN(_12722_)
  );
  AND2_X1 _47402_ (
    .A1(_12720_),
    .A2(_12722_),
    .ZN(_12723_)
  );
  INV_X1 _47403_ (
    .A(_12723_),
    .ZN(_00506_)
  );
  AND2_X1 _47404_ (
    .A1(_21256_),
    .A2(_12687_),
    .ZN(_12724_)
  );
  AND2_X1 _47405_ (
    .A1(_12643_),
    .A2(_12724_),
    .ZN(_12725_)
  );
  INV_X1 _47406_ (
    .A(_12725_),
    .ZN(_12726_)
  );
  AND2_X1 _47407_ (
    .A1(_12628_),
    .A2(_12725_),
    .ZN(_12727_)
  );
  INV_X1 _47408_ (
    .A(_12727_),
    .ZN(_12728_)
  );
  AND2_X1 _47409_ (
    .A1(\cpuregs[27] [31]),
    .A2(_12726_),
    .ZN(_12729_)
  );
  INV_X1 _47410_ (
    .A(_12729_),
    .ZN(_12730_)
  );
  AND2_X1 _47411_ (
    .A1(_12728_),
    .A2(_12730_),
    .ZN(_12731_)
  );
  INV_X1 _47412_ (
    .A(_12731_),
    .ZN(_00507_)
  );
  AND2_X1 _47413_ (
    .A1(_12703_),
    .A2(_12724_),
    .ZN(_12732_)
  );
  INV_X1 _47414_ (
    .A(_12732_),
    .ZN(_12733_)
  );
  AND2_X1 _47415_ (
    .A1(_12628_),
    .A2(_12732_),
    .ZN(_12734_)
  );
  INV_X1 _47416_ (
    .A(_12734_),
    .ZN(_12735_)
  );
  AND2_X1 _47417_ (
    .A1(\cpuregs[26] [31]),
    .A2(_12733_),
    .ZN(_12736_)
  );
  INV_X1 _47418_ (
    .A(_12736_),
    .ZN(_12737_)
  );
  AND2_X1 _47419_ (
    .A1(_12735_),
    .A2(_12737_),
    .ZN(_12738_)
  );
  INV_X1 _47420_ (
    .A(_12738_),
    .ZN(_00508_)
  );
  AND2_X1 _47421_ (
    .A1(_12557_),
    .A2(_12724_),
    .ZN(_12739_)
  );
  INV_X1 _47422_ (
    .A(_12739_),
    .ZN(_12740_)
  );
  AND2_X1 _47423_ (
    .A1(_12628_),
    .A2(_12739_),
    .ZN(_12741_)
  );
  INV_X1 _47424_ (
    .A(_12741_),
    .ZN(_12742_)
  );
  AND2_X1 _47425_ (
    .A1(\cpuregs[25] [31]),
    .A2(_12740_),
    .ZN(_12743_)
  );
  INV_X1 _47426_ (
    .A(_12743_),
    .ZN(_12744_)
  );
  AND2_X1 _47427_ (
    .A1(_12742_),
    .A2(_12744_),
    .ZN(_12745_)
  );
  INV_X1 _47428_ (
    .A(_12745_),
    .ZN(_00509_)
  );
  AND2_X1 _47429_ (
    .A1(_12637_),
    .A2(_12724_),
    .ZN(_12746_)
  );
  INV_X1 _47430_ (
    .A(_12746_),
    .ZN(_12747_)
  );
  AND2_X1 _47431_ (
    .A1(_12628_),
    .A2(_12746_),
    .ZN(_12748_)
  );
  INV_X1 _47432_ (
    .A(_12748_),
    .ZN(_12749_)
  );
  AND2_X1 _47433_ (
    .A1(\cpuregs[24] [31]),
    .A2(_12747_),
    .ZN(_12750_)
  );
  INV_X1 _47434_ (
    .A(_12750_),
    .ZN(_12751_)
  );
  AND2_X1 _47435_ (
    .A1(_12749_),
    .A2(_12751_),
    .ZN(_12752_)
  );
  INV_X1 _47436_ (
    .A(_12752_),
    .ZN(_00510_)
  );
  AND2_X1 _47437_ (
    .A1(_21257_),
    .A2(_12646_),
    .ZN(_12753_)
  );
  AND2_X1 _47438_ (
    .A1(latched_rd[2]),
    .A2(_12753_),
    .ZN(_12754_)
  );
  AND2_X1 _47439_ (
    .A1(_12643_),
    .A2(_12754_),
    .ZN(_12755_)
  );
  INV_X1 _47440_ (
    .A(_12755_),
    .ZN(_12756_)
  );
  AND2_X1 _47441_ (
    .A1(_12628_),
    .A2(_12755_),
    .ZN(_12757_)
  );
  INV_X1 _47442_ (
    .A(_12757_),
    .ZN(_12758_)
  );
  AND2_X1 _47443_ (
    .A1(\cpuregs[23] [31]),
    .A2(_12756_),
    .ZN(_12759_)
  );
  INV_X1 _47444_ (
    .A(_12759_),
    .ZN(_12760_)
  );
  AND2_X1 _47445_ (
    .A1(_12758_),
    .A2(_12760_),
    .ZN(_12761_)
  );
  INV_X1 _47446_ (
    .A(_12761_),
    .ZN(_00511_)
  );
  AND2_X1 _47447_ (
    .A1(_12703_),
    .A2(_12754_),
    .ZN(_12762_)
  );
  INV_X1 _47448_ (
    .A(_12762_),
    .ZN(_12763_)
  );
  AND2_X1 _47449_ (
    .A1(_12628_),
    .A2(_12762_),
    .ZN(_12764_)
  );
  INV_X1 _47450_ (
    .A(_12764_),
    .ZN(_12765_)
  );
  AND2_X1 _47451_ (
    .A1(\cpuregs[22] [31]),
    .A2(_12763_),
    .ZN(_12766_)
  );
  INV_X1 _47452_ (
    .A(_12766_),
    .ZN(_12767_)
  );
  AND2_X1 _47453_ (
    .A1(_12765_),
    .A2(_12767_),
    .ZN(_12768_)
  );
  INV_X1 _47454_ (
    .A(_12768_),
    .ZN(_00512_)
  );
  AND2_X1 _47455_ (
    .A1(_12557_),
    .A2(_12754_),
    .ZN(_12769_)
  );
  INV_X1 _47456_ (
    .A(_12769_),
    .ZN(_12770_)
  );
  AND2_X1 _47457_ (
    .A1(_12628_),
    .A2(_12769_),
    .ZN(_12771_)
  );
  INV_X1 _47458_ (
    .A(_12771_),
    .ZN(_12772_)
  );
  AND2_X1 _47459_ (
    .A1(\cpuregs[21] [31]),
    .A2(_12770_),
    .ZN(_12773_)
  );
  INV_X1 _47460_ (
    .A(_12773_),
    .ZN(_12774_)
  );
  AND2_X1 _47461_ (
    .A1(_12772_),
    .A2(_12774_),
    .ZN(_12775_)
  );
  INV_X1 _47462_ (
    .A(_12775_),
    .ZN(_00513_)
  );
  AND2_X1 _47463_ (
    .A1(_12637_),
    .A2(_12754_),
    .ZN(_12776_)
  );
  INV_X1 _47464_ (
    .A(_12776_),
    .ZN(_12777_)
  );
  AND2_X1 _47465_ (
    .A1(_12628_),
    .A2(_12776_),
    .ZN(_12778_)
  );
  INV_X1 _47466_ (
    .A(_12778_),
    .ZN(_12779_)
  );
  AND2_X1 _47467_ (
    .A1(\cpuregs[20] [31]),
    .A2(_12777_),
    .ZN(_12780_)
  );
  INV_X1 _47468_ (
    .A(_12780_),
    .ZN(_12781_)
  );
  AND2_X1 _47469_ (
    .A1(_12779_),
    .A2(_12781_),
    .ZN(_12782_)
  );
  INV_X1 _47470_ (
    .A(_12782_),
    .ZN(_00514_)
  );
  AND2_X1 _47471_ (
    .A1(_12557_),
    .A2(_12679_),
    .ZN(_12783_)
  );
  INV_X1 _47472_ (
    .A(_12783_),
    .ZN(_12784_)
  );
  AND2_X1 _47473_ (
    .A1(_12628_),
    .A2(_12783_),
    .ZN(_12785_)
  );
  INV_X1 _47474_ (
    .A(_12785_),
    .ZN(_12786_)
  );
  AND2_X1 _47475_ (
    .A1(\cpuregs[1] [31]),
    .A2(_12784_),
    .ZN(_12787_)
  );
  INV_X1 _47476_ (
    .A(_12787_),
    .ZN(_12788_)
  );
  AND2_X1 _47477_ (
    .A1(_12786_),
    .A2(_12788_),
    .ZN(_12789_)
  );
  INV_X1 _47478_ (
    .A(_12789_),
    .ZN(_00515_)
  );
  AND2_X1 _47479_ (
    .A1(_21256_),
    .A2(_12753_),
    .ZN(_12790_)
  );
  AND2_X1 _47480_ (
    .A1(_12643_),
    .A2(_12790_),
    .ZN(_12791_)
  );
  INV_X1 _47481_ (
    .A(_12791_),
    .ZN(_12792_)
  );
  AND2_X1 _47482_ (
    .A1(_12628_),
    .A2(_12791_),
    .ZN(_12793_)
  );
  INV_X1 _47483_ (
    .A(_12793_),
    .ZN(_12794_)
  );
  AND2_X1 _47484_ (
    .A1(\cpuregs[19] [31]),
    .A2(_12792_),
    .ZN(_12795_)
  );
  INV_X1 _47485_ (
    .A(_12795_),
    .ZN(_12796_)
  );
  AND2_X1 _47486_ (
    .A1(_12794_),
    .A2(_12796_),
    .ZN(_12797_)
  );
  INV_X1 _47487_ (
    .A(_12797_),
    .ZN(_00516_)
  );
  AND2_X1 _47488_ (
    .A1(_12703_),
    .A2(_12790_),
    .ZN(_12798_)
  );
  INV_X1 _47489_ (
    .A(_12798_),
    .ZN(_12799_)
  );
  AND2_X1 _47490_ (
    .A1(_12628_),
    .A2(_12798_),
    .ZN(_12800_)
  );
  INV_X1 _47491_ (
    .A(_12800_),
    .ZN(_12801_)
  );
  AND2_X1 _47492_ (
    .A1(\cpuregs[18] [31]),
    .A2(_12799_),
    .ZN(_12802_)
  );
  INV_X1 _47493_ (
    .A(_12802_),
    .ZN(_12803_)
  );
  AND2_X1 _47494_ (
    .A1(_12801_),
    .A2(_12803_),
    .ZN(_12804_)
  );
  INV_X1 _47495_ (
    .A(_12804_),
    .ZN(_00517_)
  );
  AND2_X1 _47496_ (
    .A1(_12557_),
    .A2(_12790_),
    .ZN(_12805_)
  );
  INV_X1 _47497_ (
    .A(_12805_),
    .ZN(_12806_)
  );
  AND2_X1 _47498_ (
    .A1(_12628_),
    .A2(_12805_),
    .ZN(_12807_)
  );
  INV_X1 _47499_ (
    .A(_12807_),
    .ZN(_12808_)
  );
  AND2_X1 _47500_ (
    .A1(\cpuregs[17] [31]),
    .A2(_12806_),
    .ZN(_12809_)
  );
  INV_X1 _47501_ (
    .A(_12809_),
    .ZN(_12810_)
  );
  AND2_X1 _47502_ (
    .A1(_12808_),
    .A2(_12810_),
    .ZN(_12811_)
  );
  INV_X1 _47503_ (
    .A(_12811_),
    .ZN(_00518_)
  );
  AND2_X1 _47504_ (
    .A1(_12637_),
    .A2(_12790_),
    .ZN(_12812_)
  );
  INV_X1 _47505_ (
    .A(_12812_),
    .ZN(_12813_)
  );
  AND2_X1 _47506_ (
    .A1(_12628_),
    .A2(_12812_),
    .ZN(_12814_)
  );
  INV_X1 _47507_ (
    .A(_12814_),
    .ZN(_12815_)
  );
  AND2_X1 _47508_ (
    .A1(\cpuregs[16] [31]),
    .A2(_12813_),
    .ZN(_12816_)
  );
  INV_X1 _47509_ (
    .A(_12816_),
    .ZN(_12817_)
  );
  AND2_X1 _47510_ (
    .A1(_12815_),
    .A2(_12817_),
    .ZN(_12818_)
  );
  INV_X1 _47511_ (
    .A(_12818_),
    .ZN(_00519_)
  );
  AND2_X1 _47512_ (
    .A1(latched_rd[2]),
    .A2(_21258_),
    .ZN(_12819_)
  );
  AND2_X1 _47513_ (
    .A1(_12547_),
    .A2(_12819_),
    .ZN(_12820_)
  );
  AND2_X1 _47514_ (
    .A1(_12643_),
    .A2(_12820_),
    .ZN(_12821_)
  );
  INV_X1 _47515_ (
    .A(_12821_),
    .ZN(_12822_)
  );
  AND2_X1 _47516_ (
    .A1(\cpuregs[15] [31]),
    .A2(_12822_),
    .ZN(_12823_)
  );
  INV_X1 _47517_ (
    .A(_12823_),
    .ZN(_12824_)
  );
  AND2_X1 _47518_ (
    .A1(_12628_),
    .A2(_12821_),
    .ZN(_12825_)
  );
  INV_X1 _47519_ (
    .A(_12825_),
    .ZN(_12826_)
  );
  AND2_X1 _47520_ (
    .A1(_12824_),
    .A2(_12826_),
    .ZN(_12827_)
  );
  INV_X1 _47521_ (
    .A(_12827_),
    .ZN(_00520_)
  );
  AND2_X1 _47522_ (
    .A1(_12657_),
    .A2(_12820_),
    .ZN(_12828_)
  );
  INV_X1 _47523_ (
    .A(_12828_),
    .ZN(_12829_)
  );
  AND2_X1 _47524_ (
    .A1(\cpuregs[14] [31]),
    .A2(_12829_),
    .ZN(_12830_)
  );
  INV_X1 _47525_ (
    .A(_12830_),
    .ZN(_12831_)
  );
  AND2_X1 _47526_ (
    .A1(_12628_),
    .A2(_12828_),
    .ZN(_12832_)
  );
  INV_X1 _47527_ (
    .A(_12832_),
    .ZN(_12833_)
  );
  AND2_X1 _47528_ (
    .A1(_12831_),
    .A2(_12833_),
    .ZN(_12834_)
  );
  INV_X1 _47529_ (
    .A(_12834_),
    .ZN(_00521_)
  );
  AND2_X1 _47530_ (
    .A1(_12557_),
    .A2(_12820_),
    .ZN(_12835_)
  );
  INV_X1 _47531_ (
    .A(_12835_),
    .ZN(_12836_)
  );
  AND2_X1 _47532_ (
    .A1(\cpuregs[13] [31]),
    .A2(_12836_),
    .ZN(_12837_)
  );
  INV_X1 _47533_ (
    .A(_12837_),
    .ZN(_12838_)
  );
  AND2_X1 _47534_ (
    .A1(_12628_),
    .A2(_12835_),
    .ZN(_12839_)
  );
  INV_X1 _47535_ (
    .A(_12839_),
    .ZN(_12840_)
  );
  AND2_X1 _47536_ (
    .A1(_12838_),
    .A2(_12840_),
    .ZN(_12841_)
  );
  INV_X1 _47537_ (
    .A(_12841_),
    .ZN(_00522_)
  );
  AND2_X1 _47538_ (
    .A1(_12549_),
    .A2(_12820_),
    .ZN(_12842_)
  );
  INV_X1 _47539_ (
    .A(_12842_),
    .ZN(_12843_)
  );
  AND2_X1 _47540_ (
    .A1(\cpuregs[12] [31]),
    .A2(_12843_),
    .ZN(_12844_)
  );
  INV_X1 _47541_ (
    .A(_12844_),
    .ZN(_12845_)
  );
  AND2_X1 _47542_ (
    .A1(_12628_),
    .A2(_12842_),
    .ZN(_12846_)
  );
  INV_X1 _47543_ (
    .A(_12846_),
    .ZN(_12847_)
  );
  AND2_X1 _47544_ (
    .A1(_12845_),
    .A2(_12847_),
    .ZN(_12848_)
  );
  INV_X1 _47545_ (
    .A(_12848_),
    .ZN(_00523_)
  );
  AND2_X1 _47546_ (
    .A1(_12558_),
    .A2(_12643_),
    .ZN(_12849_)
  );
  INV_X1 _47547_ (
    .A(_12849_),
    .ZN(_12850_)
  );
  AND2_X1 _47548_ (
    .A1(_12628_),
    .A2(_12849_),
    .ZN(_12851_)
  );
  INV_X1 _47549_ (
    .A(_12851_),
    .ZN(_12852_)
  );
  AND2_X1 _47550_ (
    .A1(\cpuregs[11] [31]),
    .A2(_12850_),
    .ZN(_12853_)
  );
  INV_X1 _47551_ (
    .A(_12853_),
    .ZN(_12854_)
  );
  AND2_X1 _47552_ (
    .A1(_12852_),
    .A2(_12854_),
    .ZN(_12855_)
  );
  INV_X1 _47553_ (
    .A(_12855_),
    .ZN(_00524_)
  );
  AND2_X1 _47554_ (
    .A1(_12558_),
    .A2(_12657_),
    .ZN(_12856_)
  );
  INV_X1 _47555_ (
    .A(_12856_),
    .ZN(_12857_)
  );
  AND2_X1 _47556_ (
    .A1(_12628_),
    .A2(_12856_),
    .ZN(_12858_)
  );
  INV_X1 _47557_ (
    .A(_12858_),
    .ZN(_12859_)
  );
  AND2_X1 _47558_ (
    .A1(\cpuregs[10] [31]),
    .A2(_12857_),
    .ZN(_12860_)
  );
  INV_X1 _47559_ (
    .A(_12860_),
    .ZN(_12861_)
  );
  AND2_X1 _47560_ (
    .A1(_12859_),
    .A2(_12861_),
    .ZN(_12862_)
  );
  INV_X1 _47561_ (
    .A(_12862_),
    .ZN(_00525_)
  );
  AND2_X1 _47562_ (
    .A1(reg_next_pc[0]),
    .A2(latched_branch),
    .ZN(_12863_)
  );
  INV_X1 _47563_ (
    .A(_12863_),
    .ZN(_12864_)
  );
  AND2_X1 _47564_ (
    .A1(_21067_),
    .A2(_22110_),
    .ZN(_12865_)
  );
  INV_X1 _47565_ (
    .A(_12865_),
    .ZN(_12866_)
  );
  AND2_X1 _47566_ (
    .A1(latched_stalu),
    .A2(_22111_),
    .ZN(_12867_)
  );
  INV_X1 _47567_ (
    .A(_12867_),
    .ZN(_12868_)
  );
  AND2_X1 _47568_ (
    .A1(_12542_),
    .A2(_12868_),
    .ZN(_12869_)
  );
  AND2_X1 _47569_ (
    .A1(_12866_),
    .A2(_12869_),
    .ZN(_12870_)
  );
  INV_X1 _47570_ (
    .A(_12870_),
    .ZN(_12871_)
  );
  AND2_X1 _47571_ (
    .A1(_12864_),
    .A2(_12871_),
    .ZN(_12872_)
  );
  INV_X1 _47572_ (
    .A(_12872_),
    .ZN(_12873_)
  );
  AND2_X1 _47573_ (
    .A1(_12555_),
    .A2(_12873_),
    .ZN(_12874_)
  );
  AND2_X1 _47574_ (
    .A1(_12755_),
    .A2(_12874_),
    .ZN(_12875_)
  );
  INV_X1 _47575_ (
    .A(_12875_),
    .ZN(_12876_)
  );
  AND2_X1 _47576_ (
    .A1(\cpuregs[23] [0]),
    .A2(_12756_),
    .ZN(_12877_)
  );
  INV_X1 _47577_ (
    .A(_12877_),
    .ZN(_12878_)
  );
  AND2_X1 _47578_ (
    .A1(_12876_),
    .A2(_12878_),
    .ZN(_12879_)
  );
  INV_X1 _47579_ (
    .A(_12879_),
    .ZN(_00527_)
  );
  AND2_X1 _47580_ (
    .A1(_02921_),
    .A2(_12542_),
    .ZN(_12880_)
  );
  INV_X1 _47581_ (
    .A(_12880_),
    .ZN(_12881_)
  );
  AND2_X1 _47582_ (
    .A1(latched_branch),
    .A2(reg_pc[1]),
    .ZN(_12882_)
  );
  INV_X1 _47583_ (
    .A(_12882_),
    .ZN(_12883_)
  );
  AND2_X1 _47584_ (
    .A1(_12881_),
    .A2(_12883_),
    .ZN(_12884_)
  );
  INV_X1 _47585_ (
    .A(_12884_),
    .ZN(_12885_)
  );
  AND2_X1 _47586_ (
    .A1(_12555_),
    .A2(_12885_),
    .ZN(_12886_)
  );
  AND2_X1 _47587_ (
    .A1(_12755_),
    .A2(_12886_),
    .ZN(_12887_)
  );
  INV_X1 _47588_ (
    .A(_12887_),
    .ZN(_12888_)
  );
  AND2_X1 _47589_ (
    .A1(\cpuregs[23] [1]),
    .A2(_12756_),
    .ZN(_12889_)
  );
  INV_X1 _47590_ (
    .A(_12889_),
    .ZN(_12890_)
  );
  AND2_X1 _47591_ (
    .A1(_12888_),
    .A2(_12890_),
    .ZN(_12891_)
  );
  INV_X1 _47592_ (
    .A(_12891_),
    .ZN(_00528_)
  );
  AND2_X1 _47593_ (
    .A1(\cpuregs[23] [2]),
    .A2(_12756_),
    .ZN(_12892_)
  );
  INV_X1 _47594_ (
    .A(_12892_),
    .ZN(_12893_)
  );
  AND2_X1 _47595_ (
    .A1(_02938_),
    .A2(_12542_),
    .ZN(_12894_)
  );
  INV_X1 _47596_ (
    .A(_12894_),
    .ZN(_12895_)
  );
  AND2_X1 _47597_ (
    .A1(latched_branch),
    .A2(_29145_[98]),
    .ZN(_12896_)
  );
  INV_X1 _47598_ (
    .A(_12896_),
    .ZN(_12897_)
  );
  AND2_X1 _47599_ (
    .A1(_12895_),
    .A2(_12897_),
    .ZN(_12898_)
  );
  INV_X1 _47600_ (
    .A(_12898_),
    .ZN(_12899_)
  );
  AND2_X1 _47601_ (
    .A1(_12555_),
    .A2(_12899_),
    .ZN(_12900_)
  );
  AND2_X1 _47602_ (
    .A1(_12755_),
    .A2(_12900_),
    .ZN(_12901_)
  );
  INV_X1 _47603_ (
    .A(_12901_),
    .ZN(_12902_)
  );
  AND2_X1 _47604_ (
    .A1(_12893_),
    .A2(_12902_),
    .ZN(_12903_)
  );
  INV_X1 _47605_ (
    .A(_12903_),
    .ZN(_00529_)
  );
  AND2_X1 _47606_ (
    .A1(_02954_),
    .A2(_12542_),
    .ZN(_12904_)
  );
  INV_X1 _47607_ (
    .A(_12904_),
    .ZN(_12905_)
  );
  AND2_X1 _47608_ (
    .A1(_21101_),
    .A2(_21102_),
    .ZN(_12906_)
  );
  INV_X1 _47609_ (
    .A(_12906_),
    .ZN(_12907_)
  );
  AND2_X1 _47610_ (
    .A1(latched_branch),
    .A2(_12564_),
    .ZN(_12908_)
  );
  AND2_X1 _47611_ (
    .A1(_12907_),
    .A2(_12908_),
    .ZN(_12909_)
  );
  INV_X1 _47612_ (
    .A(_12909_),
    .ZN(_12910_)
  );
  AND2_X1 _47613_ (
    .A1(_12905_),
    .A2(_12910_),
    .ZN(_12911_)
  );
  INV_X1 _47614_ (
    .A(_12911_),
    .ZN(_12912_)
  );
  AND2_X1 _47615_ (
    .A1(_12555_),
    .A2(_12912_),
    .ZN(_12913_)
  );
  AND2_X1 _47616_ (
    .A1(_12755_),
    .A2(_12913_),
    .ZN(_12914_)
  );
  INV_X1 _47617_ (
    .A(_12914_),
    .ZN(_12915_)
  );
  AND2_X1 _47618_ (
    .A1(\cpuregs[23] [3]),
    .A2(_12756_),
    .ZN(_12916_)
  );
  INV_X1 _47619_ (
    .A(_12916_),
    .ZN(_12917_)
  );
  AND2_X1 _47620_ (
    .A1(_12915_),
    .A2(_12917_),
    .ZN(_12918_)
  );
  INV_X1 _47621_ (
    .A(_12918_),
    .ZN(_00530_)
  );
  AND2_X1 _47622_ (
    .A1(_02970_),
    .A2(_12542_),
    .ZN(_12919_)
  );
  INV_X1 _47623_ (
    .A(_12919_),
    .ZN(_12920_)
  );
  AND2_X1 _47624_ (
    .A1(_21100_),
    .A2(_12564_),
    .ZN(_12921_)
  );
  INV_X1 _47625_ (
    .A(_12921_),
    .ZN(_12922_)
  );
  AND2_X1 _47626_ (
    .A1(latched_branch),
    .A2(_12566_),
    .ZN(_12923_)
  );
  AND2_X1 _47627_ (
    .A1(_12922_),
    .A2(_12923_),
    .ZN(_12924_)
  );
  INV_X1 _47628_ (
    .A(_12924_),
    .ZN(_12925_)
  );
  AND2_X1 _47629_ (
    .A1(_12920_),
    .A2(_12925_),
    .ZN(_12926_)
  );
  INV_X1 _47630_ (
    .A(_12926_),
    .ZN(_12927_)
  );
  AND2_X1 _47631_ (
    .A1(_12555_),
    .A2(_12927_),
    .ZN(_12928_)
  );
  AND2_X1 _47632_ (
    .A1(_12755_),
    .A2(_12928_),
    .ZN(_12929_)
  );
  INV_X1 _47633_ (
    .A(_12929_),
    .ZN(_12930_)
  );
  AND2_X1 _47634_ (
    .A1(\cpuregs[23] [4]),
    .A2(_12756_),
    .ZN(_12931_)
  );
  INV_X1 _47635_ (
    .A(_12931_),
    .ZN(_12932_)
  );
  AND2_X1 _47636_ (
    .A1(_12930_),
    .A2(_12932_),
    .ZN(_12933_)
  );
  INV_X1 _47637_ (
    .A(_12933_),
    .ZN(_00531_)
  );
  AND2_X1 _47638_ (
    .A1(_02986_),
    .A2(_12542_),
    .ZN(_12934_)
  );
  INV_X1 _47639_ (
    .A(_12934_),
    .ZN(_12935_)
  );
  AND2_X1 _47640_ (
    .A1(_21099_),
    .A2(_12566_),
    .ZN(_12936_)
  );
  INV_X1 _47641_ (
    .A(_12936_),
    .ZN(_12937_)
  );
  AND2_X1 _47642_ (
    .A1(latched_branch),
    .A2(_12568_),
    .ZN(_12938_)
  );
  AND2_X1 _47643_ (
    .A1(_12937_),
    .A2(_12938_),
    .ZN(_12939_)
  );
  INV_X1 _47644_ (
    .A(_12939_),
    .ZN(_12940_)
  );
  AND2_X1 _47645_ (
    .A1(_12935_),
    .A2(_12940_),
    .ZN(_12941_)
  );
  INV_X1 _47646_ (
    .A(_12941_),
    .ZN(_12942_)
  );
  AND2_X1 _47647_ (
    .A1(_12555_),
    .A2(_12942_),
    .ZN(_12943_)
  );
  AND2_X1 _47648_ (
    .A1(_12755_),
    .A2(_12943_),
    .ZN(_12944_)
  );
  INV_X1 _47649_ (
    .A(_12944_),
    .ZN(_12945_)
  );
  AND2_X1 _47650_ (
    .A1(\cpuregs[23] [5]),
    .A2(_12756_),
    .ZN(_12946_)
  );
  INV_X1 _47651_ (
    .A(_12946_),
    .ZN(_12947_)
  );
  AND2_X1 _47652_ (
    .A1(_12945_),
    .A2(_12947_),
    .ZN(_12948_)
  );
  INV_X1 _47653_ (
    .A(_12948_),
    .ZN(_00532_)
  );
  AND2_X1 _47654_ (
    .A1(_03002_),
    .A2(_12542_),
    .ZN(_12949_)
  );
  INV_X1 _47655_ (
    .A(_12949_),
    .ZN(_12950_)
  );
  AND2_X1 _47656_ (
    .A1(_21098_),
    .A2(_12568_),
    .ZN(_12951_)
  );
  INV_X1 _47657_ (
    .A(_12951_),
    .ZN(_12952_)
  );
  AND2_X1 _47658_ (
    .A1(latched_branch),
    .A2(_12570_),
    .ZN(_12953_)
  );
  AND2_X1 _47659_ (
    .A1(_12952_),
    .A2(_12953_),
    .ZN(_12954_)
  );
  INV_X1 _47660_ (
    .A(_12954_),
    .ZN(_12955_)
  );
  AND2_X1 _47661_ (
    .A1(_12950_),
    .A2(_12955_),
    .ZN(_12956_)
  );
  INV_X1 _47662_ (
    .A(_12956_),
    .ZN(_12957_)
  );
  AND2_X1 _47663_ (
    .A1(_12555_),
    .A2(_12957_),
    .ZN(_12958_)
  );
  AND2_X1 _47664_ (
    .A1(_12755_),
    .A2(_12958_),
    .ZN(_12959_)
  );
  INV_X1 _47665_ (
    .A(_12959_),
    .ZN(_12960_)
  );
  AND2_X1 _47666_ (
    .A1(\cpuregs[23] [6]),
    .A2(_12756_),
    .ZN(_12961_)
  );
  INV_X1 _47667_ (
    .A(_12961_),
    .ZN(_12962_)
  );
  AND2_X1 _47668_ (
    .A1(_12960_),
    .A2(_12962_),
    .ZN(_12963_)
  );
  INV_X1 _47669_ (
    .A(_12963_),
    .ZN(_00533_)
  );
  AND2_X1 _47670_ (
    .A1(_03018_),
    .A2(_12542_),
    .ZN(_12964_)
  );
  INV_X1 _47671_ (
    .A(_12964_),
    .ZN(_12965_)
  );
  AND2_X1 _47672_ (
    .A1(_21097_),
    .A2(_12570_),
    .ZN(_12966_)
  );
  INV_X1 _47673_ (
    .A(_12966_),
    .ZN(_12967_)
  );
  AND2_X1 _47674_ (
    .A1(latched_branch),
    .A2(_12572_),
    .ZN(_12968_)
  );
  AND2_X1 _47675_ (
    .A1(_12967_),
    .A2(_12968_),
    .ZN(_12969_)
  );
  INV_X1 _47676_ (
    .A(_12969_),
    .ZN(_12970_)
  );
  AND2_X1 _47677_ (
    .A1(_12965_),
    .A2(_12970_),
    .ZN(_12971_)
  );
  INV_X1 _47678_ (
    .A(_12971_),
    .ZN(_12972_)
  );
  AND2_X1 _47679_ (
    .A1(_12555_),
    .A2(_12972_),
    .ZN(_12973_)
  );
  AND2_X1 _47680_ (
    .A1(_12755_),
    .A2(_12973_),
    .ZN(_12974_)
  );
  INV_X1 _47681_ (
    .A(_12974_),
    .ZN(_12975_)
  );
  AND2_X1 _47682_ (
    .A1(\cpuregs[23] [7]),
    .A2(_12756_),
    .ZN(_12976_)
  );
  INV_X1 _47683_ (
    .A(_12976_),
    .ZN(_12977_)
  );
  AND2_X1 _47684_ (
    .A1(_12975_),
    .A2(_12977_),
    .ZN(_12978_)
  );
  INV_X1 _47685_ (
    .A(_12978_),
    .ZN(_00534_)
  );
  AND2_X1 _47686_ (
    .A1(_03034_),
    .A2(_12542_),
    .ZN(_12979_)
  );
  INV_X1 _47687_ (
    .A(_12979_),
    .ZN(_12980_)
  );
  AND2_X1 _47688_ (
    .A1(_21096_),
    .A2(_12572_),
    .ZN(_12981_)
  );
  INV_X1 _47689_ (
    .A(_12981_),
    .ZN(_12982_)
  );
  AND2_X1 _47690_ (
    .A1(latched_branch),
    .A2(_12574_),
    .ZN(_12983_)
  );
  AND2_X1 _47691_ (
    .A1(_12982_),
    .A2(_12983_),
    .ZN(_12984_)
  );
  INV_X1 _47692_ (
    .A(_12984_),
    .ZN(_12985_)
  );
  AND2_X1 _47693_ (
    .A1(_12980_),
    .A2(_12985_),
    .ZN(_12986_)
  );
  INV_X1 _47694_ (
    .A(_12986_),
    .ZN(_12987_)
  );
  AND2_X1 _47695_ (
    .A1(_12555_),
    .A2(_12987_),
    .ZN(_12988_)
  );
  AND2_X1 _47696_ (
    .A1(_12755_),
    .A2(_12988_),
    .ZN(_12989_)
  );
  INV_X1 _47697_ (
    .A(_12989_),
    .ZN(_12990_)
  );
  AND2_X1 _47698_ (
    .A1(\cpuregs[23] [8]),
    .A2(_12756_),
    .ZN(_12991_)
  );
  INV_X1 _47699_ (
    .A(_12991_),
    .ZN(_12992_)
  );
  AND2_X1 _47700_ (
    .A1(_12990_),
    .A2(_12992_),
    .ZN(_12993_)
  );
  INV_X1 _47701_ (
    .A(_12993_),
    .ZN(_00535_)
  );
  AND2_X1 _47702_ (
    .A1(_03050_),
    .A2(_12542_),
    .ZN(_12994_)
  );
  INV_X1 _47703_ (
    .A(_12994_),
    .ZN(_12995_)
  );
  AND2_X1 _47704_ (
    .A1(_21095_),
    .A2(_12574_),
    .ZN(_12996_)
  );
  INV_X1 _47705_ (
    .A(_12996_),
    .ZN(_12997_)
  );
  AND2_X1 _47706_ (
    .A1(latched_branch),
    .A2(_12576_),
    .ZN(_12998_)
  );
  AND2_X1 _47707_ (
    .A1(_12997_),
    .A2(_12998_),
    .ZN(_12999_)
  );
  INV_X1 _47708_ (
    .A(_12999_),
    .ZN(_13000_)
  );
  AND2_X1 _47709_ (
    .A1(_12995_),
    .A2(_13000_),
    .ZN(_13001_)
  );
  INV_X1 _47710_ (
    .A(_13001_),
    .ZN(_13002_)
  );
  AND2_X1 _47711_ (
    .A1(_12555_),
    .A2(_13002_),
    .ZN(_13003_)
  );
  AND2_X1 _47712_ (
    .A1(_12755_),
    .A2(_13003_),
    .ZN(_13004_)
  );
  INV_X1 _47713_ (
    .A(_13004_),
    .ZN(_13005_)
  );
  AND2_X1 _47714_ (
    .A1(\cpuregs[23] [9]),
    .A2(_12756_),
    .ZN(_13006_)
  );
  INV_X1 _47715_ (
    .A(_13006_),
    .ZN(_13007_)
  );
  AND2_X1 _47716_ (
    .A1(_13005_),
    .A2(_13007_),
    .ZN(_13008_)
  );
  INV_X1 _47717_ (
    .A(_13008_),
    .ZN(_00536_)
  );
  AND2_X1 _47718_ (
    .A1(_03066_),
    .A2(_12542_),
    .ZN(_13009_)
  );
  INV_X1 _47719_ (
    .A(_13009_),
    .ZN(_13010_)
  );
  AND2_X1 _47720_ (
    .A1(_21094_),
    .A2(_12576_),
    .ZN(_13011_)
  );
  INV_X1 _47721_ (
    .A(_13011_),
    .ZN(_13012_)
  );
  AND2_X1 _47722_ (
    .A1(latched_branch),
    .A2(_12578_),
    .ZN(_13013_)
  );
  AND2_X1 _47723_ (
    .A1(_13012_),
    .A2(_13013_),
    .ZN(_13014_)
  );
  INV_X1 _47724_ (
    .A(_13014_),
    .ZN(_13015_)
  );
  AND2_X1 _47725_ (
    .A1(_13010_),
    .A2(_13015_),
    .ZN(_13016_)
  );
  INV_X1 _47726_ (
    .A(_13016_),
    .ZN(_13017_)
  );
  AND2_X1 _47727_ (
    .A1(_12555_),
    .A2(_13017_),
    .ZN(_13018_)
  );
  AND2_X1 _47728_ (
    .A1(_12755_),
    .A2(_13018_),
    .ZN(_13019_)
  );
  INV_X1 _47729_ (
    .A(_13019_),
    .ZN(_13020_)
  );
  AND2_X1 _47730_ (
    .A1(\cpuregs[23] [10]),
    .A2(_12756_),
    .ZN(_13021_)
  );
  INV_X1 _47731_ (
    .A(_13021_),
    .ZN(_13022_)
  );
  AND2_X1 _47732_ (
    .A1(_13020_),
    .A2(_13022_),
    .ZN(_13023_)
  );
  INV_X1 _47733_ (
    .A(_13023_),
    .ZN(_00537_)
  );
  AND2_X1 _47734_ (
    .A1(_03082_),
    .A2(_12542_),
    .ZN(_13024_)
  );
  INV_X1 _47735_ (
    .A(_13024_),
    .ZN(_13025_)
  );
  AND2_X1 _47736_ (
    .A1(_21093_),
    .A2(_12578_),
    .ZN(_13026_)
  );
  INV_X1 _47737_ (
    .A(_13026_),
    .ZN(_13027_)
  );
  AND2_X1 _47738_ (
    .A1(latched_branch),
    .A2(_12580_),
    .ZN(_13028_)
  );
  AND2_X1 _47739_ (
    .A1(_13027_),
    .A2(_13028_),
    .ZN(_13029_)
  );
  INV_X1 _47740_ (
    .A(_13029_),
    .ZN(_13030_)
  );
  AND2_X1 _47741_ (
    .A1(_13025_),
    .A2(_13030_),
    .ZN(_13031_)
  );
  INV_X1 _47742_ (
    .A(_13031_),
    .ZN(_13032_)
  );
  AND2_X1 _47743_ (
    .A1(_12555_),
    .A2(_13032_),
    .ZN(_13033_)
  );
  AND2_X1 _47744_ (
    .A1(_12755_),
    .A2(_13033_),
    .ZN(_13034_)
  );
  INV_X1 _47745_ (
    .A(_13034_),
    .ZN(_13035_)
  );
  AND2_X1 _47746_ (
    .A1(\cpuregs[23] [11]),
    .A2(_12756_),
    .ZN(_13036_)
  );
  INV_X1 _47747_ (
    .A(_13036_),
    .ZN(_13037_)
  );
  AND2_X1 _47748_ (
    .A1(_13035_),
    .A2(_13037_),
    .ZN(_13038_)
  );
  INV_X1 _47749_ (
    .A(_13038_),
    .ZN(_00538_)
  );
  AND2_X1 _47750_ (
    .A1(_03098_),
    .A2(_12542_),
    .ZN(_13039_)
  );
  INV_X1 _47751_ (
    .A(_13039_),
    .ZN(_13040_)
  );
  AND2_X1 _47752_ (
    .A1(_21092_),
    .A2(_12580_),
    .ZN(_13041_)
  );
  INV_X1 _47753_ (
    .A(_13041_),
    .ZN(_13042_)
  );
  AND2_X1 _47754_ (
    .A1(latched_branch),
    .A2(_12582_),
    .ZN(_13043_)
  );
  AND2_X1 _47755_ (
    .A1(_13042_),
    .A2(_13043_),
    .ZN(_13044_)
  );
  INV_X1 _47756_ (
    .A(_13044_),
    .ZN(_13045_)
  );
  AND2_X1 _47757_ (
    .A1(_13040_),
    .A2(_13045_),
    .ZN(_13046_)
  );
  INV_X1 _47758_ (
    .A(_13046_),
    .ZN(_13047_)
  );
  AND2_X1 _47759_ (
    .A1(_12555_),
    .A2(_13047_),
    .ZN(_13048_)
  );
  AND2_X1 _47760_ (
    .A1(_12755_),
    .A2(_13048_),
    .ZN(_13049_)
  );
  INV_X1 _47761_ (
    .A(_13049_),
    .ZN(_13050_)
  );
  AND2_X1 _47762_ (
    .A1(\cpuregs[23] [12]),
    .A2(_12756_),
    .ZN(_13051_)
  );
  INV_X1 _47763_ (
    .A(_13051_),
    .ZN(_13052_)
  );
  AND2_X1 _47764_ (
    .A1(_13050_),
    .A2(_13052_),
    .ZN(_13053_)
  );
  INV_X1 _47765_ (
    .A(_13053_),
    .ZN(_00539_)
  );
  AND2_X1 _47766_ (
    .A1(_03114_),
    .A2(_12542_),
    .ZN(_13054_)
  );
  INV_X1 _47767_ (
    .A(_13054_),
    .ZN(_13055_)
  );
  AND2_X1 _47768_ (
    .A1(_21091_),
    .A2(_12582_),
    .ZN(_13056_)
  );
  INV_X1 _47769_ (
    .A(_13056_),
    .ZN(_13057_)
  );
  AND2_X1 _47770_ (
    .A1(latched_branch),
    .A2(_12584_),
    .ZN(_13058_)
  );
  AND2_X1 _47771_ (
    .A1(_13057_),
    .A2(_13058_),
    .ZN(_13059_)
  );
  INV_X1 _47772_ (
    .A(_13059_),
    .ZN(_13060_)
  );
  AND2_X1 _47773_ (
    .A1(_13055_),
    .A2(_13060_),
    .ZN(_13061_)
  );
  INV_X1 _47774_ (
    .A(_13061_),
    .ZN(_13062_)
  );
  AND2_X1 _47775_ (
    .A1(_12555_),
    .A2(_13062_),
    .ZN(_13063_)
  );
  AND2_X1 _47776_ (
    .A1(_12755_),
    .A2(_13063_),
    .ZN(_13064_)
  );
  INV_X1 _47777_ (
    .A(_13064_),
    .ZN(_13065_)
  );
  AND2_X1 _47778_ (
    .A1(\cpuregs[23] [13]),
    .A2(_12756_),
    .ZN(_13066_)
  );
  INV_X1 _47779_ (
    .A(_13066_),
    .ZN(_13067_)
  );
  AND2_X1 _47780_ (
    .A1(_13065_),
    .A2(_13067_),
    .ZN(_13068_)
  );
  INV_X1 _47781_ (
    .A(_13068_),
    .ZN(_00540_)
  );
  AND2_X1 _47782_ (
    .A1(_03130_),
    .A2(_12542_),
    .ZN(_13069_)
  );
  INV_X1 _47783_ (
    .A(_13069_),
    .ZN(_13070_)
  );
  AND2_X1 _47784_ (
    .A1(_21090_),
    .A2(_12584_),
    .ZN(_13071_)
  );
  INV_X1 _47785_ (
    .A(_13071_),
    .ZN(_13072_)
  );
  AND2_X1 _47786_ (
    .A1(latched_branch),
    .A2(_12586_),
    .ZN(_13073_)
  );
  AND2_X1 _47787_ (
    .A1(_13072_),
    .A2(_13073_),
    .ZN(_13074_)
  );
  INV_X1 _47788_ (
    .A(_13074_),
    .ZN(_13075_)
  );
  AND2_X1 _47789_ (
    .A1(_13070_),
    .A2(_13075_),
    .ZN(_13076_)
  );
  INV_X1 _47790_ (
    .A(_13076_),
    .ZN(_13077_)
  );
  AND2_X1 _47791_ (
    .A1(_12555_),
    .A2(_13077_),
    .ZN(_13078_)
  );
  AND2_X1 _47792_ (
    .A1(_12755_),
    .A2(_13078_),
    .ZN(_13079_)
  );
  INV_X1 _47793_ (
    .A(_13079_),
    .ZN(_13080_)
  );
  AND2_X1 _47794_ (
    .A1(\cpuregs[23] [14]),
    .A2(_12756_),
    .ZN(_13081_)
  );
  INV_X1 _47795_ (
    .A(_13081_),
    .ZN(_13082_)
  );
  AND2_X1 _47796_ (
    .A1(_13080_),
    .A2(_13082_),
    .ZN(_13083_)
  );
  INV_X1 _47797_ (
    .A(_13083_),
    .ZN(_00541_)
  );
  AND2_X1 _47798_ (
    .A1(_03146_),
    .A2(_12542_),
    .ZN(_13084_)
  );
  INV_X1 _47799_ (
    .A(_13084_),
    .ZN(_13085_)
  );
  AND2_X1 _47800_ (
    .A1(_21089_),
    .A2(_12586_),
    .ZN(_13086_)
  );
  INV_X1 _47801_ (
    .A(_13086_),
    .ZN(_13087_)
  );
  AND2_X1 _47802_ (
    .A1(latched_branch),
    .A2(_12588_),
    .ZN(_13088_)
  );
  AND2_X1 _47803_ (
    .A1(_13087_),
    .A2(_13088_),
    .ZN(_13089_)
  );
  INV_X1 _47804_ (
    .A(_13089_),
    .ZN(_13090_)
  );
  AND2_X1 _47805_ (
    .A1(_13085_),
    .A2(_13090_),
    .ZN(_13091_)
  );
  INV_X1 _47806_ (
    .A(_13091_),
    .ZN(_13092_)
  );
  AND2_X1 _47807_ (
    .A1(_12555_),
    .A2(_13092_),
    .ZN(_13093_)
  );
  AND2_X1 _47808_ (
    .A1(_12755_),
    .A2(_13093_),
    .ZN(_13094_)
  );
  INV_X1 _47809_ (
    .A(_13094_),
    .ZN(_13095_)
  );
  AND2_X1 _47810_ (
    .A1(\cpuregs[23] [15]),
    .A2(_12756_),
    .ZN(_13096_)
  );
  INV_X1 _47811_ (
    .A(_13096_),
    .ZN(_13097_)
  );
  AND2_X1 _47812_ (
    .A1(_13095_),
    .A2(_13097_),
    .ZN(_13098_)
  );
  INV_X1 _47813_ (
    .A(_13098_),
    .ZN(_00542_)
  );
  AND2_X1 _47814_ (
    .A1(_03162_),
    .A2(_12542_),
    .ZN(_13099_)
  );
  INV_X1 _47815_ (
    .A(_13099_),
    .ZN(_13100_)
  );
  AND2_X1 _47816_ (
    .A1(_21088_),
    .A2(_12588_),
    .ZN(_13101_)
  );
  INV_X1 _47817_ (
    .A(_13101_),
    .ZN(_13102_)
  );
  AND2_X1 _47818_ (
    .A1(latched_branch),
    .A2(_12590_),
    .ZN(_13103_)
  );
  AND2_X1 _47819_ (
    .A1(_13102_),
    .A2(_13103_),
    .ZN(_13104_)
  );
  INV_X1 _47820_ (
    .A(_13104_),
    .ZN(_13105_)
  );
  AND2_X1 _47821_ (
    .A1(_13100_),
    .A2(_13105_),
    .ZN(_13106_)
  );
  INV_X1 _47822_ (
    .A(_13106_),
    .ZN(_13107_)
  );
  AND2_X1 _47823_ (
    .A1(_12555_),
    .A2(_13107_),
    .ZN(_13108_)
  );
  AND2_X1 _47824_ (
    .A1(_12755_),
    .A2(_13108_),
    .ZN(_13109_)
  );
  INV_X1 _47825_ (
    .A(_13109_),
    .ZN(_13110_)
  );
  AND2_X1 _47826_ (
    .A1(\cpuregs[23] [16]),
    .A2(_12756_),
    .ZN(_13111_)
  );
  INV_X1 _47827_ (
    .A(_13111_),
    .ZN(_13112_)
  );
  AND2_X1 _47828_ (
    .A1(_13110_),
    .A2(_13112_),
    .ZN(_13113_)
  );
  INV_X1 _47829_ (
    .A(_13113_),
    .ZN(_00543_)
  );
  AND2_X1 _47830_ (
    .A1(_03178_),
    .A2(_12542_),
    .ZN(_13114_)
  );
  INV_X1 _47831_ (
    .A(_13114_),
    .ZN(_13115_)
  );
  AND2_X1 _47832_ (
    .A1(_21087_),
    .A2(_12590_),
    .ZN(_13116_)
  );
  INV_X1 _47833_ (
    .A(_13116_),
    .ZN(_13117_)
  );
  AND2_X1 _47834_ (
    .A1(latched_branch),
    .A2(_12592_),
    .ZN(_13118_)
  );
  AND2_X1 _47835_ (
    .A1(_13117_),
    .A2(_13118_),
    .ZN(_13119_)
  );
  INV_X1 _47836_ (
    .A(_13119_),
    .ZN(_13120_)
  );
  AND2_X1 _47837_ (
    .A1(_13115_),
    .A2(_13120_),
    .ZN(_13121_)
  );
  INV_X1 _47838_ (
    .A(_13121_),
    .ZN(_13122_)
  );
  AND2_X1 _47839_ (
    .A1(_12555_),
    .A2(_13122_),
    .ZN(_13123_)
  );
  INV_X1 _47840_ (
    .A(_13123_),
    .ZN(_13124_)
  );
  AND2_X1 _47841_ (
    .A1(_12755_),
    .A2(_13123_),
    .ZN(_13125_)
  );
  INV_X1 _47842_ (
    .A(_13125_),
    .ZN(_13126_)
  );
  AND2_X1 _47843_ (
    .A1(\cpuregs[23] [17]),
    .A2(_12756_),
    .ZN(_13127_)
  );
  INV_X1 _47844_ (
    .A(_13127_),
    .ZN(_13128_)
  );
  AND2_X1 _47845_ (
    .A1(_13126_),
    .A2(_13128_),
    .ZN(_13129_)
  );
  INV_X1 _47846_ (
    .A(_13129_),
    .ZN(_00544_)
  );
  AND2_X1 _47847_ (
    .A1(_03194_),
    .A2(_12542_),
    .ZN(_13130_)
  );
  INV_X1 _47848_ (
    .A(_13130_),
    .ZN(_13131_)
  );
  AND2_X1 _47849_ (
    .A1(_21086_),
    .A2(_12592_),
    .ZN(_13132_)
  );
  INV_X1 _47850_ (
    .A(_13132_),
    .ZN(_13133_)
  );
  AND2_X1 _47851_ (
    .A1(latched_branch),
    .A2(_12594_),
    .ZN(_13134_)
  );
  AND2_X1 _47852_ (
    .A1(_13133_),
    .A2(_13134_),
    .ZN(_13135_)
  );
  INV_X1 _47853_ (
    .A(_13135_),
    .ZN(_13136_)
  );
  AND2_X1 _47854_ (
    .A1(_13131_),
    .A2(_13136_),
    .ZN(_13137_)
  );
  INV_X1 _47855_ (
    .A(_13137_),
    .ZN(_13138_)
  );
  AND2_X1 _47856_ (
    .A1(_12555_),
    .A2(_13138_),
    .ZN(_13139_)
  );
  AND2_X1 _47857_ (
    .A1(_12755_),
    .A2(_13139_),
    .ZN(_13140_)
  );
  INV_X1 _47858_ (
    .A(_13140_),
    .ZN(_13141_)
  );
  AND2_X1 _47859_ (
    .A1(\cpuregs[23] [18]),
    .A2(_12756_),
    .ZN(_13142_)
  );
  INV_X1 _47860_ (
    .A(_13142_),
    .ZN(_13143_)
  );
  AND2_X1 _47861_ (
    .A1(_13141_),
    .A2(_13143_),
    .ZN(_13144_)
  );
  INV_X1 _47862_ (
    .A(_13144_),
    .ZN(_00545_)
  );
  AND2_X1 _47863_ (
    .A1(_03210_),
    .A2(_12542_),
    .ZN(_13145_)
  );
  INV_X1 _47864_ (
    .A(_13145_),
    .ZN(_13146_)
  );
  AND2_X1 _47865_ (
    .A1(_21085_),
    .A2(_12594_),
    .ZN(_13147_)
  );
  INV_X1 _47866_ (
    .A(_13147_),
    .ZN(_13148_)
  );
  AND2_X1 _47867_ (
    .A1(latched_branch),
    .A2(_12596_),
    .ZN(_13149_)
  );
  AND2_X1 _47868_ (
    .A1(_13148_),
    .A2(_13149_),
    .ZN(_13150_)
  );
  INV_X1 _47869_ (
    .A(_13150_),
    .ZN(_13151_)
  );
  AND2_X1 _47870_ (
    .A1(_13146_),
    .A2(_13151_),
    .ZN(_13152_)
  );
  INV_X1 _47871_ (
    .A(_13152_),
    .ZN(_13153_)
  );
  AND2_X1 _47872_ (
    .A1(_12555_),
    .A2(_13153_),
    .ZN(_13154_)
  );
  AND2_X1 _47873_ (
    .A1(_12755_),
    .A2(_13154_),
    .ZN(_13155_)
  );
  INV_X1 _47874_ (
    .A(_13155_),
    .ZN(_13156_)
  );
  AND2_X1 _47875_ (
    .A1(\cpuregs[23] [19]),
    .A2(_12756_),
    .ZN(_13157_)
  );
  INV_X1 _47876_ (
    .A(_13157_),
    .ZN(_13158_)
  );
  AND2_X1 _47877_ (
    .A1(_13156_),
    .A2(_13158_),
    .ZN(_13159_)
  );
  INV_X1 _47878_ (
    .A(_13159_),
    .ZN(_00546_)
  );
  AND2_X1 _47879_ (
    .A1(_03226_),
    .A2(_12542_),
    .ZN(_13160_)
  );
  INV_X1 _47880_ (
    .A(_13160_),
    .ZN(_13161_)
  );
  AND2_X1 _47881_ (
    .A1(_21084_),
    .A2(_12596_),
    .ZN(_13162_)
  );
  INV_X1 _47882_ (
    .A(_13162_),
    .ZN(_13163_)
  );
  AND2_X1 _47883_ (
    .A1(latched_branch),
    .A2(_12598_),
    .ZN(_13164_)
  );
  AND2_X1 _47884_ (
    .A1(_13163_),
    .A2(_13164_),
    .ZN(_13165_)
  );
  INV_X1 _47885_ (
    .A(_13165_),
    .ZN(_13166_)
  );
  AND2_X1 _47886_ (
    .A1(_13161_),
    .A2(_13166_),
    .ZN(_13167_)
  );
  INV_X1 _47887_ (
    .A(_13167_),
    .ZN(_13168_)
  );
  AND2_X1 _47888_ (
    .A1(_12555_),
    .A2(_13168_),
    .ZN(_13169_)
  );
  AND2_X1 _47889_ (
    .A1(_12755_),
    .A2(_13169_),
    .ZN(_13170_)
  );
  INV_X1 _47890_ (
    .A(_13170_),
    .ZN(_13171_)
  );
  AND2_X1 _47891_ (
    .A1(\cpuregs[23] [20]),
    .A2(_12756_),
    .ZN(_13172_)
  );
  INV_X1 _47892_ (
    .A(_13172_),
    .ZN(_13173_)
  );
  AND2_X1 _47893_ (
    .A1(_13171_),
    .A2(_13173_),
    .ZN(_13174_)
  );
  INV_X1 _47894_ (
    .A(_13174_),
    .ZN(_00547_)
  );
  AND2_X1 _47895_ (
    .A1(_03242_),
    .A2(_12542_),
    .ZN(_13175_)
  );
  INV_X1 _47896_ (
    .A(_13175_),
    .ZN(_13176_)
  );
  AND2_X1 _47897_ (
    .A1(_21083_),
    .A2(_12598_),
    .ZN(_13177_)
  );
  INV_X1 _47898_ (
    .A(_13177_),
    .ZN(_13178_)
  );
  AND2_X1 _47899_ (
    .A1(latched_branch),
    .A2(_12600_),
    .ZN(_13179_)
  );
  AND2_X1 _47900_ (
    .A1(_13178_),
    .A2(_13179_),
    .ZN(_13180_)
  );
  INV_X1 _47901_ (
    .A(_13180_),
    .ZN(_13181_)
  );
  AND2_X1 _47902_ (
    .A1(_13176_),
    .A2(_13181_),
    .ZN(_13182_)
  );
  INV_X1 _47903_ (
    .A(_13182_),
    .ZN(_13183_)
  );
  AND2_X1 _47904_ (
    .A1(_12555_),
    .A2(_13183_),
    .ZN(_13184_)
  );
  AND2_X1 _47905_ (
    .A1(_12755_),
    .A2(_13184_),
    .ZN(_13185_)
  );
  INV_X1 _47906_ (
    .A(_13185_),
    .ZN(_13186_)
  );
  AND2_X1 _47907_ (
    .A1(\cpuregs[23] [21]),
    .A2(_12756_),
    .ZN(_13187_)
  );
  INV_X1 _47908_ (
    .A(_13187_),
    .ZN(_13188_)
  );
  AND2_X1 _47909_ (
    .A1(_13186_),
    .A2(_13188_),
    .ZN(_13189_)
  );
  INV_X1 _47910_ (
    .A(_13189_),
    .ZN(_00548_)
  );
  AND2_X1 _47911_ (
    .A1(_03258_),
    .A2(_12542_),
    .ZN(_13190_)
  );
  INV_X1 _47912_ (
    .A(_13190_),
    .ZN(_13191_)
  );
  AND2_X1 _47913_ (
    .A1(_21082_),
    .A2(_12600_),
    .ZN(_13192_)
  );
  INV_X1 _47914_ (
    .A(_13192_),
    .ZN(_13193_)
  );
  AND2_X1 _47915_ (
    .A1(latched_branch),
    .A2(_12602_),
    .ZN(_13194_)
  );
  AND2_X1 _47916_ (
    .A1(_13193_),
    .A2(_13194_),
    .ZN(_13195_)
  );
  INV_X1 _47917_ (
    .A(_13195_),
    .ZN(_13196_)
  );
  AND2_X1 _47918_ (
    .A1(_13191_),
    .A2(_13196_),
    .ZN(_13197_)
  );
  INV_X1 _47919_ (
    .A(_13197_),
    .ZN(_13198_)
  );
  AND2_X1 _47920_ (
    .A1(_12555_),
    .A2(_13198_),
    .ZN(_13199_)
  );
  AND2_X1 _47921_ (
    .A1(_12755_),
    .A2(_13199_),
    .ZN(_13200_)
  );
  INV_X1 _47922_ (
    .A(_13200_),
    .ZN(_13201_)
  );
  AND2_X1 _47923_ (
    .A1(\cpuregs[23] [22]),
    .A2(_12756_),
    .ZN(_13202_)
  );
  INV_X1 _47924_ (
    .A(_13202_),
    .ZN(_13203_)
  );
  AND2_X1 _47925_ (
    .A1(_13201_),
    .A2(_13203_),
    .ZN(_13204_)
  );
  INV_X1 _47926_ (
    .A(_13204_),
    .ZN(_00549_)
  );
  AND2_X1 _47927_ (
    .A1(_03274_),
    .A2(_12542_),
    .ZN(_13205_)
  );
  INV_X1 _47928_ (
    .A(_13205_),
    .ZN(_13206_)
  );
  AND2_X1 _47929_ (
    .A1(_21081_),
    .A2(_12602_),
    .ZN(_13207_)
  );
  INV_X1 _47930_ (
    .A(_13207_),
    .ZN(_13208_)
  );
  AND2_X1 _47931_ (
    .A1(latched_branch),
    .A2(_12604_),
    .ZN(_13209_)
  );
  AND2_X1 _47932_ (
    .A1(_13208_),
    .A2(_13209_),
    .ZN(_13210_)
  );
  INV_X1 _47933_ (
    .A(_13210_),
    .ZN(_13211_)
  );
  AND2_X1 _47934_ (
    .A1(_13206_),
    .A2(_13211_),
    .ZN(_13212_)
  );
  INV_X1 _47935_ (
    .A(_13212_),
    .ZN(_13213_)
  );
  AND2_X1 _47936_ (
    .A1(_12555_),
    .A2(_13213_),
    .ZN(_13214_)
  );
  AND2_X1 _47937_ (
    .A1(_12755_),
    .A2(_13214_),
    .ZN(_13215_)
  );
  INV_X1 _47938_ (
    .A(_13215_),
    .ZN(_13216_)
  );
  AND2_X1 _47939_ (
    .A1(\cpuregs[23] [23]),
    .A2(_12756_),
    .ZN(_13217_)
  );
  INV_X1 _47940_ (
    .A(_13217_),
    .ZN(_13218_)
  );
  AND2_X1 _47941_ (
    .A1(_13216_),
    .A2(_13218_),
    .ZN(_13219_)
  );
  INV_X1 _47942_ (
    .A(_13219_),
    .ZN(_00550_)
  );
  AND2_X1 _47943_ (
    .A1(_03290_),
    .A2(_12542_),
    .ZN(_13220_)
  );
  INV_X1 _47944_ (
    .A(_13220_),
    .ZN(_13221_)
  );
  AND2_X1 _47945_ (
    .A1(_21080_),
    .A2(_12604_),
    .ZN(_13222_)
  );
  INV_X1 _47946_ (
    .A(_13222_),
    .ZN(_13223_)
  );
  AND2_X1 _47947_ (
    .A1(latched_branch),
    .A2(_12606_),
    .ZN(_13224_)
  );
  AND2_X1 _47948_ (
    .A1(_13223_),
    .A2(_13224_),
    .ZN(_13225_)
  );
  INV_X1 _47949_ (
    .A(_13225_),
    .ZN(_13226_)
  );
  AND2_X1 _47950_ (
    .A1(_13221_),
    .A2(_13226_),
    .ZN(_13227_)
  );
  INV_X1 _47951_ (
    .A(_13227_),
    .ZN(_13228_)
  );
  AND2_X1 _47952_ (
    .A1(_12555_),
    .A2(_13228_),
    .ZN(_13229_)
  );
  AND2_X1 _47953_ (
    .A1(_12755_),
    .A2(_13229_),
    .ZN(_13230_)
  );
  INV_X1 _47954_ (
    .A(_13230_),
    .ZN(_13231_)
  );
  AND2_X1 _47955_ (
    .A1(\cpuregs[23] [24]),
    .A2(_12756_),
    .ZN(_13232_)
  );
  INV_X1 _47956_ (
    .A(_13232_),
    .ZN(_13233_)
  );
  AND2_X1 _47957_ (
    .A1(_13231_),
    .A2(_13233_),
    .ZN(_13234_)
  );
  INV_X1 _47958_ (
    .A(_13234_),
    .ZN(_00551_)
  );
  AND2_X1 _47959_ (
    .A1(_03306_),
    .A2(_12542_),
    .ZN(_13235_)
  );
  INV_X1 _47960_ (
    .A(_13235_),
    .ZN(_13236_)
  );
  AND2_X1 _47961_ (
    .A1(_21079_),
    .A2(_12606_),
    .ZN(_13237_)
  );
  INV_X1 _47962_ (
    .A(_13237_),
    .ZN(_13238_)
  );
  AND2_X1 _47963_ (
    .A1(latched_branch),
    .A2(_12608_),
    .ZN(_13239_)
  );
  AND2_X1 _47964_ (
    .A1(_13238_),
    .A2(_13239_),
    .ZN(_13240_)
  );
  INV_X1 _47965_ (
    .A(_13240_),
    .ZN(_13241_)
  );
  AND2_X1 _47966_ (
    .A1(_13236_),
    .A2(_13241_),
    .ZN(_13242_)
  );
  INV_X1 _47967_ (
    .A(_13242_),
    .ZN(_13243_)
  );
  AND2_X1 _47968_ (
    .A1(_12555_),
    .A2(_13243_),
    .ZN(_13244_)
  );
  AND2_X1 _47969_ (
    .A1(_12755_),
    .A2(_13244_),
    .ZN(_13245_)
  );
  INV_X1 _47970_ (
    .A(_13245_),
    .ZN(_13246_)
  );
  AND2_X1 _47971_ (
    .A1(\cpuregs[23] [25]),
    .A2(_12756_),
    .ZN(_13247_)
  );
  INV_X1 _47972_ (
    .A(_13247_),
    .ZN(_13248_)
  );
  AND2_X1 _47973_ (
    .A1(_13246_),
    .A2(_13248_),
    .ZN(_13249_)
  );
  INV_X1 _47974_ (
    .A(_13249_),
    .ZN(_00552_)
  );
  AND2_X1 _47975_ (
    .A1(_03322_),
    .A2(_12542_),
    .ZN(_13250_)
  );
  INV_X1 _47976_ (
    .A(_13250_),
    .ZN(_13251_)
  );
  AND2_X1 _47977_ (
    .A1(_21078_),
    .A2(_12608_),
    .ZN(_13252_)
  );
  INV_X1 _47978_ (
    .A(_13252_),
    .ZN(_13253_)
  );
  AND2_X1 _47979_ (
    .A1(latched_branch),
    .A2(_12610_),
    .ZN(_13254_)
  );
  AND2_X1 _47980_ (
    .A1(_13253_),
    .A2(_13254_),
    .ZN(_13255_)
  );
  INV_X1 _47981_ (
    .A(_13255_),
    .ZN(_13256_)
  );
  AND2_X1 _47982_ (
    .A1(_13251_),
    .A2(_13256_),
    .ZN(_13257_)
  );
  INV_X1 _47983_ (
    .A(_13257_),
    .ZN(_13258_)
  );
  AND2_X1 _47984_ (
    .A1(_12555_),
    .A2(_13258_),
    .ZN(_13259_)
  );
  AND2_X1 _47985_ (
    .A1(_12755_),
    .A2(_13259_),
    .ZN(_13260_)
  );
  INV_X1 _47986_ (
    .A(_13260_),
    .ZN(_13261_)
  );
  AND2_X1 _47987_ (
    .A1(\cpuregs[23] [26]),
    .A2(_12756_),
    .ZN(_13262_)
  );
  INV_X1 _47988_ (
    .A(_13262_),
    .ZN(_13263_)
  );
  AND2_X1 _47989_ (
    .A1(_13261_),
    .A2(_13263_),
    .ZN(_13264_)
  );
  INV_X1 _47990_ (
    .A(_13264_),
    .ZN(_00553_)
  );
  AND2_X1 _47991_ (
    .A1(_03338_),
    .A2(_12542_),
    .ZN(_13265_)
  );
  INV_X1 _47992_ (
    .A(_13265_),
    .ZN(_13266_)
  );
  AND2_X1 _47993_ (
    .A1(_21077_),
    .A2(_12610_),
    .ZN(_13267_)
  );
  INV_X1 _47994_ (
    .A(_13267_),
    .ZN(_13268_)
  );
  AND2_X1 _47995_ (
    .A1(latched_branch),
    .A2(_12612_),
    .ZN(_13269_)
  );
  AND2_X1 _47996_ (
    .A1(_13268_),
    .A2(_13269_),
    .ZN(_13270_)
  );
  INV_X1 _47997_ (
    .A(_13270_),
    .ZN(_13271_)
  );
  AND2_X1 _47998_ (
    .A1(_13266_),
    .A2(_13271_),
    .ZN(_13272_)
  );
  INV_X1 _47999_ (
    .A(_13272_),
    .ZN(_13273_)
  );
  AND2_X1 _48000_ (
    .A1(_12555_),
    .A2(_13273_),
    .ZN(_13274_)
  );
  AND2_X1 _48001_ (
    .A1(_12755_),
    .A2(_13274_),
    .ZN(_13275_)
  );
  INV_X1 _48002_ (
    .A(_13275_),
    .ZN(_13276_)
  );
  AND2_X1 _48003_ (
    .A1(\cpuregs[23] [27]),
    .A2(_12756_),
    .ZN(_13277_)
  );
  INV_X1 _48004_ (
    .A(_13277_),
    .ZN(_13278_)
  );
  AND2_X1 _48005_ (
    .A1(_13276_),
    .A2(_13278_),
    .ZN(_13279_)
  );
  INV_X1 _48006_ (
    .A(_13279_),
    .ZN(_00554_)
  );
  AND2_X1 _48007_ (
    .A1(_03354_),
    .A2(_12542_),
    .ZN(_13280_)
  );
  INV_X1 _48008_ (
    .A(_13280_),
    .ZN(_13281_)
  );
  AND2_X1 _48009_ (
    .A1(_21076_),
    .A2(_12612_),
    .ZN(_13282_)
  );
  INV_X1 _48010_ (
    .A(_13282_),
    .ZN(_13283_)
  );
  AND2_X1 _48011_ (
    .A1(latched_branch),
    .A2(_12614_),
    .ZN(_13284_)
  );
  AND2_X1 _48012_ (
    .A1(_13283_),
    .A2(_13284_),
    .ZN(_13285_)
  );
  INV_X1 _48013_ (
    .A(_13285_),
    .ZN(_13286_)
  );
  AND2_X1 _48014_ (
    .A1(_13281_),
    .A2(_13286_),
    .ZN(_13287_)
  );
  INV_X1 _48015_ (
    .A(_13287_),
    .ZN(_13288_)
  );
  AND2_X1 _48016_ (
    .A1(_12555_),
    .A2(_13288_),
    .ZN(_13289_)
  );
  AND2_X1 _48017_ (
    .A1(_12755_),
    .A2(_13289_),
    .ZN(_13290_)
  );
  INV_X1 _48018_ (
    .A(_13290_),
    .ZN(_13291_)
  );
  AND2_X1 _48019_ (
    .A1(\cpuregs[23] [28]),
    .A2(_12756_),
    .ZN(_13292_)
  );
  INV_X1 _48020_ (
    .A(_13292_),
    .ZN(_13293_)
  );
  AND2_X1 _48021_ (
    .A1(_13291_),
    .A2(_13293_),
    .ZN(_13294_)
  );
  INV_X1 _48022_ (
    .A(_13294_),
    .ZN(_00555_)
  );
  AND2_X1 _48023_ (
    .A1(_03370_),
    .A2(_12542_),
    .ZN(_13295_)
  );
  INV_X1 _48024_ (
    .A(_13295_),
    .ZN(_13296_)
  );
  AND2_X1 _48025_ (
    .A1(_21075_),
    .A2(_12614_),
    .ZN(_13297_)
  );
  INV_X1 _48026_ (
    .A(_13297_),
    .ZN(_13298_)
  );
  AND2_X1 _48027_ (
    .A1(latched_branch),
    .A2(_12616_),
    .ZN(_13299_)
  );
  AND2_X1 _48028_ (
    .A1(_13298_),
    .A2(_13299_),
    .ZN(_13300_)
  );
  INV_X1 _48029_ (
    .A(_13300_),
    .ZN(_13301_)
  );
  AND2_X1 _48030_ (
    .A1(_13296_),
    .A2(_13301_),
    .ZN(_13302_)
  );
  INV_X1 _48031_ (
    .A(_13302_),
    .ZN(_13303_)
  );
  AND2_X1 _48032_ (
    .A1(_12555_),
    .A2(_13303_),
    .ZN(_13304_)
  );
  AND2_X1 _48033_ (
    .A1(_12755_),
    .A2(_13304_),
    .ZN(_13305_)
  );
  INV_X1 _48034_ (
    .A(_13305_),
    .ZN(_13306_)
  );
  AND2_X1 _48035_ (
    .A1(\cpuregs[23] [29]),
    .A2(_12756_),
    .ZN(_13307_)
  );
  INV_X1 _48036_ (
    .A(_13307_),
    .ZN(_13308_)
  );
  AND2_X1 _48037_ (
    .A1(_13306_),
    .A2(_13308_),
    .ZN(_13309_)
  );
  INV_X1 _48038_ (
    .A(_13309_),
    .ZN(_00556_)
  );
  AND2_X1 _48039_ (
    .A1(_03386_),
    .A2(_12542_),
    .ZN(_13310_)
  );
  INV_X1 _48040_ (
    .A(_13310_),
    .ZN(_13311_)
  );
  AND2_X1 _48041_ (
    .A1(_21074_),
    .A2(_12616_),
    .ZN(_13312_)
  );
  INV_X1 _48042_ (
    .A(_13312_),
    .ZN(_13313_)
  );
  AND2_X1 _48043_ (
    .A1(latched_branch),
    .A2(_12618_),
    .ZN(_13314_)
  );
  AND2_X1 _48044_ (
    .A1(_13313_),
    .A2(_13314_),
    .ZN(_13315_)
  );
  INV_X1 _48045_ (
    .A(_13315_),
    .ZN(_13316_)
  );
  AND2_X1 _48046_ (
    .A1(_13311_),
    .A2(_13316_),
    .ZN(_13317_)
  );
  INV_X1 _48047_ (
    .A(_13317_),
    .ZN(_13318_)
  );
  AND2_X1 _48048_ (
    .A1(_12555_),
    .A2(_13318_),
    .ZN(_13319_)
  );
  AND2_X1 _48049_ (
    .A1(_12755_),
    .A2(_13319_),
    .ZN(_13320_)
  );
  INV_X1 _48050_ (
    .A(_13320_),
    .ZN(_13321_)
  );
  AND2_X1 _48051_ (
    .A1(\cpuregs[23] [30]),
    .A2(_12756_),
    .ZN(_13322_)
  );
  INV_X1 _48052_ (
    .A(_13322_),
    .ZN(_13323_)
  );
  AND2_X1 _48053_ (
    .A1(_13321_),
    .A2(_13323_),
    .ZN(_13324_)
  );
  INV_X1 _48054_ (
    .A(_13324_),
    .ZN(_00557_)
  );
  AND2_X1 _48055_ (
    .A1(_12828_),
    .A2(_12874_),
    .ZN(_13325_)
  );
  INV_X1 _48056_ (
    .A(_13325_),
    .ZN(_13326_)
  );
  AND2_X1 _48057_ (
    .A1(\cpuregs[14] [0]),
    .A2(_12829_),
    .ZN(_13327_)
  );
  INV_X1 _48058_ (
    .A(_13327_),
    .ZN(_13328_)
  );
  AND2_X1 _48059_ (
    .A1(_13326_),
    .A2(_13328_),
    .ZN(_13329_)
  );
  INV_X1 _48060_ (
    .A(_13329_),
    .ZN(_00558_)
  );
  AND2_X1 _48061_ (
    .A1(_12828_),
    .A2(_12886_),
    .ZN(_13330_)
  );
  INV_X1 _48062_ (
    .A(_13330_),
    .ZN(_13331_)
  );
  AND2_X1 _48063_ (
    .A1(\cpuregs[14] [1]),
    .A2(_12829_),
    .ZN(_13332_)
  );
  INV_X1 _48064_ (
    .A(_13332_),
    .ZN(_13333_)
  );
  AND2_X1 _48065_ (
    .A1(_13331_),
    .A2(_13333_),
    .ZN(_13334_)
  );
  INV_X1 _48066_ (
    .A(_13334_),
    .ZN(_00559_)
  );
  AND2_X1 _48067_ (
    .A1(_12828_),
    .A2(_12900_),
    .ZN(_13335_)
  );
  INV_X1 _48068_ (
    .A(_13335_),
    .ZN(_13336_)
  );
  AND2_X1 _48069_ (
    .A1(\cpuregs[14] [2]),
    .A2(_12829_),
    .ZN(_13337_)
  );
  INV_X1 _48070_ (
    .A(_13337_),
    .ZN(_13338_)
  );
  AND2_X1 _48071_ (
    .A1(_13336_),
    .A2(_13338_),
    .ZN(_13339_)
  );
  INV_X1 _48072_ (
    .A(_13339_),
    .ZN(_00560_)
  );
  AND2_X1 _48073_ (
    .A1(_12828_),
    .A2(_12913_),
    .ZN(_13340_)
  );
  INV_X1 _48074_ (
    .A(_13340_),
    .ZN(_13341_)
  );
  AND2_X1 _48075_ (
    .A1(\cpuregs[14] [3]),
    .A2(_12829_),
    .ZN(_13342_)
  );
  INV_X1 _48076_ (
    .A(_13342_),
    .ZN(_13343_)
  );
  AND2_X1 _48077_ (
    .A1(_13341_),
    .A2(_13343_),
    .ZN(_13344_)
  );
  INV_X1 _48078_ (
    .A(_13344_),
    .ZN(_00561_)
  );
  AND2_X1 _48079_ (
    .A1(_12828_),
    .A2(_12928_),
    .ZN(_13345_)
  );
  INV_X1 _48080_ (
    .A(_13345_),
    .ZN(_13346_)
  );
  AND2_X1 _48081_ (
    .A1(\cpuregs[14] [4]),
    .A2(_12829_),
    .ZN(_13347_)
  );
  INV_X1 _48082_ (
    .A(_13347_),
    .ZN(_13348_)
  );
  AND2_X1 _48083_ (
    .A1(_13346_),
    .A2(_13348_),
    .ZN(_13349_)
  );
  INV_X1 _48084_ (
    .A(_13349_),
    .ZN(_00562_)
  );
  AND2_X1 _48085_ (
    .A1(_12828_),
    .A2(_12943_),
    .ZN(_13350_)
  );
  INV_X1 _48086_ (
    .A(_13350_),
    .ZN(_13351_)
  );
  AND2_X1 _48087_ (
    .A1(\cpuregs[14] [5]),
    .A2(_12829_),
    .ZN(_13352_)
  );
  INV_X1 _48088_ (
    .A(_13352_),
    .ZN(_13353_)
  );
  AND2_X1 _48089_ (
    .A1(_13351_),
    .A2(_13353_),
    .ZN(_13354_)
  );
  INV_X1 _48090_ (
    .A(_13354_),
    .ZN(_00563_)
  );
  AND2_X1 _48091_ (
    .A1(_12828_),
    .A2(_12958_),
    .ZN(_13355_)
  );
  INV_X1 _48092_ (
    .A(_13355_),
    .ZN(_13356_)
  );
  AND2_X1 _48093_ (
    .A1(\cpuregs[14] [6]),
    .A2(_12829_),
    .ZN(_13357_)
  );
  INV_X1 _48094_ (
    .A(_13357_),
    .ZN(_13358_)
  );
  AND2_X1 _48095_ (
    .A1(_13356_),
    .A2(_13358_),
    .ZN(_13359_)
  );
  INV_X1 _48096_ (
    .A(_13359_),
    .ZN(_00564_)
  );
  AND2_X1 _48097_ (
    .A1(_12828_),
    .A2(_12973_),
    .ZN(_13360_)
  );
  INV_X1 _48098_ (
    .A(_13360_),
    .ZN(_13361_)
  );
  AND2_X1 _48099_ (
    .A1(\cpuregs[14] [7]),
    .A2(_12829_),
    .ZN(_13362_)
  );
  INV_X1 _48100_ (
    .A(_13362_),
    .ZN(_13363_)
  );
  AND2_X1 _48101_ (
    .A1(_13361_),
    .A2(_13363_),
    .ZN(_13364_)
  );
  INV_X1 _48102_ (
    .A(_13364_),
    .ZN(_00565_)
  );
  AND2_X1 _48103_ (
    .A1(_12828_),
    .A2(_12988_),
    .ZN(_13365_)
  );
  INV_X1 _48104_ (
    .A(_13365_),
    .ZN(_13366_)
  );
  AND2_X1 _48105_ (
    .A1(\cpuregs[14] [8]),
    .A2(_12829_),
    .ZN(_13367_)
  );
  INV_X1 _48106_ (
    .A(_13367_),
    .ZN(_13368_)
  );
  AND2_X1 _48107_ (
    .A1(_13366_),
    .A2(_13368_),
    .ZN(_13369_)
  );
  INV_X1 _48108_ (
    .A(_13369_),
    .ZN(_00566_)
  );
  AND2_X1 _48109_ (
    .A1(_12828_),
    .A2(_13003_),
    .ZN(_13370_)
  );
  INV_X1 _48110_ (
    .A(_13370_),
    .ZN(_13371_)
  );
  AND2_X1 _48111_ (
    .A1(\cpuregs[14] [9]),
    .A2(_12829_),
    .ZN(_13372_)
  );
  INV_X1 _48112_ (
    .A(_13372_),
    .ZN(_13373_)
  );
  AND2_X1 _48113_ (
    .A1(_13371_),
    .A2(_13373_),
    .ZN(_13374_)
  );
  INV_X1 _48114_ (
    .A(_13374_),
    .ZN(_00567_)
  );
  AND2_X1 _48115_ (
    .A1(_12828_),
    .A2(_13018_),
    .ZN(_13375_)
  );
  INV_X1 _48116_ (
    .A(_13375_),
    .ZN(_13376_)
  );
  AND2_X1 _48117_ (
    .A1(\cpuregs[14] [10]),
    .A2(_12829_),
    .ZN(_13377_)
  );
  INV_X1 _48118_ (
    .A(_13377_),
    .ZN(_13378_)
  );
  AND2_X1 _48119_ (
    .A1(_13376_),
    .A2(_13378_),
    .ZN(_13379_)
  );
  INV_X1 _48120_ (
    .A(_13379_),
    .ZN(_00568_)
  );
  AND2_X1 _48121_ (
    .A1(_12828_),
    .A2(_13033_),
    .ZN(_13380_)
  );
  INV_X1 _48122_ (
    .A(_13380_),
    .ZN(_13381_)
  );
  AND2_X1 _48123_ (
    .A1(\cpuregs[14] [11]),
    .A2(_12829_),
    .ZN(_13382_)
  );
  INV_X1 _48124_ (
    .A(_13382_),
    .ZN(_13383_)
  );
  AND2_X1 _48125_ (
    .A1(_13381_),
    .A2(_13383_),
    .ZN(_13384_)
  );
  INV_X1 _48126_ (
    .A(_13384_),
    .ZN(_00569_)
  );
  AND2_X1 _48127_ (
    .A1(_12828_),
    .A2(_13048_),
    .ZN(_13385_)
  );
  INV_X1 _48128_ (
    .A(_13385_),
    .ZN(_13386_)
  );
  AND2_X1 _48129_ (
    .A1(\cpuregs[14] [12]),
    .A2(_12829_),
    .ZN(_13387_)
  );
  INV_X1 _48130_ (
    .A(_13387_),
    .ZN(_13388_)
  );
  AND2_X1 _48131_ (
    .A1(_13386_),
    .A2(_13388_),
    .ZN(_13389_)
  );
  INV_X1 _48132_ (
    .A(_13389_),
    .ZN(_00570_)
  );
  AND2_X1 _48133_ (
    .A1(_12828_),
    .A2(_13063_),
    .ZN(_13390_)
  );
  INV_X1 _48134_ (
    .A(_13390_),
    .ZN(_13391_)
  );
  AND2_X1 _48135_ (
    .A1(\cpuregs[14] [13]),
    .A2(_12829_),
    .ZN(_13392_)
  );
  INV_X1 _48136_ (
    .A(_13392_),
    .ZN(_13393_)
  );
  AND2_X1 _48137_ (
    .A1(_13391_),
    .A2(_13393_),
    .ZN(_13394_)
  );
  INV_X1 _48138_ (
    .A(_13394_),
    .ZN(_00571_)
  );
  AND2_X1 _48139_ (
    .A1(\cpuregs[14] [14]),
    .A2(_12829_),
    .ZN(_13395_)
  );
  INV_X1 _48140_ (
    .A(_13395_),
    .ZN(_13396_)
  );
  AND2_X1 _48141_ (
    .A1(_12828_),
    .A2(_13078_),
    .ZN(_13397_)
  );
  INV_X1 _48142_ (
    .A(_13397_),
    .ZN(_13398_)
  );
  AND2_X1 _48143_ (
    .A1(_13396_),
    .A2(_13398_),
    .ZN(_13399_)
  );
  INV_X1 _48144_ (
    .A(_13399_),
    .ZN(_00572_)
  );
  AND2_X1 _48145_ (
    .A1(_12828_),
    .A2(_13093_),
    .ZN(_13400_)
  );
  INV_X1 _48146_ (
    .A(_13400_),
    .ZN(_13401_)
  );
  AND2_X1 _48147_ (
    .A1(\cpuregs[14] [15]),
    .A2(_12829_),
    .ZN(_13402_)
  );
  INV_X1 _48148_ (
    .A(_13402_),
    .ZN(_13403_)
  );
  AND2_X1 _48149_ (
    .A1(_13401_),
    .A2(_13403_),
    .ZN(_13404_)
  );
  INV_X1 _48150_ (
    .A(_13404_),
    .ZN(_00573_)
  );
  AND2_X1 _48151_ (
    .A1(_12828_),
    .A2(_13108_),
    .ZN(_13405_)
  );
  INV_X1 _48152_ (
    .A(_13405_),
    .ZN(_13406_)
  );
  AND2_X1 _48153_ (
    .A1(\cpuregs[14] [16]),
    .A2(_12829_),
    .ZN(_13407_)
  );
  INV_X1 _48154_ (
    .A(_13407_),
    .ZN(_13408_)
  );
  AND2_X1 _48155_ (
    .A1(_13406_),
    .A2(_13408_),
    .ZN(_13409_)
  );
  INV_X1 _48156_ (
    .A(_13409_),
    .ZN(_00574_)
  );
  AND2_X1 _48157_ (
    .A1(\cpuregs[14] [17]),
    .A2(_12829_),
    .ZN(_13410_)
  );
  INV_X1 _48158_ (
    .A(_13410_),
    .ZN(_13411_)
  );
  AND2_X1 _48159_ (
    .A1(_12828_),
    .A2(_13123_),
    .ZN(_13412_)
  );
  INV_X1 _48160_ (
    .A(_13412_),
    .ZN(_13413_)
  );
  AND2_X1 _48161_ (
    .A1(_13411_),
    .A2(_13413_),
    .ZN(_13414_)
  );
  INV_X1 _48162_ (
    .A(_13414_),
    .ZN(_00575_)
  );
  AND2_X1 _48163_ (
    .A1(\cpuregs[14] [18]),
    .A2(_12829_),
    .ZN(_13415_)
  );
  INV_X1 _48164_ (
    .A(_13415_),
    .ZN(_13416_)
  );
  AND2_X1 _48165_ (
    .A1(_12828_),
    .A2(_13139_),
    .ZN(_13417_)
  );
  INV_X1 _48166_ (
    .A(_13417_),
    .ZN(_13418_)
  );
  AND2_X1 _48167_ (
    .A1(_13416_),
    .A2(_13418_),
    .ZN(_13419_)
  );
  INV_X1 _48168_ (
    .A(_13419_),
    .ZN(_00576_)
  );
  AND2_X1 _48169_ (
    .A1(\cpuregs[14] [19]),
    .A2(_12829_),
    .ZN(_13420_)
  );
  INV_X1 _48170_ (
    .A(_13420_),
    .ZN(_13421_)
  );
  AND2_X1 _48171_ (
    .A1(_12828_),
    .A2(_13154_),
    .ZN(_13422_)
  );
  INV_X1 _48172_ (
    .A(_13422_),
    .ZN(_13423_)
  );
  AND2_X1 _48173_ (
    .A1(_13421_),
    .A2(_13423_),
    .ZN(_13424_)
  );
  INV_X1 _48174_ (
    .A(_13424_),
    .ZN(_00577_)
  );
  AND2_X1 _48175_ (
    .A1(\cpuregs[14] [20]),
    .A2(_12829_),
    .ZN(_13425_)
  );
  INV_X1 _48176_ (
    .A(_13425_),
    .ZN(_13426_)
  );
  AND2_X1 _48177_ (
    .A1(_12828_),
    .A2(_13169_),
    .ZN(_13427_)
  );
  INV_X1 _48178_ (
    .A(_13427_),
    .ZN(_13428_)
  );
  AND2_X1 _48179_ (
    .A1(_13426_),
    .A2(_13428_),
    .ZN(_13429_)
  );
  INV_X1 _48180_ (
    .A(_13429_),
    .ZN(_00578_)
  );
  AND2_X1 _48181_ (
    .A1(\cpuregs[14] [21]),
    .A2(_12829_),
    .ZN(_13430_)
  );
  INV_X1 _48182_ (
    .A(_13430_),
    .ZN(_13431_)
  );
  AND2_X1 _48183_ (
    .A1(_12828_),
    .A2(_13184_),
    .ZN(_13432_)
  );
  INV_X1 _48184_ (
    .A(_13432_),
    .ZN(_13433_)
  );
  AND2_X1 _48185_ (
    .A1(_13431_),
    .A2(_13433_),
    .ZN(_13434_)
  );
  INV_X1 _48186_ (
    .A(_13434_),
    .ZN(_00579_)
  );
  AND2_X1 _48187_ (
    .A1(\cpuregs[14] [22]),
    .A2(_12829_),
    .ZN(_13435_)
  );
  INV_X1 _48188_ (
    .A(_13435_),
    .ZN(_13436_)
  );
  AND2_X1 _48189_ (
    .A1(_12828_),
    .A2(_13199_),
    .ZN(_13437_)
  );
  INV_X1 _48190_ (
    .A(_13437_),
    .ZN(_13438_)
  );
  AND2_X1 _48191_ (
    .A1(_13436_),
    .A2(_13438_),
    .ZN(_13439_)
  );
  INV_X1 _48192_ (
    .A(_13439_),
    .ZN(_00580_)
  );
  AND2_X1 _48193_ (
    .A1(\cpuregs[14] [23]),
    .A2(_12829_),
    .ZN(_13440_)
  );
  INV_X1 _48194_ (
    .A(_13440_),
    .ZN(_13441_)
  );
  AND2_X1 _48195_ (
    .A1(_12828_),
    .A2(_13214_),
    .ZN(_13442_)
  );
  INV_X1 _48196_ (
    .A(_13442_),
    .ZN(_13443_)
  );
  AND2_X1 _48197_ (
    .A1(_13441_),
    .A2(_13443_),
    .ZN(_13444_)
  );
  INV_X1 _48198_ (
    .A(_13444_),
    .ZN(_00581_)
  );
  AND2_X1 _48199_ (
    .A1(\cpuregs[14] [24]),
    .A2(_12829_),
    .ZN(_13445_)
  );
  INV_X1 _48200_ (
    .A(_13445_),
    .ZN(_13446_)
  );
  AND2_X1 _48201_ (
    .A1(_12828_),
    .A2(_13229_),
    .ZN(_13447_)
  );
  INV_X1 _48202_ (
    .A(_13447_),
    .ZN(_13448_)
  );
  AND2_X1 _48203_ (
    .A1(_13446_),
    .A2(_13448_),
    .ZN(_13449_)
  );
  INV_X1 _48204_ (
    .A(_13449_),
    .ZN(_00582_)
  );
  AND2_X1 _48205_ (
    .A1(\cpuregs[14] [25]),
    .A2(_12829_),
    .ZN(_13450_)
  );
  INV_X1 _48206_ (
    .A(_13450_),
    .ZN(_13451_)
  );
  AND2_X1 _48207_ (
    .A1(_12828_),
    .A2(_13244_),
    .ZN(_13452_)
  );
  INV_X1 _48208_ (
    .A(_13452_),
    .ZN(_13453_)
  );
  AND2_X1 _48209_ (
    .A1(_13451_),
    .A2(_13453_),
    .ZN(_13454_)
  );
  INV_X1 _48210_ (
    .A(_13454_),
    .ZN(_00583_)
  );
  AND2_X1 _48211_ (
    .A1(\cpuregs[14] [26]),
    .A2(_12829_),
    .ZN(_13455_)
  );
  INV_X1 _48212_ (
    .A(_13455_),
    .ZN(_13456_)
  );
  AND2_X1 _48213_ (
    .A1(_12828_),
    .A2(_13259_),
    .ZN(_13457_)
  );
  INV_X1 _48214_ (
    .A(_13457_),
    .ZN(_13458_)
  );
  AND2_X1 _48215_ (
    .A1(_13456_),
    .A2(_13458_),
    .ZN(_13459_)
  );
  INV_X1 _48216_ (
    .A(_13459_),
    .ZN(_00584_)
  );
  AND2_X1 _48217_ (
    .A1(\cpuregs[14] [27]),
    .A2(_12829_),
    .ZN(_13460_)
  );
  INV_X1 _48218_ (
    .A(_13460_),
    .ZN(_13461_)
  );
  AND2_X1 _48219_ (
    .A1(_12828_),
    .A2(_13274_),
    .ZN(_13462_)
  );
  INV_X1 _48220_ (
    .A(_13462_),
    .ZN(_13463_)
  );
  AND2_X1 _48221_ (
    .A1(_13461_),
    .A2(_13463_),
    .ZN(_13464_)
  );
  INV_X1 _48222_ (
    .A(_13464_),
    .ZN(_00585_)
  );
  AND2_X1 _48223_ (
    .A1(\cpuregs[14] [28]),
    .A2(_12829_),
    .ZN(_13465_)
  );
  INV_X1 _48224_ (
    .A(_13465_),
    .ZN(_13466_)
  );
  AND2_X1 _48225_ (
    .A1(_12828_),
    .A2(_13289_),
    .ZN(_13467_)
  );
  INV_X1 _48226_ (
    .A(_13467_),
    .ZN(_13468_)
  );
  AND2_X1 _48227_ (
    .A1(_13466_),
    .A2(_13468_),
    .ZN(_13469_)
  );
  INV_X1 _48228_ (
    .A(_13469_),
    .ZN(_00586_)
  );
  AND2_X1 _48229_ (
    .A1(\cpuregs[14] [29]),
    .A2(_12829_),
    .ZN(_13470_)
  );
  INV_X1 _48230_ (
    .A(_13470_),
    .ZN(_13471_)
  );
  AND2_X1 _48231_ (
    .A1(_12828_),
    .A2(_13304_),
    .ZN(_13472_)
  );
  INV_X1 _48232_ (
    .A(_13472_),
    .ZN(_13473_)
  );
  AND2_X1 _48233_ (
    .A1(_13471_),
    .A2(_13473_),
    .ZN(_13474_)
  );
  INV_X1 _48234_ (
    .A(_13474_),
    .ZN(_00587_)
  );
  AND2_X1 _48235_ (
    .A1(\cpuregs[14] [30]),
    .A2(_12829_),
    .ZN(_13475_)
  );
  INV_X1 _48236_ (
    .A(_13475_),
    .ZN(_13476_)
  );
  AND2_X1 _48237_ (
    .A1(_12828_),
    .A2(_13319_),
    .ZN(_13477_)
  );
  INV_X1 _48238_ (
    .A(_13477_),
    .ZN(_13478_)
  );
  AND2_X1 _48239_ (
    .A1(_13476_),
    .A2(_13478_),
    .ZN(_13479_)
  );
  INV_X1 _48240_ (
    .A(_13479_),
    .ZN(_00588_)
  );
  AND2_X1 _48241_ (
    .A1(_12821_),
    .A2(_12874_),
    .ZN(_13480_)
  );
  INV_X1 _48242_ (
    .A(_13480_),
    .ZN(_13481_)
  );
  AND2_X1 _48243_ (
    .A1(\cpuregs[15] [0]),
    .A2(_12822_),
    .ZN(_13482_)
  );
  INV_X1 _48244_ (
    .A(_13482_),
    .ZN(_13483_)
  );
  AND2_X1 _48245_ (
    .A1(_13481_),
    .A2(_13483_),
    .ZN(_13484_)
  );
  INV_X1 _48246_ (
    .A(_13484_),
    .ZN(_00589_)
  );
  AND2_X1 _48247_ (
    .A1(_12821_),
    .A2(_12886_),
    .ZN(_13485_)
  );
  INV_X1 _48248_ (
    .A(_13485_),
    .ZN(_13486_)
  );
  AND2_X1 _48249_ (
    .A1(\cpuregs[15] [1]),
    .A2(_12822_),
    .ZN(_13487_)
  );
  INV_X1 _48250_ (
    .A(_13487_),
    .ZN(_13488_)
  );
  AND2_X1 _48251_ (
    .A1(_13486_),
    .A2(_13488_),
    .ZN(_13489_)
  );
  INV_X1 _48252_ (
    .A(_13489_),
    .ZN(_00590_)
  );
  AND2_X1 _48253_ (
    .A1(_12821_),
    .A2(_12900_),
    .ZN(_13490_)
  );
  INV_X1 _48254_ (
    .A(_13490_),
    .ZN(_13491_)
  );
  AND2_X1 _48255_ (
    .A1(\cpuregs[15] [2]),
    .A2(_12822_),
    .ZN(_13492_)
  );
  INV_X1 _48256_ (
    .A(_13492_),
    .ZN(_13493_)
  );
  AND2_X1 _48257_ (
    .A1(_13491_),
    .A2(_13493_),
    .ZN(_13494_)
  );
  INV_X1 _48258_ (
    .A(_13494_),
    .ZN(_00591_)
  );
  AND2_X1 _48259_ (
    .A1(_12821_),
    .A2(_12913_),
    .ZN(_13495_)
  );
  INV_X1 _48260_ (
    .A(_13495_),
    .ZN(_13496_)
  );
  AND2_X1 _48261_ (
    .A1(\cpuregs[15] [3]),
    .A2(_12822_),
    .ZN(_13497_)
  );
  INV_X1 _48262_ (
    .A(_13497_),
    .ZN(_13498_)
  );
  AND2_X1 _48263_ (
    .A1(_13496_),
    .A2(_13498_),
    .ZN(_13499_)
  );
  INV_X1 _48264_ (
    .A(_13499_),
    .ZN(_00592_)
  );
  AND2_X1 _48265_ (
    .A1(_12821_),
    .A2(_12928_),
    .ZN(_13500_)
  );
  INV_X1 _48266_ (
    .A(_13500_),
    .ZN(_13501_)
  );
  AND2_X1 _48267_ (
    .A1(\cpuregs[15] [4]),
    .A2(_12822_),
    .ZN(_13502_)
  );
  INV_X1 _48268_ (
    .A(_13502_),
    .ZN(_13503_)
  );
  AND2_X1 _48269_ (
    .A1(_13501_),
    .A2(_13503_),
    .ZN(_13504_)
  );
  INV_X1 _48270_ (
    .A(_13504_),
    .ZN(_00593_)
  );
  AND2_X1 _48271_ (
    .A1(_12821_),
    .A2(_12943_),
    .ZN(_13505_)
  );
  INV_X1 _48272_ (
    .A(_13505_),
    .ZN(_13506_)
  );
  AND2_X1 _48273_ (
    .A1(\cpuregs[15] [5]),
    .A2(_12822_),
    .ZN(_13507_)
  );
  INV_X1 _48274_ (
    .A(_13507_),
    .ZN(_13508_)
  );
  AND2_X1 _48275_ (
    .A1(_13506_),
    .A2(_13508_),
    .ZN(_13509_)
  );
  INV_X1 _48276_ (
    .A(_13509_),
    .ZN(_00594_)
  );
  AND2_X1 _48277_ (
    .A1(_12821_),
    .A2(_12958_),
    .ZN(_13510_)
  );
  INV_X1 _48278_ (
    .A(_13510_),
    .ZN(_13511_)
  );
  AND2_X1 _48279_ (
    .A1(\cpuregs[15] [6]),
    .A2(_12822_),
    .ZN(_13512_)
  );
  INV_X1 _48280_ (
    .A(_13512_),
    .ZN(_13513_)
  );
  AND2_X1 _48281_ (
    .A1(_13511_),
    .A2(_13513_),
    .ZN(_13514_)
  );
  INV_X1 _48282_ (
    .A(_13514_),
    .ZN(_00595_)
  );
  AND2_X1 _48283_ (
    .A1(_12821_),
    .A2(_12973_),
    .ZN(_13515_)
  );
  INV_X1 _48284_ (
    .A(_13515_),
    .ZN(_13516_)
  );
  AND2_X1 _48285_ (
    .A1(\cpuregs[15] [7]),
    .A2(_12822_),
    .ZN(_13517_)
  );
  INV_X1 _48286_ (
    .A(_13517_),
    .ZN(_13518_)
  );
  AND2_X1 _48287_ (
    .A1(_13516_),
    .A2(_13518_),
    .ZN(_13519_)
  );
  INV_X1 _48288_ (
    .A(_13519_),
    .ZN(_00596_)
  );
  AND2_X1 _48289_ (
    .A1(_12821_),
    .A2(_12988_),
    .ZN(_13520_)
  );
  INV_X1 _48290_ (
    .A(_13520_),
    .ZN(_13521_)
  );
  AND2_X1 _48291_ (
    .A1(\cpuregs[15] [8]),
    .A2(_12822_),
    .ZN(_13522_)
  );
  INV_X1 _48292_ (
    .A(_13522_),
    .ZN(_13523_)
  );
  AND2_X1 _48293_ (
    .A1(_13521_),
    .A2(_13523_),
    .ZN(_13524_)
  );
  INV_X1 _48294_ (
    .A(_13524_),
    .ZN(_00597_)
  );
  AND2_X1 _48295_ (
    .A1(_12821_),
    .A2(_13003_),
    .ZN(_13525_)
  );
  INV_X1 _48296_ (
    .A(_13525_),
    .ZN(_13526_)
  );
  AND2_X1 _48297_ (
    .A1(\cpuregs[15] [9]),
    .A2(_12822_),
    .ZN(_13527_)
  );
  INV_X1 _48298_ (
    .A(_13527_),
    .ZN(_13528_)
  );
  AND2_X1 _48299_ (
    .A1(_13526_),
    .A2(_13528_),
    .ZN(_13529_)
  );
  INV_X1 _48300_ (
    .A(_13529_),
    .ZN(_00598_)
  );
  AND2_X1 _48301_ (
    .A1(_12821_),
    .A2(_13018_),
    .ZN(_13530_)
  );
  INV_X1 _48302_ (
    .A(_13530_),
    .ZN(_13531_)
  );
  AND2_X1 _48303_ (
    .A1(\cpuregs[15] [10]),
    .A2(_12822_),
    .ZN(_13532_)
  );
  INV_X1 _48304_ (
    .A(_13532_),
    .ZN(_13533_)
  );
  AND2_X1 _48305_ (
    .A1(_13531_),
    .A2(_13533_),
    .ZN(_13534_)
  );
  INV_X1 _48306_ (
    .A(_13534_),
    .ZN(_00599_)
  );
  AND2_X1 _48307_ (
    .A1(_12821_),
    .A2(_13033_),
    .ZN(_13535_)
  );
  INV_X1 _48308_ (
    .A(_13535_),
    .ZN(_13536_)
  );
  AND2_X1 _48309_ (
    .A1(\cpuregs[15] [11]),
    .A2(_12822_),
    .ZN(_13537_)
  );
  INV_X1 _48310_ (
    .A(_13537_),
    .ZN(_13538_)
  );
  AND2_X1 _48311_ (
    .A1(_13536_),
    .A2(_13538_),
    .ZN(_13539_)
  );
  INV_X1 _48312_ (
    .A(_13539_),
    .ZN(_00600_)
  );
  AND2_X1 _48313_ (
    .A1(_12821_),
    .A2(_13048_),
    .ZN(_13540_)
  );
  INV_X1 _48314_ (
    .A(_13540_),
    .ZN(_13541_)
  );
  AND2_X1 _48315_ (
    .A1(\cpuregs[15] [12]),
    .A2(_12822_),
    .ZN(_13542_)
  );
  INV_X1 _48316_ (
    .A(_13542_),
    .ZN(_13543_)
  );
  AND2_X1 _48317_ (
    .A1(_13541_),
    .A2(_13543_),
    .ZN(_13544_)
  );
  INV_X1 _48318_ (
    .A(_13544_),
    .ZN(_00601_)
  );
  AND2_X1 _48319_ (
    .A1(_12821_),
    .A2(_13063_),
    .ZN(_13545_)
  );
  INV_X1 _48320_ (
    .A(_13545_),
    .ZN(_13546_)
  );
  AND2_X1 _48321_ (
    .A1(\cpuregs[15] [13]),
    .A2(_12822_),
    .ZN(_13547_)
  );
  INV_X1 _48322_ (
    .A(_13547_),
    .ZN(_13548_)
  );
  AND2_X1 _48323_ (
    .A1(_13546_),
    .A2(_13548_),
    .ZN(_13549_)
  );
  INV_X1 _48324_ (
    .A(_13549_),
    .ZN(_00602_)
  );
  AND2_X1 _48325_ (
    .A1(_12821_),
    .A2(_13078_),
    .ZN(_13550_)
  );
  INV_X1 _48326_ (
    .A(_13550_),
    .ZN(_13551_)
  );
  AND2_X1 _48327_ (
    .A1(\cpuregs[15] [14]),
    .A2(_12822_),
    .ZN(_13552_)
  );
  INV_X1 _48328_ (
    .A(_13552_),
    .ZN(_13553_)
  );
  AND2_X1 _48329_ (
    .A1(_13551_),
    .A2(_13553_),
    .ZN(_13554_)
  );
  INV_X1 _48330_ (
    .A(_13554_),
    .ZN(_00603_)
  );
  AND2_X1 _48331_ (
    .A1(_12821_),
    .A2(_13093_),
    .ZN(_13555_)
  );
  INV_X1 _48332_ (
    .A(_13555_),
    .ZN(_13556_)
  );
  AND2_X1 _48333_ (
    .A1(\cpuregs[15] [15]),
    .A2(_12822_),
    .ZN(_13557_)
  );
  INV_X1 _48334_ (
    .A(_13557_),
    .ZN(_13558_)
  );
  AND2_X1 _48335_ (
    .A1(_13556_),
    .A2(_13558_),
    .ZN(_13559_)
  );
  INV_X1 _48336_ (
    .A(_13559_),
    .ZN(_00604_)
  );
  AND2_X1 _48337_ (
    .A1(_12821_),
    .A2(_13108_),
    .ZN(_13560_)
  );
  INV_X1 _48338_ (
    .A(_13560_),
    .ZN(_13561_)
  );
  AND2_X1 _48339_ (
    .A1(\cpuregs[15] [16]),
    .A2(_12822_),
    .ZN(_13562_)
  );
  INV_X1 _48340_ (
    .A(_13562_),
    .ZN(_13563_)
  );
  AND2_X1 _48341_ (
    .A1(_13561_),
    .A2(_13563_),
    .ZN(_13564_)
  );
  INV_X1 _48342_ (
    .A(_13564_),
    .ZN(_00605_)
  );
  AND2_X1 _48343_ (
    .A1(_21404_),
    .A2(_12822_),
    .ZN(_13565_)
  );
  INV_X1 _48344_ (
    .A(_13565_),
    .ZN(_13566_)
  );
  AND2_X1 _48345_ (
    .A1(_12821_),
    .A2(_13124_),
    .ZN(_13567_)
  );
  INV_X1 _48346_ (
    .A(_13567_),
    .ZN(_13568_)
  );
  AND2_X1 _48347_ (
    .A1(_13566_),
    .A2(_13568_),
    .ZN(_00606_)
  );
  AND2_X1 _48348_ (
    .A1(\cpuregs[15] [18]),
    .A2(_12822_),
    .ZN(_13569_)
  );
  INV_X1 _48349_ (
    .A(_13569_),
    .ZN(_13570_)
  );
  AND2_X1 _48350_ (
    .A1(_12821_),
    .A2(_13139_),
    .ZN(_13571_)
  );
  INV_X1 _48351_ (
    .A(_13571_),
    .ZN(_13572_)
  );
  AND2_X1 _48352_ (
    .A1(_13570_),
    .A2(_13572_),
    .ZN(_13573_)
  );
  INV_X1 _48353_ (
    .A(_13573_),
    .ZN(_00607_)
  );
  AND2_X1 _48354_ (
    .A1(\cpuregs[15] [19]),
    .A2(_12822_),
    .ZN(_13574_)
  );
  INV_X1 _48355_ (
    .A(_13574_),
    .ZN(_13575_)
  );
  AND2_X1 _48356_ (
    .A1(_12821_),
    .A2(_13154_),
    .ZN(_13576_)
  );
  INV_X1 _48357_ (
    .A(_13576_),
    .ZN(_13577_)
  );
  AND2_X1 _48358_ (
    .A1(_13575_),
    .A2(_13577_),
    .ZN(_13578_)
  );
  INV_X1 _48359_ (
    .A(_13578_),
    .ZN(_00608_)
  );
  AND2_X1 _48360_ (
    .A1(\cpuregs[15] [20]),
    .A2(_12822_),
    .ZN(_13579_)
  );
  INV_X1 _48361_ (
    .A(_13579_),
    .ZN(_13580_)
  );
  AND2_X1 _48362_ (
    .A1(_12821_),
    .A2(_13169_),
    .ZN(_13581_)
  );
  INV_X1 _48363_ (
    .A(_13581_),
    .ZN(_13582_)
  );
  AND2_X1 _48364_ (
    .A1(_13580_),
    .A2(_13582_),
    .ZN(_13583_)
  );
  INV_X1 _48365_ (
    .A(_13583_),
    .ZN(_00609_)
  );
  AND2_X1 _48366_ (
    .A1(\cpuregs[15] [21]),
    .A2(_12822_),
    .ZN(_13584_)
  );
  INV_X1 _48367_ (
    .A(_13584_),
    .ZN(_13585_)
  );
  AND2_X1 _48368_ (
    .A1(_12821_),
    .A2(_13184_),
    .ZN(_13586_)
  );
  INV_X1 _48369_ (
    .A(_13586_),
    .ZN(_13587_)
  );
  AND2_X1 _48370_ (
    .A1(_13585_),
    .A2(_13587_),
    .ZN(_13588_)
  );
  INV_X1 _48371_ (
    .A(_13588_),
    .ZN(_00610_)
  );
  AND2_X1 _48372_ (
    .A1(\cpuregs[15] [22]),
    .A2(_12822_),
    .ZN(_13589_)
  );
  INV_X1 _48373_ (
    .A(_13589_),
    .ZN(_13590_)
  );
  AND2_X1 _48374_ (
    .A1(_12821_),
    .A2(_13199_),
    .ZN(_13591_)
  );
  INV_X1 _48375_ (
    .A(_13591_),
    .ZN(_13592_)
  );
  AND2_X1 _48376_ (
    .A1(_13590_),
    .A2(_13592_),
    .ZN(_13593_)
  );
  INV_X1 _48377_ (
    .A(_13593_),
    .ZN(_00611_)
  );
  AND2_X1 _48378_ (
    .A1(\cpuregs[15] [23]),
    .A2(_12822_),
    .ZN(_13594_)
  );
  INV_X1 _48379_ (
    .A(_13594_),
    .ZN(_13595_)
  );
  AND2_X1 _48380_ (
    .A1(_12821_),
    .A2(_13214_),
    .ZN(_13596_)
  );
  INV_X1 _48381_ (
    .A(_13596_),
    .ZN(_13597_)
  );
  AND2_X1 _48382_ (
    .A1(_13595_),
    .A2(_13597_),
    .ZN(_13598_)
  );
  INV_X1 _48383_ (
    .A(_13598_),
    .ZN(_00612_)
  );
  AND2_X1 _48384_ (
    .A1(\cpuregs[15] [24]),
    .A2(_12822_),
    .ZN(_13599_)
  );
  INV_X1 _48385_ (
    .A(_13599_),
    .ZN(_13600_)
  );
  AND2_X1 _48386_ (
    .A1(_12821_),
    .A2(_13229_),
    .ZN(_13601_)
  );
  INV_X1 _48387_ (
    .A(_13601_),
    .ZN(_13602_)
  );
  AND2_X1 _48388_ (
    .A1(_13600_),
    .A2(_13602_),
    .ZN(_13603_)
  );
  INV_X1 _48389_ (
    .A(_13603_),
    .ZN(_00613_)
  );
  AND2_X1 _48390_ (
    .A1(\cpuregs[15] [25]),
    .A2(_12822_),
    .ZN(_13604_)
  );
  INV_X1 _48391_ (
    .A(_13604_),
    .ZN(_13605_)
  );
  AND2_X1 _48392_ (
    .A1(_12821_),
    .A2(_13244_),
    .ZN(_13606_)
  );
  INV_X1 _48393_ (
    .A(_13606_),
    .ZN(_13607_)
  );
  AND2_X1 _48394_ (
    .A1(_13605_),
    .A2(_13607_),
    .ZN(_13608_)
  );
  INV_X1 _48395_ (
    .A(_13608_),
    .ZN(_00614_)
  );
  AND2_X1 _48396_ (
    .A1(\cpuregs[15] [26]),
    .A2(_12822_),
    .ZN(_13609_)
  );
  INV_X1 _48397_ (
    .A(_13609_),
    .ZN(_13610_)
  );
  AND2_X1 _48398_ (
    .A1(_12821_),
    .A2(_13259_),
    .ZN(_13611_)
  );
  INV_X1 _48399_ (
    .A(_13611_),
    .ZN(_13612_)
  );
  AND2_X1 _48400_ (
    .A1(_13610_),
    .A2(_13612_),
    .ZN(_13613_)
  );
  INV_X1 _48401_ (
    .A(_13613_),
    .ZN(_00615_)
  );
  AND2_X1 _48402_ (
    .A1(\cpuregs[15] [27]),
    .A2(_12822_),
    .ZN(_13614_)
  );
  INV_X1 _48403_ (
    .A(_13614_),
    .ZN(_13615_)
  );
  AND2_X1 _48404_ (
    .A1(_12821_),
    .A2(_13274_),
    .ZN(_13616_)
  );
  INV_X1 _48405_ (
    .A(_13616_),
    .ZN(_13617_)
  );
  AND2_X1 _48406_ (
    .A1(_13615_),
    .A2(_13617_),
    .ZN(_13618_)
  );
  INV_X1 _48407_ (
    .A(_13618_),
    .ZN(_00616_)
  );
  AND2_X1 _48408_ (
    .A1(\cpuregs[15] [28]),
    .A2(_12822_),
    .ZN(_13619_)
  );
  INV_X1 _48409_ (
    .A(_13619_),
    .ZN(_13620_)
  );
  AND2_X1 _48410_ (
    .A1(_12821_),
    .A2(_13289_),
    .ZN(_13621_)
  );
  INV_X1 _48411_ (
    .A(_13621_),
    .ZN(_13622_)
  );
  AND2_X1 _48412_ (
    .A1(_13620_),
    .A2(_13622_),
    .ZN(_13623_)
  );
  INV_X1 _48413_ (
    .A(_13623_),
    .ZN(_00617_)
  );
  AND2_X1 _48414_ (
    .A1(\cpuregs[15] [29]),
    .A2(_12822_),
    .ZN(_13624_)
  );
  INV_X1 _48415_ (
    .A(_13624_),
    .ZN(_13625_)
  );
  AND2_X1 _48416_ (
    .A1(_12821_),
    .A2(_13304_),
    .ZN(_13626_)
  );
  INV_X1 _48417_ (
    .A(_13626_),
    .ZN(_13627_)
  );
  AND2_X1 _48418_ (
    .A1(_13625_),
    .A2(_13627_),
    .ZN(_13628_)
  );
  INV_X1 _48419_ (
    .A(_13628_),
    .ZN(_00618_)
  );
  AND2_X1 _48420_ (
    .A1(\cpuregs[15] [30]),
    .A2(_12822_),
    .ZN(_13629_)
  );
  INV_X1 _48421_ (
    .A(_13629_),
    .ZN(_13630_)
  );
  AND2_X1 _48422_ (
    .A1(_12821_),
    .A2(_13319_),
    .ZN(_13631_)
  );
  INV_X1 _48423_ (
    .A(_13631_),
    .ZN(_13632_)
  );
  AND2_X1 _48424_ (
    .A1(_13630_),
    .A2(_13632_),
    .ZN(_13633_)
  );
  INV_X1 _48425_ (
    .A(_13633_),
    .ZN(_00619_)
  );
  AND2_X1 _48426_ (
    .A1(_12762_),
    .A2(_12872_),
    .ZN(_13634_)
  );
  INV_X1 _48427_ (
    .A(_13634_),
    .ZN(_13635_)
  );
  AND2_X1 _48428_ (
    .A1(_21408_),
    .A2(_12763_),
    .ZN(_13636_)
  );
  INV_X1 _48429_ (
    .A(_13636_),
    .ZN(_13637_)
  );
  AND2_X1 _48430_ (
    .A1(_13635_),
    .A2(_13637_),
    .ZN(_00620_)
  );
  AND2_X1 _48431_ (
    .A1(_12762_),
    .A2(_12884_),
    .ZN(_13638_)
  );
  INV_X1 _48432_ (
    .A(_13638_),
    .ZN(_13639_)
  );
  AND2_X1 _48433_ (
    .A1(_21409_),
    .A2(_12763_),
    .ZN(_13640_)
  );
  INV_X1 _48434_ (
    .A(_13640_),
    .ZN(_13641_)
  );
  AND2_X1 _48435_ (
    .A1(_13639_),
    .A2(_13641_),
    .ZN(_00621_)
  );
  AND2_X1 _48436_ (
    .A1(_12762_),
    .A2(_12898_),
    .ZN(_13642_)
  );
  INV_X1 _48437_ (
    .A(_13642_),
    .ZN(_13643_)
  );
  AND2_X1 _48438_ (
    .A1(_21410_),
    .A2(_12763_),
    .ZN(_13644_)
  );
  INV_X1 _48439_ (
    .A(_13644_),
    .ZN(_13645_)
  );
  AND2_X1 _48440_ (
    .A1(_13643_),
    .A2(_13645_),
    .ZN(_00622_)
  );
  AND2_X1 _48441_ (
    .A1(_12762_),
    .A2(_12911_),
    .ZN(_13646_)
  );
  INV_X1 _48442_ (
    .A(_13646_),
    .ZN(_13647_)
  );
  AND2_X1 _48443_ (
    .A1(_21411_),
    .A2(_12763_),
    .ZN(_13648_)
  );
  INV_X1 _48444_ (
    .A(_13648_),
    .ZN(_13649_)
  );
  AND2_X1 _48445_ (
    .A1(_13647_),
    .A2(_13649_),
    .ZN(_00623_)
  );
  AND2_X1 _48446_ (
    .A1(_12762_),
    .A2(_12928_),
    .ZN(_13650_)
  );
  INV_X1 _48447_ (
    .A(_13650_),
    .ZN(_13651_)
  );
  AND2_X1 _48448_ (
    .A1(\cpuregs[22] [4]),
    .A2(_12763_),
    .ZN(_13652_)
  );
  INV_X1 _48449_ (
    .A(_13652_),
    .ZN(_13653_)
  );
  AND2_X1 _48450_ (
    .A1(_13651_),
    .A2(_13653_),
    .ZN(_13654_)
  );
  INV_X1 _48451_ (
    .A(_13654_),
    .ZN(_00624_)
  );
  AND2_X1 _48452_ (
    .A1(_12762_),
    .A2(_12941_),
    .ZN(_13655_)
  );
  INV_X1 _48453_ (
    .A(_13655_),
    .ZN(_13656_)
  );
  AND2_X1 _48454_ (
    .A1(_21413_),
    .A2(_12763_),
    .ZN(_13657_)
  );
  INV_X1 _48455_ (
    .A(_13657_),
    .ZN(_13658_)
  );
  AND2_X1 _48456_ (
    .A1(_13656_),
    .A2(_13658_),
    .ZN(_00625_)
  );
  AND2_X1 _48457_ (
    .A1(_12762_),
    .A2(_12956_),
    .ZN(_13659_)
  );
  INV_X1 _48458_ (
    .A(_13659_),
    .ZN(_13660_)
  );
  AND2_X1 _48459_ (
    .A1(_21414_),
    .A2(_12763_),
    .ZN(_13661_)
  );
  INV_X1 _48460_ (
    .A(_13661_),
    .ZN(_13662_)
  );
  AND2_X1 _48461_ (
    .A1(_13660_),
    .A2(_13662_),
    .ZN(_00626_)
  );
  AND2_X1 _48462_ (
    .A1(_12762_),
    .A2(_12971_),
    .ZN(_13663_)
  );
  INV_X1 _48463_ (
    .A(_13663_),
    .ZN(_13664_)
  );
  AND2_X1 _48464_ (
    .A1(_21415_),
    .A2(_12763_),
    .ZN(_13665_)
  );
  INV_X1 _48465_ (
    .A(_13665_),
    .ZN(_13666_)
  );
  AND2_X1 _48466_ (
    .A1(_13664_),
    .A2(_13666_),
    .ZN(_00627_)
  );
  AND2_X1 _48467_ (
    .A1(_12762_),
    .A2(_12986_),
    .ZN(_13667_)
  );
  INV_X1 _48468_ (
    .A(_13667_),
    .ZN(_13668_)
  );
  AND2_X1 _48469_ (
    .A1(_21416_),
    .A2(_12763_),
    .ZN(_13669_)
  );
  INV_X1 _48470_ (
    .A(_13669_),
    .ZN(_13670_)
  );
  AND2_X1 _48471_ (
    .A1(_13668_),
    .A2(_13670_),
    .ZN(_00628_)
  );
  AND2_X1 _48472_ (
    .A1(_12762_),
    .A2(_13001_),
    .ZN(_13671_)
  );
  INV_X1 _48473_ (
    .A(_13671_),
    .ZN(_13672_)
  );
  AND2_X1 _48474_ (
    .A1(_21417_),
    .A2(_12763_),
    .ZN(_13673_)
  );
  INV_X1 _48475_ (
    .A(_13673_),
    .ZN(_13674_)
  );
  AND2_X1 _48476_ (
    .A1(_13672_),
    .A2(_13674_),
    .ZN(_00629_)
  );
  AND2_X1 _48477_ (
    .A1(_12762_),
    .A2(_13016_),
    .ZN(_13675_)
  );
  INV_X1 _48478_ (
    .A(_13675_),
    .ZN(_13676_)
  );
  AND2_X1 _48479_ (
    .A1(_21418_),
    .A2(_12763_),
    .ZN(_13677_)
  );
  INV_X1 _48480_ (
    .A(_13677_),
    .ZN(_13678_)
  );
  AND2_X1 _48481_ (
    .A1(_13676_),
    .A2(_13678_),
    .ZN(_00630_)
  );
  AND2_X1 _48482_ (
    .A1(_12762_),
    .A2(_13033_),
    .ZN(_13679_)
  );
  INV_X1 _48483_ (
    .A(_13679_),
    .ZN(_13680_)
  );
  AND2_X1 _48484_ (
    .A1(\cpuregs[22] [11]),
    .A2(_12763_),
    .ZN(_13681_)
  );
  INV_X1 _48485_ (
    .A(_13681_),
    .ZN(_13682_)
  );
  AND2_X1 _48486_ (
    .A1(_13680_),
    .A2(_13682_),
    .ZN(_13683_)
  );
  INV_X1 _48487_ (
    .A(_13683_),
    .ZN(_00631_)
  );
  AND2_X1 _48488_ (
    .A1(_12762_),
    .A2(_13046_),
    .ZN(_13684_)
  );
  INV_X1 _48489_ (
    .A(_13684_),
    .ZN(_13685_)
  );
  AND2_X1 _48490_ (
    .A1(_21419_),
    .A2(_12763_),
    .ZN(_13686_)
  );
  INV_X1 _48491_ (
    .A(_13686_),
    .ZN(_13687_)
  );
  AND2_X1 _48492_ (
    .A1(_13685_),
    .A2(_13687_),
    .ZN(_00632_)
  );
  AND2_X1 _48493_ (
    .A1(_12762_),
    .A2(_13061_),
    .ZN(_13688_)
  );
  INV_X1 _48494_ (
    .A(_13688_),
    .ZN(_13689_)
  );
  AND2_X1 _48495_ (
    .A1(_21420_),
    .A2(_12763_),
    .ZN(_13690_)
  );
  INV_X1 _48496_ (
    .A(_13690_),
    .ZN(_13691_)
  );
  AND2_X1 _48497_ (
    .A1(_13689_),
    .A2(_13691_),
    .ZN(_00633_)
  );
  AND2_X1 _48498_ (
    .A1(_12762_),
    .A2(_13076_),
    .ZN(_13692_)
  );
  INV_X1 _48499_ (
    .A(_13692_),
    .ZN(_13693_)
  );
  AND2_X1 _48500_ (
    .A1(_21421_),
    .A2(_12763_),
    .ZN(_13694_)
  );
  INV_X1 _48501_ (
    .A(_13694_),
    .ZN(_13695_)
  );
  AND2_X1 _48502_ (
    .A1(_13693_),
    .A2(_13695_),
    .ZN(_00634_)
  );
  AND2_X1 _48503_ (
    .A1(_12762_),
    .A2(_13091_),
    .ZN(_13696_)
  );
  INV_X1 _48504_ (
    .A(_13696_),
    .ZN(_13697_)
  );
  AND2_X1 _48505_ (
    .A1(_21422_),
    .A2(_12763_),
    .ZN(_13698_)
  );
  INV_X1 _48506_ (
    .A(_13698_),
    .ZN(_13699_)
  );
  AND2_X1 _48507_ (
    .A1(_13697_),
    .A2(_13699_),
    .ZN(_00635_)
  );
  AND2_X1 _48508_ (
    .A1(_12762_),
    .A2(_13108_),
    .ZN(_13700_)
  );
  INV_X1 _48509_ (
    .A(_13700_),
    .ZN(_13701_)
  );
  AND2_X1 _48510_ (
    .A1(\cpuregs[22] [16]),
    .A2(_12763_),
    .ZN(_13702_)
  );
  INV_X1 _48511_ (
    .A(_13702_),
    .ZN(_13703_)
  );
  AND2_X1 _48512_ (
    .A1(_13701_),
    .A2(_13703_),
    .ZN(_13704_)
  );
  INV_X1 _48513_ (
    .A(_13704_),
    .ZN(_00636_)
  );
  AND2_X1 _48514_ (
    .A1(_12762_),
    .A2(_13121_),
    .ZN(_13705_)
  );
  INV_X1 _48515_ (
    .A(_13705_),
    .ZN(_13706_)
  );
  AND2_X1 _48516_ (
    .A1(_21424_),
    .A2(_12763_),
    .ZN(_13707_)
  );
  INV_X1 _48517_ (
    .A(_13707_),
    .ZN(_13708_)
  );
  AND2_X1 _48518_ (
    .A1(_13706_),
    .A2(_13708_),
    .ZN(_00637_)
  );
  AND2_X1 _48519_ (
    .A1(_12762_),
    .A2(_13139_),
    .ZN(_13709_)
  );
  INV_X1 _48520_ (
    .A(_13709_),
    .ZN(_13710_)
  );
  AND2_X1 _48521_ (
    .A1(\cpuregs[22] [18]),
    .A2(_12763_),
    .ZN(_13711_)
  );
  INV_X1 _48522_ (
    .A(_13711_),
    .ZN(_13712_)
  );
  AND2_X1 _48523_ (
    .A1(_13710_),
    .A2(_13712_),
    .ZN(_13713_)
  );
  INV_X1 _48524_ (
    .A(_13713_),
    .ZN(_00638_)
  );
  AND2_X1 _48525_ (
    .A1(_21425_),
    .A2(_12763_),
    .ZN(_13714_)
  );
  INV_X1 _48526_ (
    .A(_13714_),
    .ZN(_13715_)
  );
  AND2_X1 _48527_ (
    .A1(_12762_),
    .A2(_13152_),
    .ZN(_13716_)
  );
  INV_X1 _48528_ (
    .A(_13716_),
    .ZN(_13717_)
  );
  AND2_X1 _48529_ (
    .A1(_13715_),
    .A2(_13717_),
    .ZN(_00639_)
  );
  AND2_X1 _48530_ (
    .A1(_12762_),
    .A2(_13169_),
    .ZN(_13718_)
  );
  INV_X1 _48531_ (
    .A(_13718_),
    .ZN(_13719_)
  );
  AND2_X1 _48532_ (
    .A1(\cpuregs[22] [20]),
    .A2(_12763_),
    .ZN(_13720_)
  );
  INV_X1 _48533_ (
    .A(_13720_),
    .ZN(_13721_)
  );
  AND2_X1 _48534_ (
    .A1(_13719_),
    .A2(_13721_),
    .ZN(_13722_)
  );
  INV_X1 _48535_ (
    .A(_13722_),
    .ZN(_00640_)
  );
  AND2_X1 _48536_ (
    .A1(_12762_),
    .A2(_13184_),
    .ZN(_13723_)
  );
  INV_X1 _48537_ (
    .A(_13723_),
    .ZN(_13724_)
  );
  AND2_X1 _48538_ (
    .A1(\cpuregs[22] [21]),
    .A2(_12763_),
    .ZN(_13725_)
  );
  INV_X1 _48539_ (
    .A(_13725_),
    .ZN(_13726_)
  );
  AND2_X1 _48540_ (
    .A1(_13724_),
    .A2(_13726_),
    .ZN(_13727_)
  );
  INV_X1 _48541_ (
    .A(_13727_),
    .ZN(_00641_)
  );
  AND2_X1 _48542_ (
    .A1(_12762_),
    .A2(_13197_),
    .ZN(_13728_)
  );
  INV_X1 _48543_ (
    .A(_13728_),
    .ZN(_13729_)
  );
  AND2_X1 _48544_ (
    .A1(_21427_),
    .A2(_12763_),
    .ZN(_13730_)
  );
  INV_X1 _48545_ (
    .A(_13730_),
    .ZN(_13731_)
  );
  AND2_X1 _48546_ (
    .A1(_13729_),
    .A2(_13731_),
    .ZN(_00642_)
  );
  AND2_X1 _48547_ (
    .A1(_12762_),
    .A2(_13212_),
    .ZN(_13732_)
  );
  INV_X1 _48548_ (
    .A(_13732_),
    .ZN(_13733_)
  );
  AND2_X1 _48549_ (
    .A1(_21428_),
    .A2(_12763_),
    .ZN(_13734_)
  );
  INV_X1 _48550_ (
    .A(_13734_),
    .ZN(_13735_)
  );
  AND2_X1 _48551_ (
    .A1(_13733_),
    .A2(_13735_),
    .ZN(_00643_)
  );
  AND2_X1 _48552_ (
    .A1(_12762_),
    .A2(_13227_),
    .ZN(_13736_)
  );
  INV_X1 _48553_ (
    .A(_13736_),
    .ZN(_13737_)
  );
  AND2_X1 _48554_ (
    .A1(_21429_),
    .A2(_12763_),
    .ZN(_13738_)
  );
  INV_X1 _48555_ (
    .A(_13738_),
    .ZN(_13739_)
  );
  AND2_X1 _48556_ (
    .A1(_13737_),
    .A2(_13739_),
    .ZN(_00644_)
  );
  AND2_X1 _48557_ (
    .A1(_12762_),
    .A2(_13242_),
    .ZN(_13740_)
  );
  INV_X1 _48558_ (
    .A(_13740_),
    .ZN(_13741_)
  );
  AND2_X1 _48559_ (
    .A1(_21430_),
    .A2(_12763_),
    .ZN(_13742_)
  );
  INV_X1 _48560_ (
    .A(_13742_),
    .ZN(_13743_)
  );
  AND2_X1 _48561_ (
    .A1(_13741_),
    .A2(_13743_),
    .ZN(_00645_)
  );
  AND2_X1 _48562_ (
    .A1(_12762_),
    .A2(_13257_),
    .ZN(_13744_)
  );
  INV_X1 _48563_ (
    .A(_13744_),
    .ZN(_13745_)
  );
  AND2_X1 _48564_ (
    .A1(_21431_),
    .A2(_12763_),
    .ZN(_13746_)
  );
  INV_X1 _48565_ (
    .A(_13746_),
    .ZN(_13747_)
  );
  AND2_X1 _48566_ (
    .A1(_13745_),
    .A2(_13747_),
    .ZN(_00646_)
  );
  AND2_X1 _48567_ (
    .A1(_12762_),
    .A2(_13272_),
    .ZN(_13748_)
  );
  INV_X1 _48568_ (
    .A(_13748_),
    .ZN(_13749_)
  );
  AND2_X1 _48569_ (
    .A1(_21432_),
    .A2(_12763_),
    .ZN(_13750_)
  );
  INV_X1 _48570_ (
    .A(_13750_),
    .ZN(_13751_)
  );
  AND2_X1 _48571_ (
    .A1(_13749_),
    .A2(_13751_),
    .ZN(_00647_)
  );
  AND2_X1 _48572_ (
    .A1(_12762_),
    .A2(_13287_),
    .ZN(_13752_)
  );
  INV_X1 _48573_ (
    .A(_13752_),
    .ZN(_13753_)
  );
  AND2_X1 _48574_ (
    .A1(_21433_),
    .A2(_12763_),
    .ZN(_13754_)
  );
  INV_X1 _48575_ (
    .A(_13754_),
    .ZN(_13755_)
  );
  AND2_X1 _48576_ (
    .A1(_13753_),
    .A2(_13755_),
    .ZN(_00648_)
  );
  AND2_X1 _48577_ (
    .A1(_12762_),
    .A2(_13302_),
    .ZN(_13756_)
  );
  INV_X1 _48578_ (
    .A(_13756_),
    .ZN(_13757_)
  );
  AND2_X1 _48579_ (
    .A1(_21434_),
    .A2(_12763_),
    .ZN(_13758_)
  );
  INV_X1 _48580_ (
    .A(_13758_),
    .ZN(_13759_)
  );
  AND2_X1 _48581_ (
    .A1(_13757_),
    .A2(_13759_),
    .ZN(_00649_)
  );
  AND2_X1 _48582_ (
    .A1(_12762_),
    .A2(_13317_),
    .ZN(_13760_)
  );
  INV_X1 _48583_ (
    .A(_13760_),
    .ZN(_13761_)
  );
  AND2_X1 _48584_ (
    .A1(_21435_),
    .A2(_12763_),
    .ZN(_13762_)
  );
  INV_X1 _48585_ (
    .A(_13762_),
    .ZN(_13763_)
  );
  AND2_X1 _48586_ (
    .A1(_13761_),
    .A2(_13763_),
    .ZN(_00650_)
  );
  AND2_X1 _48587_ (
    .A1(_12812_),
    .A2(_12874_),
    .ZN(_13764_)
  );
  INV_X1 _48588_ (
    .A(_13764_),
    .ZN(_13765_)
  );
  AND2_X1 _48589_ (
    .A1(\cpuregs[16] [0]),
    .A2(_12813_),
    .ZN(_13766_)
  );
  INV_X1 _48590_ (
    .A(_13766_),
    .ZN(_13767_)
  );
  AND2_X1 _48591_ (
    .A1(_13765_),
    .A2(_13767_),
    .ZN(_13768_)
  );
  INV_X1 _48592_ (
    .A(_13768_),
    .ZN(_00651_)
  );
  AND2_X1 _48593_ (
    .A1(\cpuregs[16] [1]),
    .A2(_12813_),
    .ZN(_13769_)
  );
  INV_X1 _48594_ (
    .A(_13769_),
    .ZN(_13770_)
  );
  AND2_X1 _48595_ (
    .A1(_12812_),
    .A2(_12886_),
    .ZN(_13771_)
  );
  INV_X1 _48596_ (
    .A(_13771_),
    .ZN(_13772_)
  );
  AND2_X1 _48597_ (
    .A1(_13770_),
    .A2(_13772_),
    .ZN(_13773_)
  );
  INV_X1 _48598_ (
    .A(_13773_),
    .ZN(_00652_)
  );
  AND2_X1 _48599_ (
    .A1(\cpuregs[16] [2]),
    .A2(_12813_),
    .ZN(_13774_)
  );
  INV_X1 _48600_ (
    .A(_13774_),
    .ZN(_13775_)
  );
  AND2_X1 _48601_ (
    .A1(_12812_),
    .A2(_12900_),
    .ZN(_13776_)
  );
  INV_X1 _48602_ (
    .A(_13776_),
    .ZN(_13777_)
  );
  AND2_X1 _48603_ (
    .A1(_13775_),
    .A2(_13777_),
    .ZN(_13778_)
  );
  INV_X1 _48604_ (
    .A(_13778_),
    .ZN(_00653_)
  );
  AND2_X1 _48605_ (
    .A1(\cpuregs[16] [3]),
    .A2(_12813_),
    .ZN(_13779_)
  );
  INV_X1 _48606_ (
    .A(_13779_),
    .ZN(_13780_)
  );
  AND2_X1 _48607_ (
    .A1(_12812_),
    .A2(_12913_),
    .ZN(_13781_)
  );
  INV_X1 _48608_ (
    .A(_13781_),
    .ZN(_13782_)
  );
  AND2_X1 _48609_ (
    .A1(_13780_),
    .A2(_13782_),
    .ZN(_13783_)
  );
  INV_X1 _48610_ (
    .A(_13783_),
    .ZN(_00654_)
  );
  AND2_X1 _48611_ (
    .A1(_12812_),
    .A2(_12928_),
    .ZN(_13784_)
  );
  INV_X1 _48612_ (
    .A(_13784_),
    .ZN(_13785_)
  );
  AND2_X1 _48613_ (
    .A1(\cpuregs[16] [4]),
    .A2(_12813_),
    .ZN(_13786_)
  );
  INV_X1 _48614_ (
    .A(_13786_),
    .ZN(_13787_)
  );
  AND2_X1 _48615_ (
    .A1(_13785_),
    .A2(_13787_),
    .ZN(_13788_)
  );
  INV_X1 _48616_ (
    .A(_13788_),
    .ZN(_00655_)
  );
  AND2_X1 _48617_ (
    .A1(\cpuregs[16] [5]),
    .A2(_12813_),
    .ZN(_13789_)
  );
  INV_X1 _48618_ (
    .A(_13789_),
    .ZN(_13790_)
  );
  AND2_X1 _48619_ (
    .A1(_12812_),
    .A2(_12943_),
    .ZN(_13791_)
  );
  INV_X1 _48620_ (
    .A(_13791_),
    .ZN(_13792_)
  );
  AND2_X1 _48621_ (
    .A1(_13790_),
    .A2(_13792_),
    .ZN(_13793_)
  );
  INV_X1 _48622_ (
    .A(_13793_),
    .ZN(_00656_)
  );
  AND2_X1 _48623_ (
    .A1(\cpuregs[16] [6]),
    .A2(_12813_),
    .ZN(_13794_)
  );
  INV_X1 _48624_ (
    .A(_13794_),
    .ZN(_13795_)
  );
  AND2_X1 _48625_ (
    .A1(_12812_),
    .A2(_12958_),
    .ZN(_13796_)
  );
  INV_X1 _48626_ (
    .A(_13796_),
    .ZN(_13797_)
  );
  AND2_X1 _48627_ (
    .A1(_13795_),
    .A2(_13797_),
    .ZN(_13798_)
  );
  INV_X1 _48628_ (
    .A(_13798_),
    .ZN(_00657_)
  );
  AND2_X1 _48629_ (
    .A1(_12812_),
    .A2(_12973_),
    .ZN(_13799_)
  );
  INV_X1 _48630_ (
    .A(_13799_),
    .ZN(_13800_)
  );
  AND2_X1 _48631_ (
    .A1(\cpuregs[16] [7]),
    .A2(_12813_),
    .ZN(_13801_)
  );
  INV_X1 _48632_ (
    .A(_13801_),
    .ZN(_13802_)
  );
  AND2_X1 _48633_ (
    .A1(_13800_),
    .A2(_13802_),
    .ZN(_13803_)
  );
  INV_X1 _48634_ (
    .A(_13803_),
    .ZN(_00658_)
  );
  AND2_X1 _48635_ (
    .A1(\cpuregs[16] [8]),
    .A2(_12813_),
    .ZN(_13804_)
  );
  INV_X1 _48636_ (
    .A(_13804_),
    .ZN(_13805_)
  );
  AND2_X1 _48637_ (
    .A1(_12812_),
    .A2(_12988_),
    .ZN(_13806_)
  );
  INV_X1 _48638_ (
    .A(_13806_),
    .ZN(_13807_)
  );
  AND2_X1 _48639_ (
    .A1(_13805_),
    .A2(_13807_),
    .ZN(_13808_)
  );
  INV_X1 _48640_ (
    .A(_13808_),
    .ZN(_00659_)
  );
  AND2_X1 _48641_ (
    .A1(\cpuregs[16] [9]),
    .A2(_12813_),
    .ZN(_13809_)
  );
  INV_X1 _48642_ (
    .A(_13809_),
    .ZN(_13810_)
  );
  AND2_X1 _48643_ (
    .A1(_12812_),
    .A2(_13003_),
    .ZN(_13811_)
  );
  INV_X1 _48644_ (
    .A(_13811_),
    .ZN(_13812_)
  );
  AND2_X1 _48645_ (
    .A1(_13810_),
    .A2(_13812_),
    .ZN(_13813_)
  );
  INV_X1 _48646_ (
    .A(_13813_),
    .ZN(_00660_)
  );
  AND2_X1 _48647_ (
    .A1(_12812_),
    .A2(_13018_),
    .ZN(_13814_)
  );
  INV_X1 _48648_ (
    .A(_13814_),
    .ZN(_13815_)
  );
  AND2_X1 _48649_ (
    .A1(\cpuregs[16] [10]),
    .A2(_12813_),
    .ZN(_13816_)
  );
  INV_X1 _48650_ (
    .A(_13816_),
    .ZN(_13817_)
  );
  AND2_X1 _48651_ (
    .A1(_13815_),
    .A2(_13817_),
    .ZN(_13818_)
  );
  INV_X1 _48652_ (
    .A(_13818_),
    .ZN(_00661_)
  );
  AND2_X1 _48653_ (
    .A1(\cpuregs[16] [11]),
    .A2(_12813_),
    .ZN(_13819_)
  );
  INV_X1 _48654_ (
    .A(_13819_),
    .ZN(_13820_)
  );
  AND2_X1 _48655_ (
    .A1(_12812_),
    .A2(_13033_),
    .ZN(_13821_)
  );
  INV_X1 _48656_ (
    .A(_13821_),
    .ZN(_13822_)
  );
  AND2_X1 _48657_ (
    .A1(_13820_),
    .A2(_13822_),
    .ZN(_13823_)
  );
  INV_X1 _48658_ (
    .A(_13823_),
    .ZN(_00662_)
  );
  AND2_X1 _48659_ (
    .A1(_12812_),
    .A2(_13048_),
    .ZN(_13824_)
  );
  INV_X1 _48660_ (
    .A(_13824_),
    .ZN(_13825_)
  );
  AND2_X1 _48661_ (
    .A1(\cpuregs[16] [12]),
    .A2(_12813_),
    .ZN(_13826_)
  );
  INV_X1 _48662_ (
    .A(_13826_),
    .ZN(_13827_)
  );
  AND2_X1 _48663_ (
    .A1(_13825_),
    .A2(_13827_),
    .ZN(_13828_)
  );
  INV_X1 _48664_ (
    .A(_13828_),
    .ZN(_00663_)
  );
  AND2_X1 _48665_ (
    .A1(\cpuregs[16] [13]),
    .A2(_12813_),
    .ZN(_13829_)
  );
  INV_X1 _48666_ (
    .A(_13829_),
    .ZN(_13830_)
  );
  AND2_X1 _48667_ (
    .A1(_12812_),
    .A2(_13063_),
    .ZN(_13831_)
  );
  INV_X1 _48668_ (
    .A(_13831_),
    .ZN(_13832_)
  );
  AND2_X1 _48669_ (
    .A1(_13830_),
    .A2(_13832_),
    .ZN(_13833_)
  );
  INV_X1 _48670_ (
    .A(_13833_),
    .ZN(_00664_)
  );
  AND2_X1 _48671_ (
    .A1(\cpuregs[16] [14]),
    .A2(_12813_),
    .ZN(_13834_)
  );
  INV_X1 _48672_ (
    .A(_13834_),
    .ZN(_13835_)
  );
  AND2_X1 _48673_ (
    .A1(_12812_),
    .A2(_13078_),
    .ZN(_13836_)
  );
  INV_X1 _48674_ (
    .A(_13836_),
    .ZN(_13837_)
  );
  AND2_X1 _48675_ (
    .A1(_13835_),
    .A2(_13837_),
    .ZN(_13838_)
  );
  INV_X1 _48676_ (
    .A(_13838_),
    .ZN(_00665_)
  );
  AND2_X1 _48677_ (
    .A1(_12812_),
    .A2(_13093_),
    .ZN(_13839_)
  );
  INV_X1 _48678_ (
    .A(_13839_),
    .ZN(_13840_)
  );
  AND2_X1 _48679_ (
    .A1(\cpuregs[16] [15]),
    .A2(_12813_),
    .ZN(_13841_)
  );
  INV_X1 _48680_ (
    .A(_13841_),
    .ZN(_13842_)
  );
  AND2_X1 _48681_ (
    .A1(_13840_),
    .A2(_13842_),
    .ZN(_13843_)
  );
  INV_X1 _48682_ (
    .A(_13843_),
    .ZN(_00666_)
  );
  AND2_X1 _48683_ (
    .A1(_12812_),
    .A2(_13108_),
    .ZN(_13844_)
  );
  INV_X1 _48684_ (
    .A(_13844_),
    .ZN(_13845_)
  );
  AND2_X1 _48685_ (
    .A1(\cpuregs[16] [16]),
    .A2(_12813_),
    .ZN(_13846_)
  );
  INV_X1 _48686_ (
    .A(_13846_),
    .ZN(_13847_)
  );
  AND2_X1 _48687_ (
    .A1(_13845_),
    .A2(_13847_),
    .ZN(_13848_)
  );
  INV_X1 _48688_ (
    .A(_13848_),
    .ZN(_00667_)
  );
  AND2_X1 _48689_ (
    .A1(_12812_),
    .A2(_13123_),
    .ZN(_13849_)
  );
  INV_X1 _48690_ (
    .A(_13849_),
    .ZN(_13850_)
  );
  AND2_X1 _48691_ (
    .A1(\cpuregs[16] [17]),
    .A2(_12813_),
    .ZN(_13851_)
  );
  INV_X1 _48692_ (
    .A(_13851_),
    .ZN(_13852_)
  );
  AND2_X1 _48693_ (
    .A1(_13850_),
    .A2(_13852_),
    .ZN(_13853_)
  );
  INV_X1 _48694_ (
    .A(_13853_),
    .ZN(_00668_)
  );
  AND2_X1 _48695_ (
    .A1(_12812_),
    .A2(_13139_),
    .ZN(_13854_)
  );
  INV_X1 _48696_ (
    .A(_13854_),
    .ZN(_13855_)
  );
  AND2_X1 _48697_ (
    .A1(\cpuregs[16] [18]),
    .A2(_12813_),
    .ZN(_13856_)
  );
  INV_X1 _48698_ (
    .A(_13856_),
    .ZN(_13857_)
  );
  AND2_X1 _48699_ (
    .A1(_13855_),
    .A2(_13857_),
    .ZN(_13858_)
  );
  INV_X1 _48700_ (
    .A(_13858_),
    .ZN(_00669_)
  );
  AND2_X1 _48701_ (
    .A1(_12812_),
    .A2(_13154_),
    .ZN(_13859_)
  );
  INV_X1 _48702_ (
    .A(_13859_),
    .ZN(_13860_)
  );
  AND2_X1 _48703_ (
    .A1(\cpuregs[16] [19]),
    .A2(_12813_),
    .ZN(_13861_)
  );
  INV_X1 _48704_ (
    .A(_13861_),
    .ZN(_13862_)
  );
  AND2_X1 _48705_ (
    .A1(_13860_),
    .A2(_13862_),
    .ZN(_13863_)
  );
  INV_X1 _48706_ (
    .A(_13863_),
    .ZN(_00670_)
  );
  AND2_X1 _48707_ (
    .A1(_12812_),
    .A2(_13169_),
    .ZN(_13864_)
  );
  INV_X1 _48708_ (
    .A(_13864_),
    .ZN(_13865_)
  );
  AND2_X1 _48709_ (
    .A1(\cpuregs[16] [20]),
    .A2(_12813_),
    .ZN(_13866_)
  );
  INV_X1 _48710_ (
    .A(_13866_),
    .ZN(_13867_)
  );
  AND2_X1 _48711_ (
    .A1(_13865_),
    .A2(_13867_),
    .ZN(_13868_)
  );
  INV_X1 _48712_ (
    .A(_13868_),
    .ZN(_00671_)
  );
  AND2_X1 _48713_ (
    .A1(_12812_),
    .A2(_13184_),
    .ZN(_13869_)
  );
  INV_X1 _48714_ (
    .A(_13869_),
    .ZN(_13870_)
  );
  AND2_X1 _48715_ (
    .A1(\cpuregs[16] [21]),
    .A2(_12813_),
    .ZN(_13871_)
  );
  INV_X1 _48716_ (
    .A(_13871_),
    .ZN(_13872_)
  );
  AND2_X1 _48717_ (
    .A1(_13870_),
    .A2(_13872_),
    .ZN(_13873_)
  );
  INV_X1 _48718_ (
    .A(_13873_),
    .ZN(_00672_)
  );
  AND2_X1 _48719_ (
    .A1(_12812_),
    .A2(_13199_),
    .ZN(_13874_)
  );
  INV_X1 _48720_ (
    .A(_13874_),
    .ZN(_13875_)
  );
  AND2_X1 _48721_ (
    .A1(\cpuregs[16] [22]),
    .A2(_12813_),
    .ZN(_13876_)
  );
  INV_X1 _48722_ (
    .A(_13876_),
    .ZN(_13877_)
  );
  AND2_X1 _48723_ (
    .A1(_13875_),
    .A2(_13877_),
    .ZN(_13878_)
  );
  INV_X1 _48724_ (
    .A(_13878_),
    .ZN(_00673_)
  );
  AND2_X1 _48725_ (
    .A1(_12812_),
    .A2(_13214_),
    .ZN(_13879_)
  );
  INV_X1 _48726_ (
    .A(_13879_),
    .ZN(_13880_)
  );
  AND2_X1 _48727_ (
    .A1(\cpuregs[16] [23]),
    .A2(_12813_),
    .ZN(_13881_)
  );
  INV_X1 _48728_ (
    .A(_13881_),
    .ZN(_13882_)
  );
  AND2_X1 _48729_ (
    .A1(_13880_),
    .A2(_13882_),
    .ZN(_13883_)
  );
  INV_X1 _48730_ (
    .A(_13883_),
    .ZN(_00674_)
  );
  AND2_X1 _48731_ (
    .A1(_12812_),
    .A2(_13229_),
    .ZN(_13884_)
  );
  INV_X1 _48732_ (
    .A(_13884_),
    .ZN(_13885_)
  );
  AND2_X1 _48733_ (
    .A1(\cpuregs[16] [24]),
    .A2(_12813_),
    .ZN(_13886_)
  );
  INV_X1 _48734_ (
    .A(_13886_),
    .ZN(_13887_)
  );
  AND2_X1 _48735_ (
    .A1(_13885_),
    .A2(_13887_),
    .ZN(_13888_)
  );
  INV_X1 _48736_ (
    .A(_13888_),
    .ZN(_00675_)
  );
  AND2_X1 _48737_ (
    .A1(_12812_),
    .A2(_13244_),
    .ZN(_13889_)
  );
  INV_X1 _48738_ (
    .A(_13889_),
    .ZN(_13890_)
  );
  AND2_X1 _48739_ (
    .A1(\cpuregs[16] [25]),
    .A2(_12813_),
    .ZN(_13891_)
  );
  INV_X1 _48740_ (
    .A(_13891_),
    .ZN(_13892_)
  );
  AND2_X1 _48741_ (
    .A1(_13890_),
    .A2(_13892_),
    .ZN(_13893_)
  );
  INV_X1 _48742_ (
    .A(_13893_),
    .ZN(_00676_)
  );
  AND2_X1 _48743_ (
    .A1(_12812_),
    .A2(_13259_),
    .ZN(_13894_)
  );
  INV_X1 _48744_ (
    .A(_13894_),
    .ZN(_13895_)
  );
  AND2_X1 _48745_ (
    .A1(\cpuregs[16] [26]),
    .A2(_12813_),
    .ZN(_13896_)
  );
  INV_X1 _48746_ (
    .A(_13896_),
    .ZN(_13897_)
  );
  AND2_X1 _48747_ (
    .A1(_13895_),
    .A2(_13897_),
    .ZN(_13898_)
  );
  INV_X1 _48748_ (
    .A(_13898_),
    .ZN(_00677_)
  );
  AND2_X1 _48749_ (
    .A1(_12812_),
    .A2(_13274_),
    .ZN(_13899_)
  );
  INV_X1 _48750_ (
    .A(_13899_),
    .ZN(_13900_)
  );
  AND2_X1 _48751_ (
    .A1(\cpuregs[16] [27]),
    .A2(_12813_),
    .ZN(_13901_)
  );
  INV_X1 _48752_ (
    .A(_13901_),
    .ZN(_13902_)
  );
  AND2_X1 _48753_ (
    .A1(_13900_),
    .A2(_13902_),
    .ZN(_13903_)
  );
  INV_X1 _48754_ (
    .A(_13903_),
    .ZN(_00678_)
  );
  AND2_X1 _48755_ (
    .A1(_12812_),
    .A2(_13289_),
    .ZN(_13904_)
  );
  INV_X1 _48756_ (
    .A(_13904_),
    .ZN(_13905_)
  );
  AND2_X1 _48757_ (
    .A1(\cpuregs[16] [28]),
    .A2(_12813_),
    .ZN(_13906_)
  );
  INV_X1 _48758_ (
    .A(_13906_),
    .ZN(_13907_)
  );
  AND2_X1 _48759_ (
    .A1(_13905_),
    .A2(_13907_),
    .ZN(_13908_)
  );
  INV_X1 _48760_ (
    .A(_13908_),
    .ZN(_00679_)
  );
  AND2_X1 _48761_ (
    .A1(_12812_),
    .A2(_13304_),
    .ZN(_13909_)
  );
  INV_X1 _48762_ (
    .A(_13909_),
    .ZN(_13910_)
  );
  AND2_X1 _48763_ (
    .A1(\cpuregs[16] [29]),
    .A2(_12813_),
    .ZN(_13911_)
  );
  INV_X1 _48764_ (
    .A(_13911_),
    .ZN(_13912_)
  );
  AND2_X1 _48765_ (
    .A1(_13910_),
    .A2(_13912_),
    .ZN(_13913_)
  );
  INV_X1 _48766_ (
    .A(_13913_),
    .ZN(_00680_)
  );
  AND2_X1 _48767_ (
    .A1(_12812_),
    .A2(_13319_),
    .ZN(_13914_)
  );
  INV_X1 _48768_ (
    .A(_13914_),
    .ZN(_13915_)
  );
  AND2_X1 _48769_ (
    .A1(\cpuregs[16] [30]),
    .A2(_12813_),
    .ZN(_13916_)
  );
  INV_X1 _48770_ (
    .A(_13916_),
    .ZN(_13917_)
  );
  AND2_X1 _48771_ (
    .A1(_13915_),
    .A2(_13917_),
    .ZN(_13918_)
  );
  INV_X1 _48772_ (
    .A(_13918_),
    .ZN(_00681_)
  );
  AND2_X1 _48773_ (
    .A1(_12805_),
    .A2(_12874_),
    .ZN(_13919_)
  );
  INV_X1 _48774_ (
    .A(_13919_),
    .ZN(_13920_)
  );
  AND2_X1 _48775_ (
    .A1(\cpuregs[17] [0]),
    .A2(_12806_),
    .ZN(_13921_)
  );
  INV_X1 _48776_ (
    .A(_13921_),
    .ZN(_13922_)
  );
  AND2_X1 _48777_ (
    .A1(_13920_),
    .A2(_13922_),
    .ZN(_13923_)
  );
  INV_X1 _48778_ (
    .A(_13923_),
    .ZN(_00682_)
  );
  AND2_X1 _48779_ (
    .A1(_12805_),
    .A2(_12886_),
    .ZN(_13924_)
  );
  INV_X1 _48780_ (
    .A(_13924_),
    .ZN(_13925_)
  );
  AND2_X1 _48781_ (
    .A1(\cpuregs[17] [1]),
    .A2(_12806_),
    .ZN(_13926_)
  );
  INV_X1 _48782_ (
    .A(_13926_),
    .ZN(_13927_)
  );
  AND2_X1 _48783_ (
    .A1(_13925_),
    .A2(_13927_),
    .ZN(_13928_)
  );
  INV_X1 _48784_ (
    .A(_13928_),
    .ZN(_00683_)
  );
  AND2_X1 _48785_ (
    .A1(_12805_),
    .A2(_12900_),
    .ZN(_13929_)
  );
  INV_X1 _48786_ (
    .A(_13929_),
    .ZN(_13930_)
  );
  AND2_X1 _48787_ (
    .A1(\cpuregs[17] [2]),
    .A2(_12806_),
    .ZN(_13931_)
  );
  INV_X1 _48788_ (
    .A(_13931_),
    .ZN(_13932_)
  );
  AND2_X1 _48789_ (
    .A1(_13930_),
    .A2(_13932_),
    .ZN(_13933_)
  );
  INV_X1 _48790_ (
    .A(_13933_),
    .ZN(_00684_)
  );
  AND2_X1 _48791_ (
    .A1(_12805_),
    .A2(_12913_),
    .ZN(_13934_)
  );
  INV_X1 _48792_ (
    .A(_13934_),
    .ZN(_13935_)
  );
  AND2_X1 _48793_ (
    .A1(\cpuregs[17] [3]),
    .A2(_12806_),
    .ZN(_13936_)
  );
  INV_X1 _48794_ (
    .A(_13936_),
    .ZN(_13937_)
  );
  AND2_X1 _48795_ (
    .A1(_13935_),
    .A2(_13937_),
    .ZN(_13938_)
  );
  INV_X1 _48796_ (
    .A(_13938_),
    .ZN(_00685_)
  );
  AND2_X1 _48797_ (
    .A1(\cpuregs[17] [4]),
    .A2(_12806_),
    .ZN(_13939_)
  );
  INV_X1 _48798_ (
    .A(_13939_),
    .ZN(_13940_)
  );
  AND2_X1 _48799_ (
    .A1(_12805_),
    .A2(_12928_),
    .ZN(_13941_)
  );
  INV_X1 _48800_ (
    .A(_13941_),
    .ZN(_13942_)
  );
  AND2_X1 _48801_ (
    .A1(_13940_),
    .A2(_13942_),
    .ZN(_13943_)
  );
  INV_X1 _48802_ (
    .A(_13943_),
    .ZN(_00686_)
  );
  AND2_X1 _48803_ (
    .A1(_12805_),
    .A2(_12943_),
    .ZN(_13944_)
  );
  INV_X1 _48804_ (
    .A(_13944_),
    .ZN(_13945_)
  );
  AND2_X1 _48805_ (
    .A1(\cpuregs[17] [5]),
    .A2(_12806_),
    .ZN(_13946_)
  );
  INV_X1 _48806_ (
    .A(_13946_),
    .ZN(_13947_)
  );
  AND2_X1 _48807_ (
    .A1(_13945_),
    .A2(_13947_),
    .ZN(_13948_)
  );
  INV_X1 _48808_ (
    .A(_13948_),
    .ZN(_00687_)
  );
  AND2_X1 _48809_ (
    .A1(_12805_),
    .A2(_12958_),
    .ZN(_13949_)
  );
  INV_X1 _48810_ (
    .A(_13949_),
    .ZN(_13950_)
  );
  AND2_X1 _48811_ (
    .A1(\cpuregs[17] [6]),
    .A2(_12806_),
    .ZN(_13951_)
  );
  INV_X1 _48812_ (
    .A(_13951_),
    .ZN(_13952_)
  );
  AND2_X1 _48813_ (
    .A1(_13950_),
    .A2(_13952_),
    .ZN(_13953_)
  );
  INV_X1 _48814_ (
    .A(_13953_),
    .ZN(_00688_)
  );
  AND2_X1 _48815_ (
    .A1(_12805_),
    .A2(_12973_),
    .ZN(_13954_)
  );
  INV_X1 _48816_ (
    .A(_13954_),
    .ZN(_13955_)
  );
  AND2_X1 _48817_ (
    .A1(\cpuregs[17] [7]),
    .A2(_12806_),
    .ZN(_13956_)
  );
  INV_X1 _48818_ (
    .A(_13956_),
    .ZN(_13957_)
  );
  AND2_X1 _48819_ (
    .A1(_13955_),
    .A2(_13957_),
    .ZN(_13958_)
  );
  INV_X1 _48820_ (
    .A(_13958_),
    .ZN(_00689_)
  );
  AND2_X1 _48821_ (
    .A1(_12805_),
    .A2(_12988_),
    .ZN(_13959_)
  );
  INV_X1 _48822_ (
    .A(_13959_),
    .ZN(_13960_)
  );
  AND2_X1 _48823_ (
    .A1(\cpuregs[17] [8]),
    .A2(_12806_),
    .ZN(_13961_)
  );
  INV_X1 _48824_ (
    .A(_13961_),
    .ZN(_13962_)
  );
  AND2_X1 _48825_ (
    .A1(_13960_),
    .A2(_13962_),
    .ZN(_13963_)
  );
  INV_X1 _48826_ (
    .A(_13963_),
    .ZN(_00690_)
  );
  AND2_X1 _48827_ (
    .A1(_12805_),
    .A2(_13003_),
    .ZN(_13964_)
  );
  INV_X1 _48828_ (
    .A(_13964_),
    .ZN(_13965_)
  );
  AND2_X1 _48829_ (
    .A1(\cpuregs[17] [9]),
    .A2(_12806_),
    .ZN(_13966_)
  );
  INV_X1 _48830_ (
    .A(_13966_),
    .ZN(_13967_)
  );
  AND2_X1 _48831_ (
    .A1(_13965_),
    .A2(_13967_),
    .ZN(_13968_)
  );
  INV_X1 _48832_ (
    .A(_13968_),
    .ZN(_00691_)
  );
  AND2_X1 _48833_ (
    .A1(_12805_),
    .A2(_13018_),
    .ZN(_13969_)
  );
  INV_X1 _48834_ (
    .A(_13969_),
    .ZN(_13970_)
  );
  AND2_X1 _48835_ (
    .A1(\cpuregs[17] [10]),
    .A2(_12806_),
    .ZN(_13971_)
  );
  INV_X1 _48836_ (
    .A(_13971_),
    .ZN(_13972_)
  );
  AND2_X1 _48837_ (
    .A1(_13970_),
    .A2(_13972_),
    .ZN(_13973_)
  );
  INV_X1 _48838_ (
    .A(_13973_),
    .ZN(_00692_)
  );
  AND2_X1 _48839_ (
    .A1(_12805_),
    .A2(_13033_),
    .ZN(_13974_)
  );
  INV_X1 _48840_ (
    .A(_13974_),
    .ZN(_13975_)
  );
  AND2_X1 _48841_ (
    .A1(\cpuregs[17] [11]),
    .A2(_12806_),
    .ZN(_13976_)
  );
  INV_X1 _48842_ (
    .A(_13976_),
    .ZN(_13977_)
  );
  AND2_X1 _48843_ (
    .A1(_13975_),
    .A2(_13977_),
    .ZN(_13978_)
  );
  INV_X1 _48844_ (
    .A(_13978_),
    .ZN(_00693_)
  );
  AND2_X1 _48845_ (
    .A1(_12805_),
    .A2(_13048_),
    .ZN(_13979_)
  );
  INV_X1 _48846_ (
    .A(_13979_),
    .ZN(_13980_)
  );
  AND2_X1 _48847_ (
    .A1(\cpuregs[17] [12]),
    .A2(_12806_),
    .ZN(_13981_)
  );
  INV_X1 _48848_ (
    .A(_13981_),
    .ZN(_13982_)
  );
  AND2_X1 _48849_ (
    .A1(_13980_),
    .A2(_13982_),
    .ZN(_13983_)
  );
  INV_X1 _48850_ (
    .A(_13983_),
    .ZN(_00694_)
  );
  AND2_X1 _48851_ (
    .A1(_12805_),
    .A2(_13063_),
    .ZN(_13984_)
  );
  INV_X1 _48852_ (
    .A(_13984_),
    .ZN(_13985_)
  );
  AND2_X1 _48853_ (
    .A1(\cpuregs[17] [13]),
    .A2(_12806_),
    .ZN(_13986_)
  );
  INV_X1 _48854_ (
    .A(_13986_),
    .ZN(_13987_)
  );
  AND2_X1 _48855_ (
    .A1(_13985_),
    .A2(_13987_),
    .ZN(_13988_)
  );
  INV_X1 _48856_ (
    .A(_13988_),
    .ZN(_00695_)
  );
  AND2_X1 _48857_ (
    .A1(_12805_),
    .A2(_13078_),
    .ZN(_13989_)
  );
  INV_X1 _48858_ (
    .A(_13989_),
    .ZN(_13990_)
  );
  AND2_X1 _48859_ (
    .A1(\cpuregs[17] [14]),
    .A2(_12806_),
    .ZN(_13991_)
  );
  INV_X1 _48860_ (
    .A(_13991_),
    .ZN(_13992_)
  );
  AND2_X1 _48861_ (
    .A1(_13990_),
    .A2(_13992_),
    .ZN(_13993_)
  );
  INV_X1 _48862_ (
    .A(_13993_),
    .ZN(_00696_)
  );
  AND2_X1 _48863_ (
    .A1(_12805_),
    .A2(_13093_),
    .ZN(_13994_)
  );
  INV_X1 _48864_ (
    .A(_13994_),
    .ZN(_13995_)
  );
  AND2_X1 _48865_ (
    .A1(\cpuregs[17] [15]),
    .A2(_12806_),
    .ZN(_13996_)
  );
  INV_X1 _48866_ (
    .A(_13996_),
    .ZN(_13997_)
  );
  AND2_X1 _48867_ (
    .A1(_13995_),
    .A2(_13997_),
    .ZN(_13998_)
  );
  INV_X1 _48868_ (
    .A(_13998_),
    .ZN(_00697_)
  );
  AND2_X1 _48869_ (
    .A1(_12805_),
    .A2(_13108_),
    .ZN(_13999_)
  );
  INV_X1 _48870_ (
    .A(_13999_),
    .ZN(_14000_)
  );
  AND2_X1 _48871_ (
    .A1(\cpuregs[17] [16]),
    .A2(_12806_),
    .ZN(_14001_)
  );
  INV_X1 _48872_ (
    .A(_14001_),
    .ZN(_14002_)
  );
  AND2_X1 _48873_ (
    .A1(_14000_),
    .A2(_14002_),
    .ZN(_14003_)
  );
  INV_X1 _48874_ (
    .A(_14003_),
    .ZN(_00698_)
  );
  AND2_X1 _48875_ (
    .A1(_12805_),
    .A2(_13123_),
    .ZN(_14004_)
  );
  INV_X1 _48876_ (
    .A(_14004_),
    .ZN(_14005_)
  );
  AND2_X1 _48877_ (
    .A1(\cpuregs[17] [17]),
    .A2(_12806_),
    .ZN(_14006_)
  );
  INV_X1 _48878_ (
    .A(_14006_),
    .ZN(_14007_)
  );
  AND2_X1 _48879_ (
    .A1(_14005_),
    .A2(_14007_),
    .ZN(_14008_)
  );
  INV_X1 _48880_ (
    .A(_14008_),
    .ZN(_00699_)
  );
  AND2_X1 _48881_ (
    .A1(_12805_),
    .A2(_13139_),
    .ZN(_14009_)
  );
  INV_X1 _48882_ (
    .A(_14009_),
    .ZN(_14010_)
  );
  AND2_X1 _48883_ (
    .A1(\cpuregs[17] [18]),
    .A2(_12806_),
    .ZN(_14011_)
  );
  INV_X1 _48884_ (
    .A(_14011_),
    .ZN(_14012_)
  );
  AND2_X1 _48885_ (
    .A1(_14010_),
    .A2(_14012_),
    .ZN(_14013_)
  );
  INV_X1 _48886_ (
    .A(_14013_),
    .ZN(_00700_)
  );
  AND2_X1 _48887_ (
    .A1(_12805_),
    .A2(_13154_),
    .ZN(_14014_)
  );
  INV_X1 _48888_ (
    .A(_14014_),
    .ZN(_14015_)
  );
  AND2_X1 _48889_ (
    .A1(\cpuregs[17] [19]),
    .A2(_12806_),
    .ZN(_14016_)
  );
  INV_X1 _48890_ (
    .A(_14016_),
    .ZN(_14017_)
  );
  AND2_X1 _48891_ (
    .A1(_14015_),
    .A2(_14017_),
    .ZN(_14018_)
  );
  INV_X1 _48892_ (
    .A(_14018_),
    .ZN(_00701_)
  );
  AND2_X1 _48893_ (
    .A1(_12805_),
    .A2(_13169_),
    .ZN(_14019_)
  );
  INV_X1 _48894_ (
    .A(_14019_),
    .ZN(_14020_)
  );
  AND2_X1 _48895_ (
    .A1(\cpuregs[17] [20]),
    .A2(_12806_),
    .ZN(_14021_)
  );
  INV_X1 _48896_ (
    .A(_14021_),
    .ZN(_14022_)
  );
  AND2_X1 _48897_ (
    .A1(_14020_),
    .A2(_14022_),
    .ZN(_14023_)
  );
  INV_X1 _48898_ (
    .A(_14023_),
    .ZN(_00702_)
  );
  AND2_X1 _48899_ (
    .A1(_12805_),
    .A2(_13184_),
    .ZN(_14024_)
  );
  INV_X1 _48900_ (
    .A(_14024_),
    .ZN(_14025_)
  );
  AND2_X1 _48901_ (
    .A1(\cpuregs[17] [21]),
    .A2(_12806_),
    .ZN(_14026_)
  );
  INV_X1 _48902_ (
    .A(_14026_),
    .ZN(_14027_)
  );
  AND2_X1 _48903_ (
    .A1(_14025_),
    .A2(_14027_),
    .ZN(_14028_)
  );
  INV_X1 _48904_ (
    .A(_14028_),
    .ZN(_00703_)
  );
  AND2_X1 _48905_ (
    .A1(_12805_),
    .A2(_13199_),
    .ZN(_14029_)
  );
  INV_X1 _48906_ (
    .A(_14029_),
    .ZN(_14030_)
  );
  AND2_X1 _48907_ (
    .A1(\cpuregs[17] [22]),
    .A2(_12806_),
    .ZN(_14031_)
  );
  INV_X1 _48908_ (
    .A(_14031_),
    .ZN(_14032_)
  );
  AND2_X1 _48909_ (
    .A1(_14030_),
    .A2(_14032_),
    .ZN(_14033_)
  );
  INV_X1 _48910_ (
    .A(_14033_),
    .ZN(_00704_)
  );
  AND2_X1 _48911_ (
    .A1(_12805_),
    .A2(_13214_),
    .ZN(_14034_)
  );
  INV_X1 _48912_ (
    .A(_14034_),
    .ZN(_14035_)
  );
  AND2_X1 _48913_ (
    .A1(\cpuregs[17] [23]),
    .A2(_12806_),
    .ZN(_14036_)
  );
  INV_X1 _48914_ (
    .A(_14036_),
    .ZN(_14037_)
  );
  AND2_X1 _48915_ (
    .A1(_14035_),
    .A2(_14037_),
    .ZN(_14038_)
  );
  INV_X1 _48916_ (
    .A(_14038_),
    .ZN(_00705_)
  );
  AND2_X1 _48917_ (
    .A1(_12805_),
    .A2(_13229_),
    .ZN(_14039_)
  );
  INV_X1 _48918_ (
    .A(_14039_),
    .ZN(_14040_)
  );
  AND2_X1 _48919_ (
    .A1(\cpuregs[17] [24]),
    .A2(_12806_),
    .ZN(_14041_)
  );
  INV_X1 _48920_ (
    .A(_14041_),
    .ZN(_14042_)
  );
  AND2_X1 _48921_ (
    .A1(_14040_),
    .A2(_14042_),
    .ZN(_14043_)
  );
  INV_X1 _48922_ (
    .A(_14043_),
    .ZN(_00706_)
  );
  AND2_X1 _48923_ (
    .A1(_12805_),
    .A2(_13244_),
    .ZN(_14044_)
  );
  INV_X1 _48924_ (
    .A(_14044_),
    .ZN(_14045_)
  );
  AND2_X1 _48925_ (
    .A1(\cpuregs[17] [25]),
    .A2(_12806_),
    .ZN(_14046_)
  );
  INV_X1 _48926_ (
    .A(_14046_),
    .ZN(_14047_)
  );
  AND2_X1 _48927_ (
    .A1(_14045_),
    .A2(_14047_),
    .ZN(_14048_)
  );
  INV_X1 _48928_ (
    .A(_14048_),
    .ZN(_00707_)
  );
  AND2_X1 _48929_ (
    .A1(_12805_),
    .A2(_13259_),
    .ZN(_14049_)
  );
  INV_X1 _48930_ (
    .A(_14049_),
    .ZN(_14050_)
  );
  AND2_X1 _48931_ (
    .A1(\cpuregs[17] [26]),
    .A2(_12806_),
    .ZN(_14051_)
  );
  INV_X1 _48932_ (
    .A(_14051_),
    .ZN(_14052_)
  );
  AND2_X1 _48933_ (
    .A1(_14050_),
    .A2(_14052_),
    .ZN(_14053_)
  );
  INV_X1 _48934_ (
    .A(_14053_),
    .ZN(_00708_)
  );
  AND2_X1 _48935_ (
    .A1(_12805_),
    .A2(_13274_),
    .ZN(_14054_)
  );
  INV_X1 _48936_ (
    .A(_14054_),
    .ZN(_14055_)
  );
  AND2_X1 _48937_ (
    .A1(\cpuregs[17] [27]),
    .A2(_12806_),
    .ZN(_14056_)
  );
  INV_X1 _48938_ (
    .A(_14056_),
    .ZN(_14057_)
  );
  AND2_X1 _48939_ (
    .A1(_14055_),
    .A2(_14057_),
    .ZN(_14058_)
  );
  INV_X1 _48940_ (
    .A(_14058_),
    .ZN(_00709_)
  );
  AND2_X1 _48941_ (
    .A1(_12805_),
    .A2(_13289_),
    .ZN(_14059_)
  );
  INV_X1 _48942_ (
    .A(_14059_),
    .ZN(_14060_)
  );
  AND2_X1 _48943_ (
    .A1(\cpuregs[17] [28]),
    .A2(_12806_),
    .ZN(_14061_)
  );
  INV_X1 _48944_ (
    .A(_14061_),
    .ZN(_14062_)
  );
  AND2_X1 _48945_ (
    .A1(_14060_),
    .A2(_14062_),
    .ZN(_14063_)
  );
  INV_X1 _48946_ (
    .A(_14063_),
    .ZN(_00710_)
  );
  AND2_X1 _48947_ (
    .A1(_12805_),
    .A2(_13304_),
    .ZN(_14064_)
  );
  INV_X1 _48948_ (
    .A(_14064_),
    .ZN(_14065_)
  );
  AND2_X1 _48949_ (
    .A1(\cpuregs[17] [29]),
    .A2(_12806_),
    .ZN(_14066_)
  );
  INV_X1 _48950_ (
    .A(_14066_),
    .ZN(_14067_)
  );
  AND2_X1 _48951_ (
    .A1(_14065_),
    .A2(_14067_),
    .ZN(_14068_)
  );
  INV_X1 _48952_ (
    .A(_14068_),
    .ZN(_00711_)
  );
  AND2_X1 _48953_ (
    .A1(_12805_),
    .A2(_13319_),
    .ZN(_14069_)
  );
  INV_X1 _48954_ (
    .A(_14069_),
    .ZN(_14070_)
  );
  AND2_X1 _48955_ (
    .A1(\cpuregs[17] [30]),
    .A2(_12806_),
    .ZN(_14071_)
  );
  INV_X1 _48956_ (
    .A(_14071_),
    .ZN(_14072_)
  );
  AND2_X1 _48957_ (
    .A1(_14070_),
    .A2(_14072_),
    .ZN(_14073_)
  );
  INV_X1 _48958_ (
    .A(_14073_),
    .ZN(_00712_)
  );
  AND2_X1 _48959_ (
    .A1(_12842_),
    .A2(_12874_),
    .ZN(_14074_)
  );
  INV_X1 _48960_ (
    .A(_14074_),
    .ZN(_14075_)
  );
  AND2_X1 _48961_ (
    .A1(\cpuregs[12] [0]),
    .A2(_12843_),
    .ZN(_14076_)
  );
  INV_X1 _48962_ (
    .A(_14076_),
    .ZN(_14077_)
  );
  AND2_X1 _48963_ (
    .A1(_14075_),
    .A2(_14077_),
    .ZN(_14078_)
  );
  INV_X1 _48964_ (
    .A(_14078_),
    .ZN(_00713_)
  );
  AND2_X1 _48965_ (
    .A1(_12842_),
    .A2(_12886_),
    .ZN(_14079_)
  );
  INV_X1 _48966_ (
    .A(_14079_),
    .ZN(_14080_)
  );
  AND2_X1 _48967_ (
    .A1(\cpuregs[12] [1]),
    .A2(_12843_),
    .ZN(_14081_)
  );
  INV_X1 _48968_ (
    .A(_14081_),
    .ZN(_14082_)
  );
  AND2_X1 _48969_ (
    .A1(_14080_),
    .A2(_14082_),
    .ZN(_14083_)
  );
  INV_X1 _48970_ (
    .A(_14083_),
    .ZN(_00714_)
  );
  AND2_X1 _48971_ (
    .A1(\cpuregs[12] [2]),
    .A2(_12843_),
    .ZN(_14084_)
  );
  INV_X1 _48972_ (
    .A(_14084_),
    .ZN(_14085_)
  );
  AND2_X1 _48973_ (
    .A1(_12842_),
    .A2(_12900_),
    .ZN(_14086_)
  );
  INV_X1 _48974_ (
    .A(_14086_),
    .ZN(_14087_)
  );
  AND2_X1 _48975_ (
    .A1(_14085_),
    .A2(_14087_),
    .ZN(_14088_)
  );
  INV_X1 _48976_ (
    .A(_14088_),
    .ZN(_00715_)
  );
  AND2_X1 _48977_ (
    .A1(_12842_),
    .A2(_12913_),
    .ZN(_14089_)
  );
  INV_X1 _48978_ (
    .A(_14089_),
    .ZN(_14090_)
  );
  AND2_X1 _48979_ (
    .A1(\cpuregs[12] [3]),
    .A2(_12843_),
    .ZN(_14091_)
  );
  INV_X1 _48980_ (
    .A(_14091_),
    .ZN(_14092_)
  );
  AND2_X1 _48981_ (
    .A1(_14090_),
    .A2(_14092_),
    .ZN(_14093_)
  );
  INV_X1 _48982_ (
    .A(_14093_),
    .ZN(_00716_)
  );
  AND2_X1 _48983_ (
    .A1(\cpuregs[12] [4]),
    .A2(_12843_),
    .ZN(_14094_)
  );
  INV_X1 _48984_ (
    .A(_14094_),
    .ZN(_14095_)
  );
  AND2_X1 _48985_ (
    .A1(_12842_),
    .A2(_12928_),
    .ZN(_14096_)
  );
  INV_X1 _48986_ (
    .A(_14096_),
    .ZN(_14097_)
  );
  AND2_X1 _48987_ (
    .A1(_14095_),
    .A2(_14097_),
    .ZN(_14098_)
  );
  INV_X1 _48988_ (
    .A(_14098_),
    .ZN(_00717_)
  );
  AND2_X1 _48989_ (
    .A1(_12842_),
    .A2(_12943_),
    .ZN(_14099_)
  );
  INV_X1 _48990_ (
    .A(_14099_),
    .ZN(_14100_)
  );
  AND2_X1 _48991_ (
    .A1(\cpuregs[12] [5]),
    .A2(_12843_),
    .ZN(_14101_)
  );
  INV_X1 _48992_ (
    .A(_14101_),
    .ZN(_14102_)
  );
  AND2_X1 _48993_ (
    .A1(_14100_),
    .A2(_14102_),
    .ZN(_14103_)
  );
  INV_X1 _48994_ (
    .A(_14103_),
    .ZN(_00718_)
  );
  AND2_X1 _48995_ (
    .A1(_12842_),
    .A2(_12958_),
    .ZN(_14104_)
  );
  INV_X1 _48996_ (
    .A(_14104_),
    .ZN(_14105_)
  );
  AND2_X1 _48997_ (
    .A1(\cpuregs[12] [6]),
    .A2(_12843_),
    .ZN(_14106_)
  );
  INV_X1 _48998_ (
    .A(_14106_),
    .ZN(_14107_)
  );
  AND2_X1 _48999_ (
    .A1(_14105_),
    .A2(_14107_),
    .ZN(_14108_)
  );
  INV_X1 _49000_ (
    .A(_14108_),
    .ZN(_00719_)
  );
  AND2_X1 _49001_ (
    .A1(_12842_),
    .A2(_12973_),
    .ZN(_14109_)
  );
  INV_X1 _49002_ (
    .A(_14109_),
    .ZN(_14110_)
  );
  AND2_X1 _49003_ (
    .A1(\cpuregs[12] [7]),
    .A2(_12843_),
    .ZN(_14111_)
  );
  INV_X1 _49004_ (
    .A(_14111_),
    .ZN(_14112_)
  );
  AND2_X1 _49005_ (
    .A1(_14110_),
    .A2(_14112_),
    .ZN(_14113_)
  );
  INV_X1 _49006_ (
    .A(_14113_),
    .ZN(_00720_)
  );
  AND2_X1 _49007_ (
    .A1(_12842_),
    .A2(_12988_),
    .ZN(_14114_)
  );
  INV_X1 _49008_ (
    .A(_14114_),
    .ZN(_14115_)
  );
  AND2_X1 _49009_ (
    .A1(\cpuregs[12] [8]),
    .A2(_12843_),
    .ZN(_14116_)
  );
  INV_X1 _49010_ (
    .A(_14116_),
    .ZN(_14117_)
  );
  AND2_X1 _49011_ (
    .A1(_14115_),
    .A2(_14117_),
    .ZN(_14118_)
  );
  INV_X1 _49012_ (
    .A(_14118_),
    .ZN(_00721_)
  );
  AND2_X1 _49013_ (
    .A1(_12842_),
    .A2(_13003_),
    .ZN(_14119_)
  );
  INV_X1 _49014_ (
    .A(_14119_),
    .ZN(_14120_)
  );
  AND2_X1 _49015_ (
    .A1(\cpuregs[12] [9]),
    .A2(_12843_),
    .ZN(_14121_)
  );
  INV_X1 _49016_ (
    .A(_14121_),
    .ZN(_14122_)
  );
  AND2_X1 _49017_ (
    .A1(_14120_),
    .A2(_14122_),
    .ZN(_14123_)
  );
  INV_X1 _49018_ (
    .A(_14123_),
    .ZN(_00722_)
  );
  AND2_X1 _49019_ (
    .A1(_12842_),
    .A2(_13018_),
    .ZN(_14124_)
  );
  INV_X1 _49020_ (
    .A(_14124_),
    .ZN(_14125_)
  );
  AND2_X1 _49021_ (
    .A1(\cpuregs[12] [10]),
    .A2(_12843_),
    .ZN(_14126_)
  );
  INV_X1 _49022_ (
    .A(_14126_),
    .ZN(_14127_)
  );
  AND2_X1 _49023_ (
    .A1(_14125_),
    .A2(_14127_),
    .ZN(_14128_)
  );
  INV_X1 _49024_ (
    .A(_14128_),
    .ZN(_00723_)
  );
  AND2_X1 _49025_ (
    .A1(_12842_),
    .A2(_13033_),
    .ZN(_14129_)
  );
  INV_X1 _49026_ (
    .A(_14129_),
    .ZN(_14130_)
  );
  AND2_X1 _49027_ (
    .A1(\cpuregs[12] [11]),
    .A2(_12843_),
    .ZN(_14131_)
  );
  INV_X1 _49028_ (
    .A(_14131_),
    .ZN(_14132_)
  );
  AND2_X1 _49029_ (
    .A1(_14130_),
    .A2(_14132_),
    .ZN(_14133_)
  );
  INV_X1 _49030_ (
    .A(_14133_),
    .ZN(_00724_)
  );
  AND2_X1 _49031_ (
    .A1(_12842_),
    .A2(_13048_),
    .ZN(_14134_)
  );
  INV_X1 _49032_ (
    .A(_14134_),
    .ZN(_14135_)
  );
  AND2_X1 _49033_ (
    .A1(\cpuregs[12] [12]),
    .A2(_12843_),
    .ZN(_14136_)
  );
  INV_X1 _49034_ (
    .A(_14136_),
    .ZN(_14137_)
  );
  AND2_X1 _49035_ (
    .A1(_14135_),
    .A2(_14137_),
    .ZN(_14138_)
  );
  INV_X1 _49036_ (
    .A(_14138_),
    .ZN(_00725_)
  );
  AND2_X1 _49037_ (
    .A1(_12842_),
    .A2(_13063_),
    .ZN(_14139_)
  );
  INV_X1 _49038_ (
    .A(_14139_),
    .ZN(_14140_)
  );
  AND2_X1 _49039_ (
    .A1(\cpuregs[12] [13]),
    .A2(_12843_),
    .ZN(_14141_)
  );
  INV_X1 _49040_ (
    .A(_14141_),
    .ZN(_14142_)
  );
  AND2_X1 _49041_ (
    .A1(_14140_),
    .A2(_14142_),
    .ZN(_14143_)
  );
  INV_X1 _49042_ (
    .A(_14143_),
    .ZN(_00726_)
  );
  AND2_X1 _49043_ (
    .A1(_12842_),
    .A2(_13078_),
    .ZN(_14144_)
  );
  INV_X1 _49044_ (
    .A(_14144_),
    .ZN(_14145_)
  );
  AND2_X1 _49045_ (
    .A1(\cpuregs[12] [14]),
    .A2(_12843_),
    .ZN(_14146_)
  );
  INV_X1 _49046_ (
    .A(_14146_),
    .ZN(_14147_)
  );
  AND2_X1 _49047_ (
    .A1(_14145_),
    .A2(_14147_),
    .ZN(_14148_)
  );
  INV_X1 _49048_ (
    .A(_14148_),
    .ZN(_00727_)
  );
  AND2_X1 _49049_ (
    .A1(_12842_),
    .A2(_13093_),
    .ZN(_14149_)
  );
  INV_X1 _49050_ (
    .A(_14149_),
    .ZN(_14150_)
  );
  AND2_X1 _49051_ (
    .A1(\cpuregs[12] [15]),
    .A2(_12843_),
    .ZN(_14151_)
  );
  INV_X1 _49052_ (
    .A(_14151_),
    .ZN(_14152_)
  );
  AND2_X1 _49053_ (
    .A1(_14150_),
    .A2(_14152_),
    .ZN(_14153_)
  );
  INV_X1 _49054_ (
    .A(_14153_),
    .ZN(_00728_)
  );
  AND2_X1 _49055_ (
    .A1(_12842_),
    .A2(_13108_),
    .ZN(_14154_)
  );
  INV_X1 _49056_ (
    .A(_14154_),
    .ZN(_14155_)
  );
  AND2_X1 _49057_ (
    .A1(\cpuregs[12] [16]),
    .A2(_12843_),
    .ZN(_14156_)
  );
  INV_X1 _49058_ (
    .A(_14156_),
    .ZN(_14157_)
  );
  AND2_X1 _49059_ (
    .A1(_14155_),
    .A2(_14157_),
    .ZN(_14158_)
  );
  INV_X1 _49060_ (
    .A(_14158_),
    .ZN(_00729_)
  );
  AND2_X1 _49061_ (
    .A1(\cpuregs[12] [17]),
    .A2(_12843_),
    .ZN(_14159_)
  );
  INV_X1 _49062_ (
    .A(_14159_),
    .ZN(_14160_)
  );
  AND2_X1 _49063_ (
    .A1(_12842_),
    .A2(_13123_),
    .ZN(_14161_)
  );
  INV_X1 _49064_ (
    .A(_14161_),
    .ZN(_14162_)
  );
  AND2_X1 _49065_ (
    .A1(_14160_),
    .A2(_14162_),
    .ZN(_14163_)
  );
  INV_X1 _49066_ (
    .A(_14163_),
    .ZN(_00730_)
  );
  AND2_X1 _49067_ (
    .A1(\cpuregs[12] [18]),
    .A2(_12843_),
    .ZN(_14164_)
  );
  INV_X1 _49068_ (
    .A(_14164_),
    .ZN(_14165_)
  );
  AND2_X1 _49069_ (
    .A1(_12842_),
    .A2(_13139_),
    .ZN(_14166_)
  );
  INV_X1 _49070_ (
    .A(_14166_),
    .ZN(_14167_)
  );
  AND2_X1 _49071_ (
    .A1(_14165_),
    .A2(_14167_),
    .ZN(_14168_)
  );
  INV_X1 _49072_ (
    .A(_14168_),
    .ZN(_00731_)
  );
  AND2_X1 _49073_ (
    .A1(\cpuregs[12] [19]),
    .A2(_12843_),
    .ZN(_14169_)
  );
  INV_X1 _49074_ (
    .A(_14169_),
    .ZN(_14170_)
  );
  AND2_X1 _49075_ (
    .A1(_12842_),
    .A2(_13154_),
    .ZN(_14171_)
  );
  INV_X1 _49076_ (
    .A(_14171_),
    .ZN(_14172_)
  );
  AND2_X1 _49077_ (
    .A1(_14170_),
    .A2(_14172_),
    .ZN(_14173_)
  );
  INV_X1 _49078_ (
    .A(_14173_),
    .ZN(_00732_)
  );
  AND2_X1 _49079_ (
    .A1(\cpuregs[12] [20]),
    .A2(_12843_),
    .ZN(_14174_)
  );
  INV_X1 _49080_ (
    .A(_14174_),
    .ZN(_14175_)
  );
  AND2_X1 _49081_ (
    .A1(_12842_),
    .A2(_13169_),
    .ZN(_14176_)
  );
  INV_X1 _49082_ (
    .A(_14176_),
    .ZN(_14177_)
  );
  AND2_X1 _49083_ (
    .A1(_14175_),
    .A2(_14177_),
    .ZN(_14178_)
  );
  INV_X1 _49084_ (
    .A(_14178_),
    .ZN(_00733_)
  );
  AND2_X1 _49085_ (
    .A1(\cpuregs[12] [21]),
    .A2(_12843_),
    .ZN(_14179_)
  );
  INV_X1 _49086_ (
    .A(_14179_),
    .ZN(_14180_)
  );
  AND2_X1 _49087_ (
    .A1(_12842_),
    .A2(_13184_),
    .ZN(_14181_)
  );
  INV_X1 _49088_ (
    .A(_14181_),
    .ZN(_14182_)
  );
  AND2_X1 _49089_ (
    .A1(_14180_),
    .A2(_14182_),
    .ZN(_14183_)
  );
  INV_X1 _49090_ (
    .A(_14183_),
    .ZN(_00734_)
  );
  AND2_X1 _49091_ (
    .A1(\cpuregs[12] [22]),
    .A2(_12843_),
    .ZN(_14184_)
  );
  INV_X1 _49092_ (
    .A(_14184_),
    .ZN(_14185_)
  );
  AND2_X1 _49093_ (
    .A1(_12842_),
    .A2(_13199_),
    .ZN(_14186_)
  );
  INV_X1 _49094_ (
    .A(_14186_),
    .ZN(_14187_)
  );
  AND2_X1 _49095_ (
    .A1(_14185_),
    .A2(_14187_),
    .ZN(_14188_)
  );
  INV_X1 _49096_ (
    .A(_14188_),
    .ZN(_00735_)
  );
  AND2_X1 _49097_ (
    .A1(\cpuregs[12] [23]),
    .A2(_12843_),
    .ZN(_14189_)
  );
  INV_X1 _49098_ (
    .A(_14189_),
    .ZN(_14190_)
  );
  AND2_X1 _49099_ (
    .A1(_12842_),
    .A2(_13214_),
    .ZN(_14191_)
  );
  INV_X1 _49100_ (
    .A(_14191_),
    .ZN(_14192_)
  );
  AND2_X1 _49101_ (
    .A1(_14190_),
    .A2(_14192_),
    .ZN(_14193_)
  );
  INV_X1 _49102_ (
    .A(_14193_),
    .ZN(_00736_)
  );
  AND2_X1 _49103_ (
    .A1(\cpuregs[12] [24]),
    .A2(_12843_),
    .ZN(_14194_)
  );
  INV_X1 _49104_ (
    .A(_14194_),
    .ZN(_14195_)
  );
  AND2_X1 _49105_ (
    .A1(_12842_),
    .A2(_13229_),
    .ZN(_14196_)
  );
  INV_X1 _49106_ (
    .A(_14196_),
    .ZN(_14197_)
  );
  AND2_X1 _49107_ (
    .A1(_14195_),
    .A2(_14197_),
    .ZN(_14198_)
  );
  INV_X1 _49108_ (
    .A(_14198_),
    .ZN(_00737_)
  );
  AND2_X1 _49109_ (
    .A1(\cpuregs[12] [25]),
    .A2(_12843_),
    .ZN(_14199_)
  );
  INV_X1 _49110_ (
    .A(_14199_),
    .ZN(_14200_)
  );
  AND2_X1 _49111_ (
    .A1(_12842_),
    .A2(_13244_),
    .ZN(_14201_)
  );
  INV_X1 _49112_ (
    .A(_14201_),
    .ZN(_14202_)
  );
  AND2_X1 _49113_ (
    .A1(_14200_),
    .A2(_14202_),
    .ZN(_14203_)
  );
  INV_X1 _49114_ (
    .A(_14203_),
    .ZN(_00738_)
  );
  AND2_X1 _49115_ (
    .A1(\cpuregs[12] [26]),
    .A2(_12843_),
    .ZN(_14204_)
  );
  INV_X1 _49116_ (
    .A(_14204_),
    .ZN(_14205_)
  );
  AND2_X1 _49117_ (
    .A1(_12842_),
    .A2(_13259_),
    .ZN(_14206_)
  );
  INV_X1 _49118_ (
    .A(_14206_),
    .ZN(_14207_)
  );
  AND2_X1 _49119_ (
    .A1(_14205_),
    .A2(_14207_),
    .ZN(_14208_)
  );
  INV_X1 _49120_ (
    .A(_14208_),
    .ZN(_00739_)
  );
  AND2_X1 _49121_ (
    .A1(\cpuregs[12] [27]),
    .A2(_12843_),
    .ZN(_14209_)
  );
  INV_X1 _49122_ (
    .A(_14209_),
    .ZN(_14210_)
  );
  AND2_X1 _49123_ (
    .A1(_12842_),
    .A2(_13274_),
    .ZN(_14211_)
  );
  INV_X1 _49124_ (
    .A(_14211_),
    .ZN(_14212_)
  );
  AND2_X1 _49125_ (
    .A1(_14210_),
    .A2(_14212_),
    .ZN(_14213_)
  );
  INV_X1 _49126_ (
    .A(_14213_),
    .ZN(_00740_)
  );
  AND2_X1 _49127_ (
    .A1(\cpuregs[12] [28]),
    .A2(_12843_),
    .ZN(_14214_)
  );
  INV_X1 _49128_ (
    .A(_14214_),
    .ZN(_14215_)
  );
  AND2_X1 _49129_ (
    .A1(_12842_),
    .A2(_13289_),
    .ZN(_14216_)
  );
  INV_X1 _49130_ (
    .A(_14216_),
    .ZN(_14217_)
  );
  AND2_X1 _49131_ (
    .A1(_14215_),
    .A2(_14217_),
    .ZN(_14218_)
  );
  INV_X1 _49132_ (
    .A(_14218_),
    .ZN(_00741_)
  );
  AND2_X1 _49133_ (
    .A1(\cpuregs[12] [29]),
    .A2(_12843_),
    .ZN(_14219_)
  );
  INV_X1 _49134_ (
    .A(_14219_),
    .ZN(_14220_)
  );
  AND2_X1 _49135_ (
    .A1(_12842_),
    .A2(_13304_),
    .ZN(_14221_)
  );
  INV_X1 _49136_ (
    .A(_14221_),
    .ZN(_14222_)
  );
  AND2_X1 _49137_ (
    .A1(_14220_),
    .A2(_14222_),
    .ZN(_14223_)
  );
  INV_X1 _49138_ (
    .A(_14223_),
    .ZN(_00742_)
  );
  AND2_X1 _49139_ (
    .A1(\cpuregs[12] [30]),
    .A2(_12843_),
    .ZN(_14224_)
  );
  INV_X1 _49140_ (
    .A(_14224_),
    .ZN(_14225_)
  );
  AND2_X1 _49141_ (
    .A1(_12842_),
    .A2(_13319_),
    .ZN(_14226_)
  );
  INV_X1 _49142_ (
    .A(_14226_),
    .ZN(_14227_)
  );
  AND2_X1 _49143_ (
    .A1(_14225_),
    .A2(_14227_),
    .ZN(_14228_)
  );
  INV_X1 _49144_ (
    .A(_14228_),
    .ZN(_00743_)
  );
  AND2_X1 _49145_ (
    .A1(_12680_),
    .A2(_12874_),
    .ZN(_14229_)
  );
  INV_X1 _49146_ (
    .A(_14229_),
    .ZN(_14230_)
  );
  AND2_X1 _49147_ (
    .A1(\cpuregs[3] [0]),
    .A2(_12681_),
    .ZN(_14231_)
  );
  INV_X1 _49148_ (
    .A(_14231_),
    .ZN(_14232_)
  );
  AND2_X1 _49149_ (
    .A1(_14230_),
    .A2(_14232_),
    .ZN(_14233_)
  );
  INV_X1 _49150_ (
    .A(_14233_),
    .ZN(_00744_)
  );
  AND2_X1 _49151_ (
    .A1(_12680_),
    .A2(_12886_),
    .ZN(_14234_)
  );
  INV_X1 _49152_ (
    .A(_14234_),
    .ZN(_14235_)
  );
  AND2_X1 _49153_ (
    .A1(\cpuregs[3] [1]),
    .A2(_12681_),
    .ZN(_14236_)
  );
  INV_X1 _49154_ (
    .A(_14236_),
    .ZN(_14237_)
  );
  AND2_X1 _49155_ (
    .A1(_14235_),
    .A2(_14237_),
    .ZN(_14238_)
  );
  INV_X1 _49156_ (
    .A(_14238_),
    .ZN(_00745_)
  );
  AND2_X1 _49157_ (
    .A1(_12680_),
    .A2(_12900_),
    .ZN(_14239_)
  );
  INV_X1 _49158_ (
    .A(_14239_),
    .ZN(_14240_)
  );
  AND2_X1 _49159_ (
    .A1(\cpuregs[3] [2]),
    .A2(_12681_),
    .ZN(_14241_)
  );
  INV_X1 _49160_ (
    .A(_14241_),
    .ZN(_14242_)
  );
  AND2_X1 _49161_ (
    .A1(_14240_),
    .A2(_14242_),
    .ZN(_14243_)
  );
  INV_X1 _49162_ (
    .A(_14243_),
    .ZN(_00746_)
  );
  AND2_X1 _49163_ (
    .A1(_12680_),
    .A2(_12913_),
    .ZN(_14244_)
  );
  INV_X1 _49164_ (
    .A(_14244_),
    .ZN(_14245_)
  );
  AND2_X1 _49165_ (
    .A1(\cpuregs[3] [3]),
    .A2(_12681_),
    .ZN(_14246_)
  );
  INV_X1 _49166_ (
    .A(_14246_),
    .ZN(_14247_)
  );
  AND2_X1 _49167_ (
    .A1(_14245_),
    .A2(_14247_),
    .ZN(_14248_)
  );
  INV_X1 _49168_ (
    .A(_14248_),
    .ZN(_00747_)
  );
  AND2_X1 _49169_ (
    .A1(_12680_),
    .A2(_12928_),
    .ZN(_14249_)
  );
  INV_X1 _49170_ (
    .A(_14249_),
    .ZN(_14250_)
  );
  AND2_X1 _49171_ (
    .A1(\cpuregs[3] [4]),
    .A2(_12681_),
    .ZN(_14251_)
  );
  INV_X1 _49172_ (
    .A(_14251_),
    .ZN(_14252_)
  );
  AND2_X1 _49173_ (
    .A1(_14250_),
    .A2(_14252_),
    .ZN(_14253_)
  );
  INV_X1 _49174_ (
    .A(_14253_),
    .ZN(_00748_)
  );
  AND2_X1 _49175_ (
    .A1(_12680_),
    .A2(_12943_),
    .ZN(_14254_)
  );
  INV_X1 _49176_ (
    .A(_14254_),
    .ZN(_14255_)
  );
  AND2_X1 _49177_ (
    .A1(\cpuregs[3] [5]),
    .A2(_12681_),
    .ZN(_14256_)
  );
  INV_X1 _49178_ (
    .A(_14256_),
    .ZN(_14257_)
  );
  AND2_X1 _49179_ (
    .A1(_14255_),
    .A2(_14257_),
    .ZN(_14258_)
  );
  INV_X1 _49180_ (
    .A(_14258_),
    .ZN(_00749_)
  );
  AND2_X1 _49181_ (
    .A1(_12680_),
    .A2(_12958_),
    .ZN(_14259_)
  );
  INV_X1 _49182_ (
    .A(_14259_),
    .ZN(_14260_)
  );
  AND2_X1 _49183_ (
    .A1(\cpuregs[3] [6]),
    .A2(_12681_),
    .ZN(_14261_)
  );
  INV_X1 _49184_ (
    .A(_14261_),
    .ZN(_14262_)
  );
  AND2_X1 _49185_ (
    .A1(_14260_),
    .A2(_14262_),
    .ZN(_14263_)
  );
  INV_X1 _49186_ (
    .A(_14263_),
    .ZN(_00750_)
  );
  AND2_X1 _49187_ (
    .A1(_12680_),
    .A2(_12973_),
    .ZN(_14264_)
  );
  INV_X1 _49188_ (
    .A(_14264_),
    .ZN(_14265_)
  );
  AND2_X1 _49189_ (
    .A1(\cpuregs[3] [7]),
    .A2(_12681_),
    .ZN(_14266_)
  );
  INV_X1 _49190_ (
    .A(_14266_),
    .ZN(_14267_)
  );
  AND2_X1 _49191_ (
    .A1(_14265_),
    .A2(_14267_),
    .ZN(_14268_)
  );
  INV_X1 _49192_ (
    .A(_14268_),
    .ZN(_00751_)
  );
  AND2_X1 _49193_ (
    .A1(_12680_),
    .A2(_12988_),
    .ZN(_14269_)
  );
  INV_X1 _49194_ (
    .A(_14269_),
    .ZN(_14270_)
  );
  AND2_X1 _49195_ (
    .A1(\cpuregs[3] [8]),
    .A2(_12681_),
    .ZN(_14271_)
  );
  INV_X1 _49196_ (
    .A(_14271_),
    .ZN(_14272_)
  );
  AND2_X1 _49197_ (
    .A1(_14270_),
    .A2(_14272_),
    .ZN(_14273_)
  );
  INV_X1 _49198_ (
    .A(_14273_),
    .ZN(_00752_)
  );
  AND2_X1 _49199_ (
    .A1(_12680_),
    .A2(_13003_),
    .ZN(_14274_)
  );
  INV_X1 _49200_ (
    .A(_14274_),
    .ZN(_14275_)
  );
  AND2_X1 _49201_ (
    .A1(\cpuregs[3] [9]),
    .A2(_12681_),
    .ZN(_14276_)
  );
  INV_X1 _49202_ (
    .A(_14276_),
    .ZN(_14277_)
  );
  AND2_X1 _49203_ (
    .A1(_14275_),
    .A2(_14277_),
    .ZN(_14278_)
  );
  INV_X1 _49204_ (
    .A(_14278_),
    .ZN(_00753_)
  );
  AND2_X1 _49205_ (
    .A1(_12680_),
    .A2(_13018_),
    .ZN(_14279_)
  );
  INV_X1 _49206_ (
    .A(_14279_),
    .ZN(_14280_)
  );
  AND2_X1 _49207_ (
    .A1(\cpuregs[3] [10]),
    .A2(_12681_),
    .ZN(_14281_)
  );
  INV_X1 _49208_ (
    .A(_14281_),
    .ZN(_14282_)
  );
  AND2_X1 _49209_ (
    .A1(_14280_),
    .A2(_14282_),
    .ZN(_14283_)
  );
  INV_X1 _49210_ (
    .A(_14283_),
    .ZN(_00754_)
  );
  AND2_X1 _49211_ (
    .A1(_12680_),
    .A2(_13033_),
    .ZN(_14284_)
  );
  INV_X1 _49212_ (
    .A(_14284_),
    .ZN(_14285_)
  );
  AND2_X1 _49213_ (
    .A1(\cpuregs[3] [11]),
    .A2(_12681_),
    .ZN(_14286_)
  );
  INV_X1 _49214_ (
    .A(_14286_),
    .ZN(_14287_)
  );
  AND2_X1 _49215_ (
    .A1(_14285_),
    .A2(_14287_),
    .ZN(_14288_)
  );
  INV_X1 _49216_ (
    .A(_14288_),
    .ZN(_00755_)
  );
  AND2_X1 _49217_ (
    .A1(_12680_),
    .A2(_13048_),
    .ZN(_14289_)
  );
  INV_X1 _49218_ (
    .A(_14289_),
    .ZN(_14290_)
  );
  AND2_X1 _49219_ (
    .A1(\cpuregs[3] [12]),
    .A2(_12681_),
    .ZN(_14291_)
  );
  INV_X1 _49220_ (
    .A(_14291_),
    .ZN(_14292_)
  );
  AND2_X1 _49221_ (
    .A1(_14290_),
    .A2(_14292_),
    .ZN(_14293_)
  );
  INV_X1 _49222_ (
    .A(_14293_),
    .ZN(_00756_)
  );
  AND2_X1 _49223_ (
    .A1(_12680_),
    .A2(_13063_),
    .ZN(_14294_)
  );
  INV_X1 _49224_ (
    .A(_14294_),
    .ZN(_14295_)
  );
  AND2_X1 _49225_ (
    .A1(\cpuregs[3] [13]),
    .A2(_12681_),
    .ZN(_14296_)
  );
  INV_X1 _49226_ (
    .A(_14296_),
    .ZN(_14297_)
  );
  AND2_X1 _49227_ (
    .A1(_14295_),
    .A2(_14297_),
    .ZN(_14298_)
  );
  INV_X1 _49228_ (
    .A(_14298_),
    .ZN(_00757_)
  );
  AND2_X1 _49229_ (
    .A1(\cpuregs[3] [14]),
    .A2(_12681_),
    .ZN(_14299_)
  );
  INV_X1 _49230_ (
    .A(_14299_),
    .ZN(_14300_)
  );
  AND2_X1 _49231_ (
    .A1(_12680_),
    .A2(_13078_),
    .ZN(_14301_)
  );
  INV_X1 _49232_ (
    .A(_14301_),
    .ZN(_14302_)
  );
  AND2_X1 _49233_ (
    .A1(_14300_),
    .A2(_14302_),
    .ZN(_14303_)
  );
  INV_X1 _49234_ (
    .A(_14303_),
    .ZN(_00758_)
  );
  AND2_X1 _49235_ (
    .A1(_12680_),
    .A2(_13093_),
    .ZN(_14304_)
  );
  INV_X1 _49236_ (
    .A(_14304_),
    .ZN(_14305_)
  );
  AND2_X1 _49237_ (
    .A1(\cpuregs[3] [15]),
    .A2(_12681_),
    .ZN(_14306_)
  );
  INV_X1 _49238_ (
    .A(_14306_),
    .ZN(_14307_)
  );
  AND2_X1 _49239_ (
    .A1(_14305_),
    .A2(_14307_),
    .ZN(_14308_)
  );
  INV_X1 _49240_ (
    .A(_14308_),
    .ZN(_00759_)
  );
  AND2_X1 _49241_ (
    .A1(_12680_),
    .A2(_13108_),
    .ZN(_14309_)
  );
  INV_X1 _49242_ (
    .A(_14309_),
    .ZN(_14310_)
  );
  AND2_X1 _49243_ (
    .A1(\cpuregs[3] [16]),
    .A2(_12681_),
    .ZN(_14311_)
  );
  INV_X1 _49244_ (
    .A(_14311_),
    .ZN(_14312_)
  );
  AND2_X1 _49245_ (
    .A1(_14310_),
    .A2(_14312_),
    .ZN(_14313_)
  );
  INV_X1 _49246_ (
    .A(_14313_),
    .ZN(_00760_)
  );
  AND2_X1 _49247_ (
    .A1(_12680_),
    .A2(_13123_),
    .ZN(_14314_)
  );
  INV_X1 _49248_ (
    .A(_14314_),
    .ZN(_14315_)
  );
  AND2_X1 _49249_ (
    .A1(\cpuregs[3] [17]),
    .A2(_12681_),
    .ZN(_14316_)
  );
  INV_X1 _49250_ (
    .A(_14316_),
    .ZN(_14317_)
  );
  AND2_X1 _49251_ (
    .A1(_14315_),
    .A2(_14317_),
    .ZN(_14318_)
  );
  INV_X1 _49252_ (
    .A(_14318_),
    .ZN(_00761_)
  );
  AND2_X1 _49253_ (
    .A1(_12680_),
    .A2(_13139_),
    .ZN(_14319_)
  );
  INV_X1 _49254_ (
    .A(_14319_),
    .ZN(_14320_)
  );
  AND2_X1 _49255_ (
    .A1(\cpuregs[3] [18]),
    .A2(_12681_),
    .ZN(_14321_)
  );
  INV_X1 _49256_ (
    .A(_14321_),
    .ZN(_14322_)
  );
  AND2_X1 _49257_ (
    .A1(_14320_),
    .A2(_14322_),
    .ZN(_14323_)
  );
  INV_X1 _49258_ (
    .A(_14323_),
    .ZN(_00762_)
  );
  AND2_X1 _49259_ (
    .A1(_12680_),
    .A2(_13154_),
    .ZN(_14324_)
  );
  INV_X1 _49260_ (
    .A(_14324_),
    .ZN(_14325_)
  );
  AND2_X1 _49261_ (
    .A1(\cpuregs[3] [19]),
    .A2(_12681_),
    .ZN(_14326_)
  );
  INV_X1 _49262_ (
    .A(_14326_),
    .ZN(_14327_)
  );
  AND2_X1 _49263_ (
    .A1(_14325_),
    .A2(_14327_),
    .ZN(_14328_)
  );
  INV_X1 _49264_ (
    .A(_14328_),
    .ZN(_00763_)
  );
  AND2_X1 _49265_ (
    .A1(_12680_),
    .A2(_13169_),
    .ZN(_14329_)
  );
  INV_X1 _49266_ (
    .A(_14329_),
    .ZN(_14330_)
  );
  AND2_X1 _49267_ (
    .A1(\cpuregs[3] [20]),
    .A2(_12681_),
    .ZN(_14331_)
  );
  INV_X1 _49268_ (
    .A(_14331_),
    .ZN(_14332_)
  );
  AND2_X1 _49269_ (
    .A1(_14330_),
    .A2(_14332_),
    .ZN(_14333_)
  );
  INV_X1 _49270_ (
    .A(_14333_),
    .ZN(_00764_)
  );
  AND2_X1 _49271_ (
    .A1(_12680_),
    .A2(_13184_),
    .ZN(_14334_)
  );
  INV_X1 _49272_ (
    .A(_14334_),
    .ZN(_14335_)
  );
  AND2_X1 _49273_ (
    .A1(\cpuregs[3] [21]),
    .A2(_12681_),
    .ZN(_14336_)
  );
  INV_X1 _49274_ (
    .A(_14336_),
    .ZN(_14337_)
  );
  AND2_X1 _49275_ (
    .A1(_14335_),
    .A2(_14337_),
    .ZN(_14338_)
  );
  INV_X1 _49276_ (
    .A(_14338_),
    .ZN(_00765_)
  );
  AND2_X1 _49277_ (
    .A1(_12680_),
    .A2(_13199_),
    .ZN(_14339_)
  );
  INV_X1 _49278_ (
    .A(_14339_),
    .ZN(_14340_)
  );
  AND2_X1 _49279_ (
    .A1(\cpuregs[3] [22]),
    .A2(_12681_),
    .ZN(_14341_)
  );
  INV_X1 _49280_ (
    .A(_14341_),
    .ZN(_14342_)
  );
  AND2_X1 _49281_ (
    .A1(_14340_),
    .A2(_14342_),
    .ZN(_14343_)
  );
  INV_X1 _49282_ (
    .A(_14343_),
    .ZN(_00766_)
  );
  AND2_X1 _49283_ (
    .A1(_12680_),
    .A2(_13214_),
    .ZN(_14344_)
  );
  INV_X1 _49284_ (
    .A(_14344_),
    .ZN(_14345_)
  );
  AND2_X1 _49285_ (
    .A1(\cpuregs[3] [23]),
    .A2(_12681_),
    .ZN(_14346_)
  );
  INV_X1 _49286_ (
    .A(_14346_),
    .ZN(_14347_)
  );
  AND2_X1 _49287_ (
    .A1(_14345_),
    .A2(_14347_),
    .ZN(_14348_)
  );
  INV_X1 _49288_ (
    .A(_14348_),
    .ZN(_00767_)
  );
  AND2_X1 _49289_ (
    .A1(_12680_),
    .A2(_13229_),
    .ZN(_14349_)
  );
  INV_X1 _49290_ (
    .A(_14349_),
    .ZN(_14350_)
  );
  AND2_X1 _49291_ (
    .A1(\cpuregs[3] [24]),
    .A2(_12681_),
    .ZN(_14351_)
  );
  INV_X1 _49292_ (
    .A(_14351_),
    .ZN(_14352_)
  );
  AND2_X1 _49293_ (
    .A1(_14350_),
    .A2(_14352_),
    .ZN(_14353_)
  );
  INV_X1 _49294_ (
    .A(_14353_),
    .ZN(_00768_)
  );
  AND2_X1 _49295_ (
    .A1(_12680_),
    .A2(_13244_),
    .ZN(_14354_)
  );
  INV_X1 _49296_ (
    .A(_14354_),
    .ZN(_14355_)
  );
  AND2_X1 _49297_ (
    .A1(\cpuregs[3] [25]),
    .A2(_12681_),
    .ZN(_14356_)
  );
  INV_X1 _49298_ (
    .A(_14356_),
    .ZN(_14357_)
  );
  AND2_X1 _49299_ (
    .A1(_14355_),
    .A2(_14357_),
    .ZN(_14358_)
  );
  INV_X1 _49300_ (
    .A(_14358_),
    .ZN(_00769_)
  );
  AND2_X1 _49301_ (
    .A1(_12680_),
    .A2(_13259_),
    .ZN(_14359_)
  );
  INV_X1 _49302_ (
    .A(_14359_),
    .ZN(_14360_)
  );
  AND2_X1 _49303_ (
    .A1(\cpuregs[3] [26]),
    .A2(_12681_),
    .ZN(_14361_)
  );
  INV_X1 _49304_ (
    .A(_14361_),
    .ZN(_14362_)
  );
  AND2_X1 _49305_ (
    .A1(_14360_),
    .A2(_14362_),
    .ZN(_14363_)
  );
  INV_X1 _49306_ (
    .A(_14363_),
    .ZN(_00770_)
  );
  AND2_X1 _49307_ (
    .A1(_12680_),
    .A2(_13274_),
    .ZN(_14364_)
  );
  INV_X1 _49308_ (
    .A(_14364_),
    .ZN(_14365_)
  );
  AND2_X1 _49309_ (
    .A1(\cpuregs[3] [27]),
    .A2(_12681_),
    .ZN(_14366_)
  );
  INV_X1 _49310_ (
    .A(_14366_),
    .ZN(_14367_)
  );
  AND2_X1 _49311_ (
    .A1(_14365_),
    .A2(_14367_),
    .ZN(_14368_)
  );
  INV_X1 _49312_ (
    .A(_14368_),
    .ZN(_00771_)
  );
  AND2_X1 _49313_ (
    .A1(_12680_),
    .A2(_13289_),
    .ZN(_14369_)
  );
  INV_X1 _49314_ (
    .A(_14369_),
    .ZN(_14370_)
  );
  AND2_X1 _49315_ (
    .A1(\cpuregs[3] [28]),
    .A2(_12681_),
    .ZN(_14371_)
  );
  INV_X1 _49316_ (
    .A(_14371_),
    .ZN(_14372_)
  );
  AND2_X1 _49317_ (
    .A1(_14370_),
    .A2(_14372_),
    .ZN(_14373_)
  );
  INV_X1 _49318_ (
    .A(_14373_),
    .ZN(_00772_)
  );
  AND2_X1 _49319_ (
    .A1(_12680_),
    .A2(_13304_),
    .ZN(_14374_)
  );
  INV_X1 _49320_ (
    .A(_14374_),
    .ZN(_14375_)
  );
  AND2_X1 _49321_ (
    .A1(\cpuregs[3] [29]),
    .A2(_12681_),
    .ZN(_14376_)
  );
  INV_X1 _49322_ (
    .A(_14376_),
    .ZN(_14377_)
  );
  AND2_X1 _49323_ (
    .A1(_14375_),
    .A2(_14377_),
    .ZN(_14378_)
  );
  INV_X1 _49324_ (
    .A(_14378_),
    .ZN(_00773_)
  );
  AND2_X1 _49325_ (
    .A1(_12680_),
    .A2(_13319_),
    .ZN(_14379_)
  );
  INV_X1 _49326_ (
    .A(_14379_),
    .ZN(_14380_)
  );
  AND2_X1 _49327_ (
    .A1(\cpuregs[3] [30]),
    .A2(_12681_),
    .ZN(_14381_)
  );
  INV_X1 _49328_ (
    .A(_14381_),
    .ZN(_14382_)
  );
  AND2_X1 _49329_ (
    .A1(_14380_),
    .A2(_14382_),
    .ZN(_14383_)
  );
  INV_X1 _49330_ (
    .A(_14383_),
    .ZN(_00774_)
  );
  AND2_X1 _49331_ (
    .A1(_12783_),
    .A2(_12874_),
    .ZN(_14384_)
  );
  INV_X1 _49332_ (
    .A(_14384_),
    .ZN(_14385_)
  );
  AND2_X1 _49333_ (
    .A1(\cpuregs[1] [0]),
    .A2(_12784_),
    .ZN(_14386_)
  );
  INV_X1 _49334_ (
    .A(_14386_),
    .ZN(_14387_)
  );
  AND2_X1 _49335_ (
    .A1(_14385_),
    .A2(_14387_),
    .ZN(_14388_)
  );
  INV_X1 _49336_ (
    .A(_14388_),
    .ZN(_00775_)
  );
  AND2_X1 _49337_ (
    .A1(_12783_),
    .A2(_12886_),
    .ZN(_14389_)
  );
  INV_X1 _49338_ (
    .A(_14389_),
    .ZN(_14390_)
  );
  AND2_X1 _49339_ (
    .A1(\cpuregs[1] [1]),
    .A2(_12784_),
    .ZN(_14391_)
  );
  INV_X1 _49340_ (
    .A(_14391_),
    .ZN(_14392_)
  );
  AND2_X1 _49341_ (
    .A1(_14390_),
    .A2(_14392_),
    .ZN(_14393_)
  );
  INV_X1 _49342_ (
    .A(_14393_),
    .ZN(_00776_)
  );
  AND2_X1 _49343_ (
    .A1(_12783_),
    .A2(_12900_),
    .ZN(_14394_)
  );
  INV_X1 _49344_ (
    .A(_14394_),
    .ZN(_14395_)
  );
  AND2_X1 _49345_ (
    .A1(\cpuregs[1] [2]),
    .A2(_12784_),
    .ZN(_14396_)
  );
  INV_X1 _49346_ (
    .A(_14396_),
    .ZN(_14397_)
  );
  AND2_X1 _49347_ (
    .A1(_14395_),
    .A2(_14397_),
    .ZN(_14398_)
  );
  INV_X1 _49348_ (
    .A(_14398_),
    .ZN(_00777_)
  );
  AND2_X1 _49349_ (
    .A1(_12783_),
    .A2(_12913_),
    .ZN(_14399_)
  );
  INV_X1 _49350_ (
    .A(_14399_),
    .ZN(_14400_)
  );
  AND2_X1 _49351_ (
    .A1(\cpuregs[1] [3]),
    .A2(_12784_),
    .ZN(_14401_)
  );
  INV_X1 _49352_ (
    .A(_14401_),
    .ZN(_14402_)
  );
  AND2_X1 _49353_ (
    .A1(_14400_),
    .A2(_14402_),
    .ZN(_14403_)
  );
  INV_X1 _49354_ (
    .A(_14403_),
    .ZN(_00778_)
  );
  AND2_X1 _49355_ (
    .A1(\cpuregs[1] [4]),
    .A2(_12784_),
    .ZN(_14404_)
  );
  INV_X1 _49356_ (
    .A(_14404_),
    .ZN(_14405_)
  );
  AND2_X1 _49357_ (
    .A1(_12783_),
    .A2(_12928_),
    .ZN(_14406_)
  );
  INV_X1 _49358_ (
    .A(_14406_),
    .ZN(_14407_)
  );
  AND2_X1 _49359_ (
    .A1(_14405_),
    .A2(_14407_),
    .ZN(_14408_)
  );
  INV_X1 _49360_ (
    .A(_14408_),
    .ZN(_00779_)
  );
  AND2_X1 _49361_ (
    .A1(_12783_),
    .A2(_12943_),
    .ZN(_14409_)
  );
  INV_X1 _49362_ (
    .A(_14409_),
    .ZN(_14410_)
  );
  AND2_X1 _49363_ (
    .A1(\cpuregs[1] [5]),
    .A2(_12784_),
    .ZN(_14411_)
  );
  INV_X1 _49364_ (
    .A(_14411_),
    .ZN(_14412_)
  );
  AND2_X1 _49365_ (
    .A1(_14410_),
    .A2(_14412_),
    .ZN(_14413_)
  );
  INV_X1 _49366_ (
    .A(_14413_),
    .ZN(_00780_)
  );
  AND2_X1 _49367_ (
    .A1(_12783_),
    .A2(_12958_),
    .ZN(_14414_)
  );
  INV_X1 _49368_ (
    .A(_14414_),
    .ZN(_14415_)
  );
  AND2_X1 _49369_ (
    .A1(\cpuregs[1] [6]),
    .A2(_12784_),
    .ZN(_14416_)
  );
  INV_X1 _49370_ (
    .A(_14416_),
    .ZN(_14417_)
  );
  AND2_X1 _49371_ (
    .A1(_14415_),
    .A2(_14417_),
    .ZN(_14418_)
  );
  INV_X1 _49372_ (
    .A(_14418_),
    .ZN(_00781_)
  );
  AND2_X1 _49373_ (
    .A1(_12783_),
    .A2(_12973_),
    .ZN(_14419_)
  );
  INV_X1 _49374_ (
    .A(_14419_),
    .ZN(_14420_)
  );
  AND2_X1 _49375_ (
    .A1(\cpuregs[1] [7]),
    .A2(_12784_),
    .ZN(_14421_)
  );
  INV_X1 _49376_ (
    .A(_14421_),
    .ZN(_14422_)
  );
  AND2_X1 _49377_ (
    .A1(_14420_),
    .A2(_14422_),
    .ZN(_14423_)
  );
  INV_X1 _49378_ (
    .A(_14423_),
    .ZN(_00782_)
  );
  AND2_X1 _49379_ (
    .A1(_12783_),
    .A2(_12988_),
    .ZN(_14424_)
  );
  INV_X1 _49380_ (
    .A(_14424_),
    .ZN(_14425_)
  );
  AND2_X1 _49381_ (
    .A1(\cpuregs[1] [8]),
    .A2(_12784_),
    .ZN(_14426_)
  );
  INV_X1 _49382_ (
    .A(_14426_),
    .ZN(_14427_)
  );
  AND2_X1 _49383_ (
    .A1(_14425_),
    .A2(_14427_),
    .ZN(_14428_)
  );
  INV_X1 _49384_ (
    .A(_14428_),
    .ZN(_00783_)
  );
  AND2_X1 _49385_ (
    .A1(_12783_),
    .A2(_13003_),
    .ZN(_14429_)
  );
  INV_X1 _49386_ (
    .A(_14429_),
    .ZN(_14430_)
  );
  AND2_X1 _49387_ (
    .A1(\cpuregs[1] [9]),
    .A2(_12784_),
    .ZN(_14431_)
  );
  INV_X1 _49388_ (
    .A(_14431_),
    .ZN(_14432_)
  );
  AND2_X1 _49389_ (
    .A1(_14430_),
    .A2(_14432_),
    .ZN(_14433_)
  );
  INV_X1 _49390_ (
    .A(_14433_),
    .ZN(_00784_)
  );
  AND2_X1 _49391_ (
    .A1(_12783_),
    .A2(_13018_),
    .ZN(_14434_)
  );
  INV_X1 _49392_ (
    .A(_14434_),
    .ZN(_14435_)
  );
  AND2_X1 _49393_ (
    .A1(\cpuregs[1] [10]),
    .A2(_12784_),
    .ZN(_14436_)
  );
  INV_X1 _49394_ (
    .A(_14436_),
    .ZN(_14437_)
  );
  AND2_X1 _49395_ (
    .A1(_14435_),
    .A2(_14437_),
    .ZN(_14438_)
  );
  INV_X1 _49396_ (
    .A(_14438_),
    .ZN(_00785_)
  );
  AND2_X1 _49397_ (
    .A1(_12783_),
    .A2(_13033_),
    .ZN(_14439_)
  );
  INV_X1 _49398_ (
    .A(_14439_),
    .ZN(_14440_)
  );
  AND2_X1 _49399_ (
    .A1(\cpuregs[1] [11]),
    .A2(_12784_),
    .ZN(_14441_)
  );
  INV_X1 _49400_ (
    .A(_14441_),
    .ZN(_14442_)
  );
  AND2_X1 _49401_ (
    .A1(_14440_),
    .A2(_14442_),
    .ZN(_14443_)
  );
  INV_X1 _49402_ (
    .A(_14443_),
    .ZN(_00786_)
  );
  AND2_X1 _49403_ (
    .A1(_12783_),
    .A2(_13048_),
    .ZN(_14444_)
  );
  INV_X1 _49404_ (
    .A(_14444_),
    .ZN(_14445_)
  );
  AND2_X1 _49405_ (
    .A1(\cpuregs[1] [12]),
    .A2(_12784_),
    .ZN(_14446_)
  );
  INV_X1 _49406_ (
    .A(_14446_),
    .ZN(_14447_)
  );
  AND2_X1 _49407_ (
    .A1(_14445_),
    .A2(_14447_),
    .ZN(_14448_)
  );
  INV_X1 _49408_ (
    .A(_14448_),
    .ZN(_00787_)
  );
  AND2_X1 _49409_ (
    .A1(_12783_),
    .A2(_13063_),
    .ZN(_14449_)
  );
  INV_X1 _49410_ (
    .A(_14449_),
    .ZN(_14450_)
  );
  AND2_X1 _49411_ (
    .A1(\cpuregs[1] [13]),
    .A2(_12784_),
    .ZN(_14451_)
  );
  INV_X1 _49412_ (
    .A(_14451_),
    .ZN(_14452_)
  );
  AND2_X1 _49413_ (
    .A1(_14450_),
    .A2(_14452_),
    .ZN(_14453_)
  );
  INV_X1 _49414_ (
    .A(_14453_),
    .ZN(_00788_)
  );
  AND2_X1 _49415_ (
    .A1(_12783_),
    .A2(_13078_),
    .ZN(_14454_)
  );
  INV_X1 _49416_ (
    .A(_14454_),
    .ZN(_14455_)
  );
  AND2_X1 _49417_ (
    .A1(\cpuregs[1] [14]),
    .A2(_12784_),
    .ZN(_14456_)
  );
  INV_X1 _49418_ (
    .A(_14456_),
    .ZN(_14457_)
  );
  AND2_X1 _49419_ (
    .A1(_14455_),
    .A2(_14457_),
    .ZN(_14458_)
  );
  INV_X1 _49420_ (
    .A(_14458_),
    .ZN(_00789_)
  );
  AND2_X1 _49421_ (
    .A1(_12783_),
    .A2(_13093_),
    .ZN(_14459_)
  );
  INV_X1 _49422_ (
    .A(_14459_),
    .ZN(_14460_)
  );
  AND2_X1 _49423_ (
    .A1(\cpuregs[1] [15]),
    .A2(_12784_),
    .ZN(_14461_)
  );
  INV_X1 _49424_ (
    .A(_14461_),
    .ZN(_14462_)
  );
  AND2_X1 _49425_ (
    .A1(_14460_),
    .A2(_14462_),
    .ZN(_14463_)
  );
  INV_X1 _49426_ (
    .A(_14463_),
    .ZN(_00790_)
  );
  AND2_X1 _49427_ (
    .A1(\cpuregs[1] [16]),
    .A2(_12784_),
    .ZN(_14464_)
  );
  INV_X1 _49428_ (
    .A(_14464_),
    .ZN(_14465_)
  );
  AND2_X1 _49429_ (
    .A1(_12783_),
    .A2(_13108_),
    .ZN(_14466_)
  );
  INV_X1 _49430_ (
    .A(_14466_),
    .ZN(_14467_)
  );
  AND2_X1 _49431_ (
    .A1(_14465_),
    .A2(_14467_),
    .ZN(_14468_)
  );
  INV_X1 _49432_ (
    .A(_14468_),
    .ZN(_00791_)
  );
  AND2_X1 _49433_ (
    .A1(_12783_),
    .A2(_13123_),
    .ZN(_14469_)
  );
  INV_X1 _49434_ (
    .A(_14469_),
    .ZN(_14470_)
  );
  AND2_X1 _49435_ (
    .A1(\cpuregs[1] [17]),
    .A2(_12784_),
    .ZN(_14471_)
  );
  INV_X1 _49436_ (
    .A(_14471_),
    .ZN(_14472_)
  );
  AND2_X1 _49437_ (
    .A1(_14470_),
    .A2(_14472_),
    .ZN(_14473_)
  );
  INV_X1 _49438_ (
    .A(_14473_),
    .ZN(_00792_)
  );
  AND2_X1 _49439_ (
    .A1(_12783_),
    .A2(_13139_),
    .ZN(_14474_)
  );
  INV_X1 _49440_ (
    .A(_14474_),
    .ZN(_14475_)
  );
  AND2_X1 _49441_ (
    .A1(\cpuregs[1] [18]),
    .A2(_12784_),
    .ZN(_14476_)
  );
  INV_X1 _49442_ (
    .A(_14476_),
    .ZN(_14477_)
  );
  AND2_X1 _49443_ (
    .A1(_14475_),
    .A2(_14477_),
    .ZN(_14478_)
  );
  INV_X1 _49444_ (
    .A(_14478_),
    .ZN(_00793_)
  );
  AND2_X1 _49445_ (
    .A1(_12783_),
    .A2(_13154_),
    .ZN(_14479_)
  );
  INV_X1 _49446_ (
    .A(_14479_),
    .ZN(_14480_)
  );
  AND2_X1 _49447_ (
    .A1(\cpuregs[1] [19]),
    .A2(_12784_),
    .ZN(_14481_)
  );
  INV_X1 _49448_ (
    .A(_14481_),
    .ZN(_14482_)
  );
  AND2_X1 _49449_ (
    .A1(_14480_),
    .A2(_14482_),
    .ZN(_14483_)
  );
  INV_X1 _49450_ (
    .A(_14483_),
    .ZN(_00794_)
  );
  AND2_X1 _49451_ (
    .A1(_12783_),
    .A2(_13169_),
    .ZN(_14484_)
  );
  INV_X1 _49452_ (
    .A(_14484_),
    .ZN(_14485_)
  );
  AND2_X1 _49453_ (
    .A1(\cpuregs[1] [20]),
    .A2(_12784_),
    .ZN(_14486_)
  );
  INV_X1 _49454_ (
    .A(_14486_),
    .ZN(_14487_)
  );
  AND2_X1 _49455_ (
    .A1(_14485_),
    .A2(_14487_),
    .ZN(_14488_)
  );
  INV_X1 _49456_ (
    .A(_14488_),
    .ZN(_00795_)
  );
  AND2_X1 _49457_ (
    .A1(_12783_),
    .A2(_13184_),
    .ZN(_14489_)
  );
  INV_X1 _49458_ (
    .A(_14489_),
    .ZN(_14490_)
  );
  AND2_X1 _49459_ (
    .A1(\cpuregs[1] [21]),
    .A2(_12784_),
    .ZN(_14491_)
  );
  INV_X1 _49460_ (
    .A(_14491_),
    .ZN(_14492_)
  );
  AND2_X1 _49461_ (
    .A1(_14490_),
    .A2(_14492_),
    .ZN(_14493_)
  );
  INV_X1 _49462_ (
    .A(_14493_),
    .ZN(_00796_)
  );
  AND2_X1 _49463_ (
    .A1(_12783_),
    .A2(_13199_),
    .ZN(_14494_)
  );
  INV_X1 _49464_ (
    .A(_14494_),
    .ZN(_14495_)
  );
  AND2_X1 _49465_ (
    .A1(\cpuregs[1] [22]),
    .A2(_12784_),
    .ZN(_14496_)
  );
  INV_X1 _49466_ (
    .A(_14496_),
    .ZN(_14497_)
  );
  AND2_X1 _49467_ (
    .A1(_14495_),
    .A2(_14497_),
    .ZN(_14498_)
  );
  INV_X1 _49468_ (
    .A(_14498_),
    .ZN(_00797_)
  );
  AND2_X1 _49469_ (
    .A1(_12783_),
    .A2(_13214_),
    .ZN(_14499_)
  );
  INV_X1 _49470_ (
    .A(_14499_),
    .ZN(_14500_)
  );
  AND2_X1 _49471_ (
    .A1(\cpuregs[1] [23]),
    .A2(_12784_),
    .ZN(_14501_)
  );
  INV_X1 _49472_ (
    .A(_14501_),
    .ZN(_14502_)
  );
  AND2_X1 _49473_ (
    .A1(_14500_),
    .A2(_14502_),
    .ZN(_14503_)
  );
  INV_X1 _49474_ (
    .A(_14503_),
    .ZN(_00798_)
  );
  AND2_X1 _49475_ (
    .A1(_12783_),
    .A2(_13229_),
    .ZN(_14504_)
  );
  INV_X1 _49476_ (
    .A(_14504_),
    .ZN(_14505_)
  );
  AND2_X1 _49477_ (
    .A1(\cpuregs[1] [24]),
    .A2(_12784_),
    .ZN(_14506_)
  );
  INV_X1 _49478_ (
    .A(_14506_),
    .ZN(_14507_)
  );
  AND2_X1 _49479_ (
    .A1(_14505_),
    .A2(_14507_),
    .ZN(_14508_)
  );
  INV_X1 _49480_ (
    .A(_14508_),
    .ZN(_00799_)
  );
  AND2_X1 _49481_ (
    .A1(_12783_),
    .A2(_13244_),
    .ZN(_14509_)
  );
  INV_X1 _49482_ (
    .A(_14509_),
    .ZN(_14510_)
  );
  AND2_X1 _49483_ (
    .A1(\cpuregs[1] [25]),
    .A2(_12784_),
    .ZN(_14511_)
  );
  INV_X1 _49484_ (
    .A(_14511_),
    .ZN(_14512_)
  );
  AND2_X1 _49485_ (
    .A1(_14510_),
    .A2(_14512_),
    .ZN(_14513_)
  );
  INV_X1 _49486_ (
    .A(_14513_),
    .ZN(_00800_)
  );
  AND2_X1 _49487_ (
    .A1(_12783_),
    .A2(_13259_),
    .ZN(_14514_)
  );
  INV_X1 _49488_ (
    .A(_14514_),
    .ZN(_14515_)
  );
  AND2_X1 _49489_ (
    .A1(\cpuregs[1] [26]),
    .A2(_12784_),
    .ZN(_14516_)
  );
  INV_X1 _49490_ (
    .A(_14516_),
    .ZN(_14517_)
  );
  AND2_X1 _49491_ (
    .A1(_14515_),
    .A2(_14517_),
    .ZN(_14518_)
  );
  INV_X1 _49492_ (
    .A(_14518_),
    .ZN(_00801_)
  );
  AND2_X1 _49493_ (
    .A1(_12783_),
    .A2(_13274_),
    .ZN(_14519_)
  );
  INV_X1 _49494_ (
    .A(_14519_),
    .ZN(_14520_)
  );
  AND2_X1 _49495_ (
    .A1(\cpuregs[1] [27]),
    .A2(_12784_),
    .ZN(_14521_)
  );
  INV_X1 _49496_ (
    .A(_14521_),
    .ZN(_14522_)
  );
  AND2_X1 _49497_ (
    .A1(_14520_),
    .A2(_14522_),
    .ZN(_14523_)
  );
  INV_X1 _49498_ (
    .A(_14523_),
    .ZN(_00802_)
  );
  AND2_X1 _49499_ (
    .A1(_12783_),
    .A2(_13289_),
    .ZN(_14524_)
  );
  INV_X1 _49500_ (
    .A(_14524_),
    .ZN(_14525_)
  );
  AND2_X1 _49501_ (
    .A1(\cpuregs[1] [28]),
    .A2(_12784_),
    .ZN(_14526_)
  );
  INV_X1 _49502_ (
    .A(_14526_),
    .ZN(_14527_)
  );
  AND2_X1 _49503_ (
    .A1(_14525_),
    .A2(_14527_),
    .ZN(_14528_)
  );
  INV_X1 _49504_ (
    .A(_14528_),
    .ZN(_00803_)
  );
  AND2_X1 _49505_ (
    .A1(_12783_),
    .A2(_13304_),
    .ZN(_14529_)
  );
  INV_X1 _49506_ (
    .A(_14529_),
    .ZN(_14530_)
  );
  AND2_X1 _49507_ (
    .A1(\cpuregs[1] [29]),
    .A2(_12784_),
    .ZN(_14531_)
  );
  INV_X1 _49508_ (
    .A(_14531_),
    .ZN(_14532_)
  );
  AND2_X1 _49509_ (
    .A1(_14530_),
    .A2(_14532_),
    .ZN(_14533_)
  );
  INV_X1 _49510_ (
    .A(_14533_),
    .ZN(_00804_)
  );
  AND2_X1 _49511_ (
    .A1(_12783_),
    .A2(_13319_),
    .ZN(_14534_)
  );
  INV_X1 _49512_ (
    .A(_14534_),
    .ZN(_14535_)
  );
  AND2_X1 _49513_ (
    .A1(\cpuregs[1] [30]),
    .A2(_12784_),
    .ZN(_14536_)
  );
  INV_X1 _49514_ (
    .A(_14536_),
    .ZN(_14537_)
  );
  AND2_X1 _49515_ (
    .A1(_14535_),
    .A2(_14537_),
    .ZN(_14538_)
  );
  INV_X1 _49516_ (
    .A(_14538_),
    .ZN(_00805_)
  );
  AND2_X1 _49517_ (
    .A1(_12704_),
    .A2(_12872_),
    .ZN(_14539_)
  );
  INV_X1 _49518_ (
    .A(_14539_),
    .ZN(_14540_)
  );
  AND2_X1 _49519_ (
    .A1(_21537_),
    .A2(_12705_),
    .ZN(_14541_)
  );
  INV_X1 _49520_ (
    .A(_14541_),
    .ZN(_14542_)
  );
  AND2_X1 _49521_ (
    .A1(_14540_),
    .A2(_14542_),
    .ZN(_00806_)
  );
  AND2_X1 _49522_ (
    .A1(_12704_),
    .A2(_12884_),
    .ZN(_14543_)
  );
  INV_X1 _49523_ (
    .A(_14543_),
    .ZN(_14544_)
  );
  AND2_X1 _49524_ (
    .A1(_21538_),
    .A2(_12705_),
    .ZN(_14545_)
  );
  INV_X1 _49525_ (
    .A(_14545_),
    .ZN(_14546_)
  );
  AND2_X1 _49526_ (
    .A1(_14544_),
    .A2(_14546_),
    .ZN(_00807_)
  );
  AND2_X1 _49527_ (
    .A1(_12704_),
    .A2(_12898_),
    .ZN(_14547_)
  );
  INV_X1 _49528_ (
    .A(_14547_),
    .ZN(_14548_)
  );
  AND2_X1 _49529_ (
    .A1(_21539_),
    .A2(_12705_),
    .ZN(_14549_)
  );
  INV_X1 _49530_ (
    .A(_14549_),
    .ZN(_14550_)
  );
  AND2_X1 _49531_ (
    .A1(_14548_),
    .A2(_14550_),
    .ZN(_00808_)
  );
  AND2_X1 _49532_ (
    .A1(_12704_),
    .A2(_12911_),
    .ZN(_14551_)
  );
  INV_X1 _49533_ (
    .A(_14551_),
    .ZN(_14552_)
  );
  AND2_X1 _49534_ (
    .A1(_21540_),
    .A2(_12705_),
    .ZN(_14553_)
  );
  INV_X1 _49535_ (
    .A(_14553_),
    .ZN(_14554_)
  );
  AND2_X1 _49536_ (
    .A1(_14552_),
    .A2(_14554_),
    .ZN(_00809_)
  );
  AND2_X1 _49537_ (
    .A1(_12704_),
    .A2(_12928_),
    .ZN(_14555_)
  );
  INV_X1 _49538_ (
    .A(_14555_),
    .ZN(_14556_)
  );
  AND2_X1 _49539_ (
    .A1(\cpuregs[2] [4]),
    .A2(_12705_),
    .ZN(_14557_)
  );
  INV_X1 _49540_ (
    .A(_14557_),
    .ZN(_14558_)
  );
  AND2_X1 _49541_ (
    .A1(_14556_),
    .A2(_14558_),
    .ZN(_14559_)
  );
  INV_X1 _49542_ (
    .A(_14559_),
    .ZN(_00810_)
  );
  AND2_X1 _49543_ (
    .A1(_12704_),
    .A2(_12941_),
    .ZN(_14560_)
  );
  INV_X1 _49544_ (
    .A(_14560_),
    .ZN(_14561_)
  );
  AND2_X1 _49545_ (
    .A1(_21542_),
    .A2(_12705_),
    .ZN(_14562_)
  );
  INV_X1 _49546_ (
    .A(_14562_),
    .ZN(_14563_)
  );
  AND2_X1 _49547_ (
    .A1(_14561_),
    .A2(_14563_),
    .ZN(_00811_)
  );
  AND2_X1 _49548_ (
    .A1(_12704_),
    .A2(_12958_),
    .ZN(_14564_)
  );
  INV_X1 _49549_ (
    .A(_14564_),
    .ZN(_14565_)
  );
  AND2_X1 _49550_ (
    .A1(\cpuregs[2] [6]),
    .A2(_12705_),
    .ZN(_14566_)
  );
  INV_X1 _49551_ (
    .A(_14566_),
    .ZN(_14567_)
  );
  AND2_X1 _49552_ (
    .A1(_14565_),
    .A2(_14567_),
    .ZN(_14568_)
  );
  INV_X1 _49553_ (
    .A(_14568_),
    .ZN(_00812_)
  );
  AND2_X1 _49554_ (
    .A1(_12704_),
    .A2(_12971_),
    .ZN(_14569_)
  );
  INV_X1 _49555_ (
    .A(_14569_),
    .ZN(_14570_)
  );
  AND2_X1 _49556_ (
    .A1(_21544_),
    .A2(_12705_),
    .ZN(_14571_)
  );
  INV_X1 _49557_ (
    .A(_14571_),
    .ZN(_14572_)
  );
  AND2_X1 _49558_ (
    .A1(_14570_),
    .A2(_14572_),
    .ZN(_00813_)
  );
  AND2_X1 _49559_ (
    .A1(_12704_),
    .A2(_12986_),
    .ZN(_14573_)
  );
  INV_X1 _49560_ (
    .A(_14573_),
    .ZN(_14574_)
  );
  AND2_X1 _49561_ (
    .A1(_21545_),
    .A2(_12705_),
    .ZN(_14575_)
  );
  INV_X1 _49562_ (
    .A(_14575_),
    .ZN(_14576_)
  );
  AND2_X1 _49563_ (
    .A1(_14574_),
    .A2(_14576_),
    .ZN(_00814_)
  );
  AND2_X1 _49564_ (
    .A1(_12704_),
    .A2(_13001_),
    .ZN(_14577_)
  );
  INV_X1 _49565_ (
    .A(_14577_),
    .ZN(_14578_)
  );
  AND2_X1 _49566_ (
    .A1(_21546_),
    .A2(_12705_),
    .ZN(_14579_)
  );
  INV_X1 _49567_ (
    .A(_14579_),
    .ZN(_14580_)
  );
  AND2_X1 _49568_ (
    .A1(_14578_),
    .A2(_14580_),
    .ZN(_00815_)
  );
  AND2_X1 _49569_ (
    .A1(_12704_),
    .A2(_13016_),
    .ZN(_14581_)
  );
  INV_X1 _49570_ (
    .A(_14581_),
    .ZN(_14582_)
  );
  AND2_X1 _49571_ (
    .A1(_21547_),
    .A2(_12705_),
    .ZN(_14583_)
  );
  INV_X1 _49572_ (
    .A(_14583_),
    .ZN(_14584_)
  );
  AND2_X1 _49573_ (
    .A1(_14582_),
    .A2(_14584_),
    .ZN(_00816_)
  );
  AND2_X1 _49574_ (
    .A1(_12704_),
    .A2(_13031_),
    .ZN(_14585_)
  );
  INV_X1 _49575_ (
    .A(_14585_),
    .ZN(_14586_)
  );
  AND2_X1 _49576_ (
    .A1(_21548_),
    .A2(_12705_),
    .ZN(_14587_)
  );
  INV_X1 _49577_ (
    .A(_14587_),
    .ZN(_14588_)
  );
  AND2_X1 _49578_ (
    .A1(_14586_),
    .A2(_14588_),
    .ZN(_00817_)
  );
  AND2_X1 _49579_ (
    .A1(_12704_),
    .A2(_13046_),
    .ZN(_14589_)
  );
  INV_X1 _49580_ (
    .A(_14589_),
    .ZN(_14590_)
  );
  AND2_X1 _49581_ (
    .A1(_21549_),
    .A2(_12705_),
    .ZN(_14591_)
  );
  INV_X1 _49582_ (
    .A(_14591_),
    .ZN(_14592_)
  );
  AND2_X1 _49583_ (
    .A1(_14590_),
    .A2(_14592_),
    .ZN(_00818_)
  );
  AND2_X1 _49584_ (
    .A1(_12704_),
    .A2(_13061_),
    .ZN(_14593_)
  );
  INV_X1 _49585_ (
    .A(_14593_),
    .ZN(_14594_)
  );
  AND2_X1 _49586_ (
    .A1(_21550_),
    .A2(_12705_),
    .ZN(_14595_)
  );
  INV_X1 _49587_ (
    .A(_14595_),
    .ZN(_14596_)
  );
  AND2_X1 _49588_ (
    .A1(_14594_),
    .A2(_14596_),
    .ZN(_00819_)
  );
  AND2_X1 _49589_ (
    .A1(\cpuregs[2] [14]),
    .A2(_12705_),
    .ZN(_14597_)
  );
  INV_X1 _49590_ (
    .A(_14597_),
    .ZN(_14598_)
  );
  AND2_X1 _49591_ (
    .A1(_12704_),
    .A2(_13078_),
    .ZN(_14599_)
  );
  INV_X1 _49592_ (
    .A(_14599_),
    .ZN(_14600_)
  );
  AND2_X1 _49593_ (
    .A1(_14598_),
    .A2(_14600_),
    .ZN(_14601_)
  );
  INV_X1 _49594_ (
    .A(_14601_),
    .ZN(_00820_)
  );
  AND2_X1 _49595_ (
    .A1(_12704_),
    .A2(_13091_),
    .ZN(_14602_)
  );
  INV_X1 _49596_ (
    .A(_14602_),
    .ZN(_14603_)
  );
  AND2_X1 _49597_ (
    .A1(_21552_),
    .A2(_12705_),
    .ZN(_14604_)
  );
  INV_X1 _49598_ (
    .A(_14604_),
    .ZN(_14605_)
  );
  AND2_X1 _49599_ (
    .A1(_14603_),
    .A2(_14605_),
    .ZN(_00821_)
  );
  AND2_X1 _49600_ (
    .A1(\cpuregs[2] [16]),
    .A2(_12705_),
    .ZN(_14606_)
  );
  INV_X1 _49601_ (
    .A(_14606_),
    .ZN(_14607_)
  );
  AND2_X1 _49602_ (
    .A1(_12704_),
    .A2(_13108_),
    .ZN(_14608_)
  );
  INV_X1 _49603_ (
    .A(_14608_),
    .ZN(_14609_)
  );
  AND2_X1 _49604_ (
    .A1(_14607_),
    .A2(_14609_),
    .ZN(_14610_)
  );
  INV_X1 _49605_ (
    .A(_14610_),
    .ZN(_00822_)
  );
  AND2_X1 _49606_ (
    .A1(_12704_),
    .A2(_13121_),
    .ZN(_14611_)
  );
  INV_X1 _49607_ (
    .A(_14611_),
    .ZN(_14612_)
  );
  AND2_X1 _49608_ (
    .A1(_21554_),
    .A2(_12705_),
    .ZN(_14613_)
  );
  INV_X1 _49609_ (
    .A(_14613_),
    .ZN(_14614_)
  );
  AND2_X1 _49610_ (
    .A1(_14612_),
    .A2(_14614_),
    .ZN(_00823_)
  );
  AND2_X1 _49611_ (
    .A1(_12704_),
    .A2(_13139_),
    .ZN(_14615_)
  );
  INV_X1 _49612_ (
    .A(_14615_),
    .ZN(_14616_)
  );
  AND2_X1 _49613_ (
    .A1(\cpuregs[2] [18]),
    .A2(_12705_),
    .ZN(_14617_)
  );
  INV_X1 _49614_ (
    .A(_14617_),
    .ZN(_14618_)
  );
  AND2_X1 _49615_ (
    .A1(_14616_),
    .A2(_14618_),
    .ZN(_14619_)
  );
  INV_X1 _49616_ (
    .A(_14619_),
    .ZN(_00824_)
  );
  AND2_X1 _49617_ (
    .A1(_12704_),
    .A2(_13152_),
    .ZN(_14620_)
  );
  INV_X1 _49618_ (
    .A(_14620_),
    .ZN(_14621_)
  );
  AND2_X1 _49619_ (
    .A1(_21556_),
    .A2(_12705_),
    .ZN(_14622_)
  );
  INV_X1 _49620_ (
    .A(_14622_),
    .ZN(_14623_)
  );
  AND2_X1 _49621_ (
    .A1(_14621_),
    .A2(_14623_),
    .ZN(_00825_)
  );
  AND2_X1 _49622_ (
    .A1(_12704_),
    .A2(_13169_),
    .ZN(_14624_)
  );
  INV_X1 _49623_ (
    .A(_14624_),
    .ZN(_14625_)
  );
  AND2_X1 _49624_ (
    .A1(\cpuregs[2] [20]),
    .A2(_12705_),
    .ZN(_14626_)
  );
  INV_X1 _49625_ (
    .A(_14626_),
    .ZN(_14627_)
  );
  AND2_X1 _49626_ (
    .A1(_14625_),
    .A2(_14627_),
    .ZN(_14628_)
  );
  INV_X1 _49627_ (
    .A(_14628_),
    .ZN(_00826_)
  );
  AND2_X1 _49628_ (
    .A1(_12704_),
    .A2(_13182_),
    .ZN(_14629_)
  );
  INV_X1 _49629_ (
    .A(_14629_),
    .ZN(_14630_)
  );
  AND2_X1 _49630_ (
    .A1(_21557_),
    .A2(_12705_),
    .ZN(_14631_)
  );
  INV_X1 _49631_ (
    .A(_14631_),
    .ZN(_14632_)
  );
  AND2_X1 _49632_ (
    .A1(_14630_),
    .A2(_14632_),
    .ZN(_00827_)
  );
  AND2_X1 _49633_ (
    .A1(_12704_),
    .A2(_13197_),
    .ZN(_14633_)
  );
  INV_X1 _49634_ (
    .A(_14633_),
    .ZN(_14634_)
  );
  AND2_X1 _49635_ (
    .A1(_21558_),
    .A2(_12705_),
    .ZN(_14635_)
  );
  INV_X1 _49636_ (
    .A(_14635_),
    .ZN(_14636_)
  );
  AND2_X1 _49637_ (
    .A1(_14634_),
    .A2(_14636_),
    .ZN(_00828_)
  );
  AND2_X1 _49638_ (
    .A1(_12704_),
    .A2(_13212_),
    .ZN(_14637_)
  );
  INV_X1 _49639_ (
    .A(_14637_),
    .ZN(_14638_)
  );
  AND2_X1 _49640_ (
    .A1(_21559_),
    .A2(_12705_),
    .ZN(_14639_)
  );
  INV_X1 _49641_ (
    .A(_14639_),
    .ZN(_14640_)
  );
  AND2_X1 _49642_ (
    .A1(_14638_),
    .A2(_14640_),
    .ZN(_00829_)
  );
  AND2_X1 _49643_ (
    .A1(_12704_),
    .A2(_13227_),
    .ZN(_14641_)
  );
  INV_X1 _49644_ (
    .A(_14641_),
    .ZN(_14642_)
  );
  AND2_X1 _49645_ (
    .A1(_21560_),
    .A2(_12705_),
    .ZN(_14643_)
  );
  INV_X1 _49646_ (
    .A(_14643_),
    .ZN(_14644_)
  );
  AND2_X1 _49647_ (
    .A1(_14642_),
    .A2(_14644_),
    .ZN(_00830_)
  );
  AND2_X1 _49648_ (
    .A1(_12704_),
    .A2(_13242_),
    .ZN(_14645_)
  );
  INV_X1 _49649_ (
    .A(_14645_),
    .ZN(_14646_)
  );
  AND2_X1 _49650_ (
    .A1(_21561_),
    .A2(_12705_),
    .ZN(_14647_)
  );
  INV_X1 _49651_ (
    .A(_14647_),
    .ZN(_14648_)
  );
  AND2_X1 _49652_ (
    .A1(_14646_),
    .A2(_14648_),
    .ZN(_00831_)
  );
  AND2_X1 _49653_ (
    .A1(_12704_),
    .A2(_13257_),
    .ZN(_14649_)
  );
  INV_X1 _49654_ (
    .A(_14649_),
    .ZN(_14650_)
  );
  AND2_X1 _49655_ (
    .A1(_21562_),
    .A2(_12705_),
    .ZN(_14651_)
  );
  INV_X1 _49656_ (
    .A(_14651_),
    .ZN(_14652_)
  );
  AND2_X1 _49657_ (
    .A1(_14650_),
    .A2(_14652_),
    .ZN(_00832_)
  );
  AND2_X1 _49658_ (
    .A1(_12704_),
    .A2(_13272_),
    .ZN(_14653_)
  );
  INV_X1 _49659_ (
    .A(_14653_),
    .ZN(_14654_)
  );
  AND2_X1 _49660_ (
    .A1(_21563_),
    .A2(_12705_),
    .ZN(_14655_)
  );
  INV_X1 _49661_ (
    .A(_14655_),
    .ZN(_14656_)
  );
  AND2_X1 _49662_ (
    .A1(_14654_),
    .A2(_14656_),
    .ZN(_00833_)
  );
  AND2_X1 _49663_ (
    .A1(_12704_),
    .A2(_13287_),
    .ZN(_14657_)
  );
  INV_X1 _49664_ (
    .A(_14657_),
    .ZN(_14658_)
  );
  AND2_X1 _49665_ (
    .A1(_21564_),
    .A2(_12705_),
    .ZN(_14659_)
  );
  INV_X1 _49666_ (
    .A(_14659_),
    .ZN(_14660_)
  );
  AND2_X1 _49667_ (
    .A1(_14658_),
    .A2(_14660_),
    .ZN(_00834_)
  );
  AND2_X1 _49668_ (
    .A1(_12704_),
    .A2(_13302_),
    .ZN(_14661_)
  );
  INV_X1 _49669_ (
    .A(_14661_),
    .ZN(_14662_)
  );
  AND2_X1 _49670_ (
    .A1(_21565_),
    .A2(_12705_),
    .ZN(_14663_)
  );
  INV_X1 _49671_ (
    .A(_14663_),
    .ZN(_14664_)
  );
  AND2_X1 _49672_ (
    .A1(_14662_),
    .A2(_14664_),
    .ZN(_00835_)
  );
  AND2_X1 _49673_ (
    .A1(_12704_),
    .A2(_13317_),
    .ZN(_14665_)
  );
  INV_X1 _49674_ (
    .A(_14665_),
    .ZN(_14666_)
  );
  AND2_X1 _49675_ (
    .A1(_21566_),
    .A2(_12705_),
    .ZN(_14667_)
  );
  INV_X1 _49676_ (
    .A(_14667_),
    .ZN(_14668_)
  );
  AND2_X1 _49677_ (
    .A1(_14666_),
    .A2(_14668_),
    .ZN(_00836_)
  );
  AND2_X1 _49678_ (
    .A1(_12746_),
    .A2(_12874_),
    .ZN(_14669_)
  );
  INV_X1 _49679_ (
    .A(_14669_),
    .ZN(_14670_)
  );
  AND2_X1 _49680_ (
    .A1(\cpuregs[24] [0]),
    .A2(_12747_),
    .ZN(_14671_)
  );
  INV_X1 _49681_ (
    .A(_14671_),
    .ZN(_14672_)
  );
  AND2_X1 _49682_ (
    .A1(_14670_),
    .A2(_14672_),
    .ZN(_14673_)
  );
  INV_X1 _49683_ (
    .A(_14673_),
    .ZN(_00837_)
  );
  AND2_X1 _49684_ (
    .A1(_12746_),
    .A2(_12886_),
    .ZN(_14674_)
  );
  INV_X1 _49685_ (
    .A(_14674_),
    .ZN(_14675_)
  );
  AND2_X1 _49686_ (
    .A1(\cpuregs[24] [1]),
    .A2(_12747_),
    .ZN(_14676_)
  );
  INV_X1 _49687_ (
    .A(_14676_),
    .ZN(_14677_)
  );
  AND2_X1 _49688_ (
    .A1(_14675_),
    .A2(_14677_),
    .ZN(_14678_)
  );
  INV_X1 _49689_ (
    .A(_14678_),
    .ZN(_00838_)
  );
  AND2_X1 _49690_ (
    .A1(\cpuregs[24] [2]),
    .A2(_12747_),
    .ZN(_14679_)
  );
  INV_X1 _49691_ (
    .A(_14679_),
    .ZN(_14680_)
  );
  AND2_X1 _49692_ (
    .A1(_12746_),
    .A2(_12900_),
    .ZN(_14681_)
  );
  INV_X1 _49693_ (
    .A(_14681_),
    .ZN(_14682_)
  );
  AND2_X1 _49694_ (
    .A1(_14680_),
    .A2(_14682_),
    .ZN(_14683_)
  );
  INV_X1 _49695_ (
    .A(_14683_),
    .ZN(_00839_)
  );
  AND2_X1 _49696_ (
    .A1(_12746_),
    .A2(_12913_),
    .ZN(_14684_)
  );
  INV_X1 _49697_ (
    .A(_14684_),
    .ZN(_14685_)
  );
  AND2_X1 _49698_ (
    .A1(\cpuregs[24] [3]),
    .A2(_12747_),
    .ZN(_14686_)
  );
  INV_X1 _49699_ (
    .A(_14686_),
    .ZN(_14687_)
  );
  AND2_X1 _49700_ (
    .A1(_14685_),
    .A2(_14687_),
    .ZN(_14688_)
  );
  INV_X1 _49701_ (
    .A(_14688_),
    .ZN(_00840_)
  );
  AND2_X1 _49702_ (
    .A1(_12746_),
    .A2(_12928_),
    .ZN(_14689_)
  );
  INV_X1 _49703_ (
    .A(_14689_),
    .ZN(_14690_)
  );
  AND2_X1 _49704_ (
    .A1(\cpuregs[24] [4]),
    .A2(_12747_),
    .ZN(_14691_)
  );
  INV_X1 _49705_ (
    .A(_14691_),
    .ZN(_14692_)
  );
  AND2_X1 _49706_ (
    .A1(_14690_),
    .A2(_14692_),
    .ZN(_14693_)
  );
  INV_X1 _49707_ (
    .A(_14693_),
    .ZN(_00841_)
  );
  AND2_X1 _49708_ (
    .A1(_12746_),
    .A2(_12943_),
    .ZN(_14694_)
  );
  INV_X1 _49709_ (
    .A(_14694_),
    .ZN(_14695_)
  );
  AND2_X1 _49710_ (
    .A1(\cpuregs[24] [5]),
    .A2(_12747_),
    .ZN(_14696_)
  );
  INV_X1 _49711_ (
    .A(_14696_),
    .ZN(_14697_)
  );
  AND2_X1 _49712_ (
    .A1(_14695_),
    .A2(_14697_),
    .ZN(_14698_)
  );
  INV_X1 _49713_ (
    .A(_14698_),
    .ZN(_00842_)
  );
  AND2_X1 _49714_ (
    .A1(_12746_),
    .A2(_12958_),
    .ZN(_14699_)
  );
  INV_X1 _49715_ (
    .A(_14699_),
    .ZN(_14700_)
  );
  AND2_X1 _49716_ (
    .A1(\cpuregs[24] [6]),
    .A2(_12747_),
    .ZN(_14701_)
  );
  INV_X1 _49717_ (
    .A(_14701_),
    .ZN(_14702_)
  );
  AND2_X1 _49718_ (
    .A1(_14700_),
    .A2(_14702_),
    .ZN(_14703_)
  );
  INV_X1 _49719_ (
    .A(_14703_),
    .ZN(_00843_)
  );
  AND2_X1 _49720_ (
    .A1(_12746_),
    .A2(_12973_),
    .ZN(_14704_)
  );
  INV_X1 _49721_ (
    .A(_14704_),
    .ZN(_14705_)
  );
  AND2_X1 _49722_ (
    .A1(\cpuregs[24] [7]),
    .A2(_12747_),
    .ZN(_14706_)
  );
  INV_X1 _49723_ (
    .A(_14706_),
    .ZN(_14707_)
  );
  AND2_X1 _49724_ (
    .A1(_14705_),
    .A2(_14707_),
    .ZN(_14708_)
  );
  INV_X1 _49725_ (
    .A(_14708_),
    .ZN(_00844_)
  );
  AND2_X1 _49726_ (
    .A1(_12746_),
    .A2(_12988_),
    .ZN(_14709_)
  );
  INV_X1 _49727_ (
    .A(_14709_),
    .ZN(_14710_)
  );
  AND2_X1 _49728_ (
    .A1(\cpuregs[24] [8]),
    .A2(_12747_),
    .ZN(_14711_)
  );
  INV_X1 _49729_ (
    .A(_14711_),
    .ZN(_14712_)
  );
  AND2_X1 _49730_ (
    .A1(_14710_),
    .A2(_14712_),
    .ZN(_14713_)
  );
  INV_X1 _49731_ (
    .A(_14713_),
    .ZN(_00845_)
  );
  AND2_X1 _49732_ (
    .A1(_12746_),
    .A2(_13003_),
    .ZN(_14714_)
  );
  INV_X1 _49733_ (
    .A(_14714_),
    .ZN(_14715_)
  );
  AND2_X1 _49734_ (
    .A1(\cpuregs[24] [9]),
    .A2(_12747_),
    .ZN(_14716_)
  );
  INV_X1 _49735_ (
    .A(_14716_),
    .ZN(_14717_)
  );
  AND2_X1 _49736_ (
    .A1(_14715_),
    .A2(_14717_),
    .ZN(_14718_)
  );
  INV_X1 _49737_ (
    .A(_14718_),
    .ZN(_00846_)
  );
  AND2_X1 _49738_ (
    .A1(_12746_),
    .A2(_13018_),
    .ZN(_14719_)
  );
  INV_X1 _49739_ (
    .A(_14719_),
    .ZN(_14720_)
  );
  AND2_X1 _49740_ (
    .A1(\cpuregs[24] [10]),
    .A2(_12747_),
    .ZN(_14721_)
  );
  INV_X1 _49741_ (
    .A(_14721_),
    .ZN(_14722_)
  );
  AND2_X1 _49742_ (
    .A1(_14720_),
    .A2(_14722_),
    .ZN(_14723_)
  );
  INV_X1 _49743_ (
    .A(_14723_),
    .ZN(_00847_)
  );
  AND2_X1 _49744_ (
    .A1(_12746_),
    .A2(_13033_),
    .ZN(_14724_)
  );
  INV_X1 _49745_ (
    .A(_14724_),
    .ZN(_14725_)
  );
  AND2_X1 _49746_ (
    .A1(\cpuregs[24] [11]),
    .A2(_12747_),
    .ZN(_14726_)
  );
  INV_X1 _49747_ (
    .A(_14726_),
    .ZN(_14727_)
  );
  AND2_X1 _49748_ (
    .A1(_14725_),
    .A2(_14727_),
    .ZN(_14728_)
  );
  INV_X1 _49749_ (
    .A(_14728_),
    .ZN(_00848_)
  );
  AND2_X1 _49750_ (
    .A1(_12746_),
    .A2(_13048_),
    .ZN(_14729_)
  );
  INV_X1 _49751_ (
    .A(_14729_),
    .ZN(_14730_)
  );
  AND2_X1 _49752_ (
    .A1(\cpuregs[24] [12]),
    .A2(_12747_),
    .ZN(_14731_)
  );
  INV_X1 _49753_ (
    .A(_14731_),
    .ZN(_14732_)
  );
  AND2_X1 _49754_ (
    .A1(_14730_),
    .A2(_14732_),
    .ZN(_14733_)
  );
  INV_X1 _49755_ (
    .A(_14733_),
    .ZN(_00849_)
  );
  AND2_X1 _49756_ (
    .A1(_12746_),
    .A2(_13063_),
    .ZN(_14734_)
  );
  INV_X1 _49757_ (
    .A(_14734_),
    .ZN(_14735_)
  );
  AND2_X1 _49758_ (
    .A1(\cpuregs[24] [13]),
    .A2(_12747_),
    .ZN(_14736_)
  );
  INV_X1 _49759_ (
    .A(_14736_),
    .ZN(_14737_)
  );
  AND2_X1 _49760_ (
    .A1(_14735_),
    .A2(_14737_),
    .ZN(_14738_)
  );
  INV_X1 _49761_ (
    .A(_14738_),
    .ZN(_00850_)
  );
  AND2_X1 _49762_ (
    .A1(_12746_),
    .A2(_13078_),
    .ZN(_14739_)
  );
  INV_X1 _49763_ (
    .A(_14739_),
    .ZN(_14740_)
  );
  AND2_X1 _49764_ (
    .A1(\cpuregs[24] [14]),
    .A2(_12747_),
    .ZN(_14741_)
  );
  INV_X1 _49765_ (
    .A(_14741_),
    .ZN(_14742_)
  );
  AND2_X1 _49766_ (
    .A1(_14740_),
    .A2(_14742_),
    .ZN(_14743_)
  );
  INV_X1 _49767_ (
    .A(_14743_),
    .ZN(_00851_)
  );
  AND2_X1 _49768_ (
    .A1(_12746_),
    .A2(_13093_),
    .ZN(_14744_)
  );
  INV_X1 _49769_ (
    .A(_14744_),
    .ZN(_14745_)
  );
  AND2_X1 _49770_ (
    .A1(\cpuregs[24] [15]),
    .A2(_12747_),
    .ZN(_14746_)
  );
  INV_X1 _49771_ (
    .A(_14746_),
    .ZN(_14747_)
  );
  AND2_X1 _49772_ (
    .A1(_14745_),
    .A2(_14747_),
    .ZN(_14748_)
  );
  INV_X1 _49773_ (
    .A(_14748_),
    .ZN(_00852_)
  );
  AND2_X1 _49774_ (
    .A1(\cpuregs[24] [16]),
    .A2(_12747_),
    .ZN(_14749_)
  );
  INV_X1 _49775_ (
    .A(_14749_),
    .ZN(_14750_)
  );
  AND2_X1 _49776_ (
    .A1(_12746_),
    .A2(_13108_),
    .ZN(_14751_)
  );
  INV_X1 _49777_ (
    .A(_14751_),
    .ZN(_14752_)
  );
  AND2_X1 _49778_ (
    .A1(_14750_),
    .A2(_14752_),
    .ZN(_14753_)
  );
  INV_X1 _49779_ (
    .A(_14753_),
    .ZN(_00853_)
  );
  AND2_X1 _49780_ (
    .A1(_12746_),
    .A2(_13123_),
    .ZN(_14754_)
  );
  INV_X1 _49781_ (
    .A(_14754_),
    .ZN(_14755_)
  );
  AND2_X1 _49782_ (
    .A1(\cpuregs[24] [17]),
    .A2(_12747_),
    .ZN(_14756_)
  );
  INV_X1 _49783_ (
    .A(_14756_),
    .ZN(_14757_)
  );
  AND2_X1 _49784_ (
    .A1(_14755_),
    .A2(_14757_),
    .ZN(_14758_)
  );
  INV_X1 _49785_ (
    .A(_14758_),
    .ZN(_00854_)
  );
  AND2_X1 _49786_ (
    .A1(_12746_),
    .A2(_13139_),
    .ZN(_14759_)
  );
  INV_X1 _49787_ (
    .A(_14759_),
    .ZN(_14760_)
  );
  AND2_X1 _49788_ (
    .A1(\cpuregs[24] [18]),
    .A2(_12747_),
    .ZN(_14761_)
  );
  INV_X1 _49789_ (
    .A(_14761_),
    .ZN(_14762_)
  );
  AND2_X1 _49790_ (
    .A1(_14760_),
    .A2(_14762_),
    .ZN(_14763_)
  );
  INV_X1 _49791_ (
    .A(_14763_),
    .ZN(_00855_)
  );
  AND2_X1 _49792_ (
    .A1(_12746_),
    .A2(_13154_),
    .ZN(_14764_)
  );
  INV_X1 _49793_ (
    .A(_14764_),
    .ZN(_14765_)
  );
  AND2_X1 _49794_ (
    .A1(\cpuregs[24] [19]),
    .A2(_12747_),
    .ZN(_14766_)
  );
  INV_X1 _49795_ (
    .A(_14766_),
    .ZN(_14767_)
  );
  AND2_X1 _49796_ (
    .A1(_14765_),
    .A2(_14767_),
    .ZN(_14768_)
  );
  INV_X1 _49797_ (
    .A(_14768_),
    .ZN(_00856_)
  );
  AND2_X1 _49798_ (
    .A1(_12746_),
    .A2(_13169_),
    .ZN(_14769_)
  );
  INV_X1 _49799_ (
    .A(_14769_),
    .ZN(_14770_)
  );
  AND2_X1 _49800_ (
    .A1(\cpuregs[24] [20]),
    .A2(_12747_),
    .ZN(_14771_)
  );
  INV_X1 _49801_ (
    .A(_14771_),
    .ZN(_14772_)
  );
  AND2_X1 _49802_ (
    .A1(_14770_),
    .A2(_14772_),
    .ZN(_14773_)
  );
  INV_X1 _49803_ (
    .A(_14773_),
    .ZN(_00857_)
  );
  AND2_X1 _49804_ (
    .A1(_12746_),
    .A2(_13184_),
    .ZN(_14774_)
  );
  INV_X1 _49805_ (
    .A(_14774_),
    .ZN(_14775_)
  );
  AND2_X1 _49806_ (
    .A1(\cpuregs[24] [21]),
    .A2(_12747_),
    .ZN(_14776_)
  );
  INV_X1 _49807_ (
    .A(_14776_),
    .ZN(_14777_)
  );
  AND2_X1 _49808_ (
    .A1(_14775_),
    .A2(_14777_),
    .ZN(_14778_)
  );
  INV_X1 _49809_ (
    .A(_14778_),
    .ZN(_00858_)
  );
  AND2_X1 _49810_ (
    .A1(_12746_),
    .A2(_13199_),
    .ZN(_14779_)
  );
  INV_X1 _49811_ (
    .A(_14779_),
    .ZN(_14780_)
  );
  AND2_X1 _49812_ (
    .A1(\cpuregs[24] [22]),
    .A2(_12747_),
    .ZN(_14781_)
  );
  INV_X1 _49813_ (
    .A(_14781_),
    .ZN(_14782_)
  );
  AND2_X1 _49814_ (
    .A1(_14780_),
    .A2(_14782_),
    .ZN(_14783_)
  );
  INV_X1 _49815_ (
    .A(_14783_),
    .ZN(_00859_)
  );
  AND2_X1 _49816_ (
    .A1(_12746_),
    .A2(_13214_),
    .ZN(_14784_)
  );
  INV_X1 _49817_ (
    .A(_14784_),
    .ZN(_14785_)
  );
  AND2_X1 _49818_ (
    .A1(\cpuregs[24] [23]),
    .A2(_12747_),
    .ZN(_14786_)
  );
  INV_X1 _49819_ (
    .A(_14786_),
    .ZN(_14787_)
  );
  AND2_X1 _49820_ (
    .A1(_14785_),
    .A2(_14787_),
    .ZN(_14788_)
  );
  INV_X1 _49821_ (
    .A(_14788_),
    .ZN(_00860_)
  );
  AND2_X1 _49822_ (
    .A1(_12746_),
    .A2(_13229_),
    .ZN(_14789_)
  );
  INV_X1 _49823_ (
    .A(_14789_),
    .ZN(_14790_)
  );
  AND2_X1 _49824_ (
    .A1(\cpuregs[24] [24]),
    .A2(_12747_),
    .ZN(_14791_)
  );
  INV_X1 _49825_ (
    .A(_14791_),
    .ZN(_14792_)
  );
  AND2_X1 _49826_ (
    .A1(_14790_),
    .A2(_14792_),
    .ZN(_14793_)
  );
  INV_X1 _49827_ (
    .A(_14793_),
    .ZN(_00861_)
  );
  AND2_X1 _49828_ (
    .A1(_12746_),
    .A2(_13244_),
    .ZN(_14794_)
  );
  INV_X1 _49829_ (
    .A(_14794_),
    .ZN(_14795_)
  );
  AND2_X1 _49830_ (
    .A1(\cpuregs[24] [25]),
    .A2(_12747_),
    .ZN(_14796_)
  );
  INV_X1 _49831_ (
    .A(_14796_),
    .ZN(_14797_)
  );
  AND2_X1 _49832_ (
    .A1(_14795_),
    .A2(_14797_),
    .ZN(_14798_)
  );
  INV_X1 _49833_ (
    .A(_14798_),
    .ZN(_00862_)
  );
  AND2_X1 _49834_ (
    .A1(_12746_),
    .A2(_13259_),
    .ZN(_14799_)
  );
  INV_X1 _49835_ (
    .A(_14799_),
    .ZN(_14800_)
  );
  AND2_X1 _49836_ (
    .A1(\cpuregs[24] [26]),
    .A2(_12747_),
    .ZN(_14801_)
  );
  INV_X1 _49837_ (
    .A(_14801_),
    .ZN(_14802_)
  );
  AND2_X1 _49838_ (
    .A1(_14800_),
    .A2(_14802_),
    .ZN(_14803_)
  );
  INV_X1 _49839_ (
    .A(_14803_),
    .ZN(_00863_)
  );
  AND2_X1 _49840_ (
    .A1(_12746_),
    .A2(_13274_),
    .ZN(_14804_)
  );
  INV_X1 _49841_ (
    .A(_14804_),
    .ZN(_14805_)
  );
  AND2_X1 _49842_ (
    .A1(\cpuregs[24] [27]),
    .A2(_12747_),
    .ZN(_14806_)
  );
  INV_X1 _49843_ (
    .A(_14806_),
    .ZN(_14807_)
  );
  AND2_X1 _49844_ (
    .A1(_14805_),
    .A2(_14807_),
    .ZN(_14808_)
  );
  INV_X1 _49845_ (
    .A(_14808_),
    .ZN(_00864_)
  );
  AND2_X1 _49846_ (
    .A1(_12746_),
    .A2(_13289_),
    .ZN(_14809_)
  );
  INV_X1 _49847_ (
    .A(_14809_),
    .ZN(_14810_)
  );
  AND2_X1 _49848_ (
    .A1(\cpuregs[24] [28]),
    .A2(_12747_),
    .ZN(_14811_)
  );
  INV_X1 _49849_ (
    .A(_14811_),
    .ZN(_14812_)
  );
  AND2_X1 _49850_ (
    .A1(_14810_),
    .A2(_14812_),
    .ZN(_14813_)
  );
  INV_X1 _49851_ (
    .A(_14813_),
    .ZN(_00865_)
  );
  AND2_X1 _49852_ (
    .A1(_12746_),
    .A2(_13304_),
    .ZN(_14814_)
  );
  INV_X1 _49853_ (
    .A(_14814_),
    .ZN(_14815_)
  );
  AND2_X1 _49854_ (
    .A1(\cpuregs[24] [29]),
    .A2(_12747_),
    .ZN(_14816_)
  );
  INV_X1 _49855_ (
    .A(_14816_),
    .ZN(_14817_)
  );
  AND2_X1 _49856_ (
    .A1(_14815_),
    .A2(_14817_),
    .ZN(_14818_)
  );
  INV_X1 _49857_ (
    .A(_14818_),
    .ZN(_00866_)
  );
  AND2_X1 _49858_ (
    .A1(_12746_),
    .A2(_13319_),
    .ZN(_14819_)
  );
  INV_X1 _49859_ (
    .A(_14819_),
    .ZN(_14820_)
  );
  AND2_X1 _49860_ (
    .A1(\cpuregs[24] [30]),
    .A2(_12747_),
    .ZN(_14821_)
  );
  INV_X1 _49861_ (
    .A(_14821_),
    .ZN(_14822_)
  );
  AND2_X1 _49862_ (
    .A1(_14820_),
    .A2(_14822_),
    .ZN(_14823_)
  );
  INV_X1 _49863_ (
    .A(_14823_),
    .ZN(_00867_)
  );
  AND2_X1 _49864_ (
    .A1(_12849_),
    .A2(_12874_),
    .ZN(_14824_)
  );
  INV_X1 _49865_ (
    .A(_14824_),
    .ZN(_14825_)
  );
  AND2_X1 _49866_ (
    .A1(\cpuregs[11] [0]),
    .A2(_12850_),
    .ZN(_14826_)
  );
  INV_X1 _49867_ (
    .A(_14826_),
    .ZN(_14827_)
  );
  AND2_X1 _49868_ (
    .A1(_14825_),
    .A2(_14827_),
    .ZN(_14828_)
  );
  INV_X1 _49869_ (
    .A(_14828_),
    .ZN(_00868_)
  );
  AND2_X1 _49870_ (
    .A1(_12849_),
    .A2(_12886_),
    .ZN(_14829_)
  );
  INV_X1 _49871_ (
    .A(_14829_),
    .ZN(_14830_)
  );
  AND2_X1 _49872_ (
    .A1(\cpuregs[11] [1]),
    .A2(_12850_),
    .ZN(_14831_)
  );
  INV_X1 _49873_ (
    .A(_14831_),
    .ZN(_14832_)
  );
  AND2_X1 _49874_ (
    .A1(_14830_),
    .A2(_14832_),
    .ZN(_14833_)
  );
  INV_X1 _49875_ (
    .A(_14833_),
    .ZN(_00869_)
  );
  AND2_X1 _49876_ (
    .A1(_12849_),
    .A2(_12900_),
    .ZN(_14834_)
  );
  INV_X1 _49877_ (
    .A(_14834_),
    .ZN(_14835_)
  );
  AND2_X1 _49878_ (
    .A1(\cpuregs[11] [2]),
    .A2(_12850_),
    .ZN(_14836_)
  );
  INV_X1 _49879_ (
    .A(_14836_),
    .ZN(_14837_)
  );
  AND2_X1 _49880_ (
    .A1(_14835_),
    .A2(_14837_),
    .ZN(_14838_)
  );
  INV_X1 _49881_ (
    .A(_14838_),
    .ZN(_00870_)
  );
  AND2_X1 _49882_ (
    .A1(\cpuregs[11] [3]),
    .A2(_12850_),
    .ZN(_14839_)
  );
  INV_X1 _49883_ (
    .A(_14839_),
    .ZN(_14840_)
  );
  AND2_X1 _49884_ (
    .A1(_12849_),
    .A2(_12913_),
    .ZN(_14841_)
  );
  INV_X1 _49885_ (
    .A(_14841_),
    .ZN(_14842_)
  );
  AND2_X1 _49886_ (
    .A1(_14840_),
    .A2(_14842_),
    .ZN(_14843_)
  );
  INV_X1 _49887_ (
    .A(_14843_),
    .ZN(_00871_)
  );
  AND2_X1 _49888_ (
    .A1(_12849_),
    .A2(_12928_),
    .ZN(_14844_)
  );
  INV_X1 _49889_ (
    .A(_14844_),
    .ZN(_14845_)
  );
  AND2_X1 _49890_ (
    .A1(\cpuregs[11] [4]),
    .A2(_12850_),
    .ZN(_14846_)
  );
  INV_X1 _49891_ (
    .A(_14846_),
    .ZN(_14847_)
  );
  AND2_X1 _49892_ (
    .A1(_14845_),
    .A2(_14847_),
    .ZN(_14848_)
  );
  INV_X1 _49893_ (
    .A(_14848_),
    .ZN(_00872_)
  );
  AND2_X1 _49894_ (
    .A1(_12849_),
    .A2(_12943_),
    .ZN(_14849_)
  );
  INV_X1 _49895_ (
    .A(_14849_),
    .ZN(_14850_)
  );
  AND2_X1 _49896_ (
    .A1(\cpuregs[11] [5]),
    .A2(_12850_),
    .ZN(_14851_)
  );
  INV_X1 _49897_ (
    .A(_14851_),
    .ZN(_14852_)
  );
  AND2_X1 _49898_ (
    .A1(_14850_),
    .A2(_14852_),
    .ZN(_14853_)
  );
  INV_X1 _49899_ (
    .A(_14853_),
    .ZN(_00873_)
  );
  AND2_X1 _49900_ (
    .A1(_12849_),
    .A2(_12958_),
    .ZN(_14854_)
  );
  INV_X1 _49901_ (
    .A(_14854_),
    .ZN(_14855_)
  );
  AND2_X1 _49902_ (
    .A1(\cpuregs[11] [6]),
    .A2(_12850_),
    .ZN(_14856_)
  );
  INV_X1 _49903_ (
    .A(_14856_),
    .ZN(_14857_)
  );
  AND2_X1 _49904_ (
    .A1(_14855_),
    .A2(_14857_),
    .ZN(_14858_)
  );
  INV_X1 _49905_ (
    .A(_14858_),
    .ZN(_00874_)
  );
  AND2_X1 _49906_ (
    .A1(_12849_),
    .A2(_12973_),
    .ZN(_14859_)
  );
  INV_X1 _49907_ (
    .A(_14859_),
    .ZN(_14860_)
  );
  AND2_X1 _49908_ (
    .A1(\cpuregs[11] [7]),
    .A2(_12850_),
    .ZN(_14861_)
  );
  INV_X1 _49909_ (
    .A(_14861_),
    .ZN(_14862_)
  );
  AND2_X1 _49910_ (
    .A1(_14860_),
    .A2(_14862_),
    .ZN(_14863_)
  );
  INV_X1 _49911_ (
    .A(_14863_),
    .ZN(_00875_)
  );
  AND2_X1 _49912_ (
    .A1(_12849_),
    .A2(_12988_),
    .ZN(_14864_)
  );
  INV_X1 _49913_ (
    .A(_14864_),
    .ZN(_14865_)
  );
  AND2_X1 _49914_ (
    .A1(\cpuregs[11] [8]),
    .A2(_12850_),
    .ZN(_14866_)
  );
  INV_X1 _49915_ (
    .A(_14866_),
    .ZN(_14867_)
  );
  AND2_X1 _49916_ (
    .A1(_14865_),
    .A2(_14867_),
    .ZN(_14868_)
  );
  INV_X1 _49917_ (
    .A(_14868_),
    .ZN(_00876_)
  );
  AND2_X1 _49918_ (
    .A1(_12849_),
    .A2(_13003_),
    .ZN(_14869_)
  );
  INV_X1 _49919_ (
    .A(_14869_),
    .ZN(_14870_)
  );
  AND2_X1 _49920_ (
    .A1(\cpuregs[11] [9]),
    .A2(_12850_),
    .ZN(_14871_)
  );
  INV_X1 _49921_ (
    .A(_14871_),
    .ZN(_14872_)
  );
  AND2_X1 _49922_ (
    .A1(_14870_),
    .A2(_14872_),
    .ZN(_14873_)
  );
  INV_X1 _49923_ (
    .A(_14873_),
    .ZN(_00877_)
  );
  AND2_X1 _49924_ (
    .A1(_12849_),
    .A2(_13018_),
    .ZN(_14874_)
  );
  INV_X1 _49925_ (
    .A(_14874_),
    .ZN(_14875_)
  );
  AND2_X1 _49926_ (
    .A1(\cpuregs[11] [10]),
    .A2(_12850_),
    .ZN(_14876_)
  );
  INV_X1 _49927_ (
    .A(_14876_),
    .ZN(_14877_)
  );
  AND2_X1 _49928_ (
    .A1(_14875_),
    .A2(_14877_),
    .ZN(_14878_)
  );
  INV_X1 _49929_ (
    .A(_14878_),
    .ZN(_00878_)
  );
  AND2_X1 _49930_ (
    .A1(_12849_),
    .A2(_13033_),
    .ZN(_14879_)
  );
  INV_X1 _49931_ (
    .A(_14879_),
    .ZN(_14880_)
  );
  AND2_X1 _49932_ (
    .A1(\cpuregs[11] [11]),
    .A2(_12850_),
    .ZN(_14881_)
  );
  INV_X1 _49933_ (
    .A(_14881_),
    .ZN(_14882_)
  );
  AND2_X1 _49934_ (
    .A1(_14880_),
    .A2(_14882_),
    .ZN(_14883_)
  );
  INV_X1 _49935_ (
    .A(_14883_),
    .ZN(_00879_)
  );
  AND2_X1 _49936_ (
    .A1(_12849_),
    .A2(_13048_),
    .ZN(_14884_)
  );
  INV_X1 _49937_ (
    .A(_14884_),
    .ZN(_14885_)
  );
  AND2_X1 _49938_ (
    .A1(\cpuregs[11] [12]),
    .A2(_12850_),
    .ZN(_14886_)
  );
  INV_X1 _49939_ (
    .A(_14886_),
    .ZN(_14887_)
  );
  AND2_X1 _49940_ (
    .A1(_14885_),
    .A2(_14887_),
    .ZN(_14888_)
  );
  INV_X1 _49941_ (
    .A(_14888_),
    .ZN(_00880_)
  );
  AND2_X1 _49942_ (
    .A1(_12849_),
    .A2(_13063_),
    .ZN(_14889_)
  );
  INV_X1 _49943_ (
    .A(_14889_),
    .ZN(_14890_)
  );
  AND2_X1 _49944_ (
    .A1(\cpuregs[11] [13]),
    .A2(_12850_),
    .ZN(_14891_)
  );
  INV_X1 _49945_ (
    .A(_14891_),
    .ZN(_14892_)
  );
  AND2_X1 _49946_ (
    .A1(_14890_),
    .A2(_14892_),
    .ZN(_14893_)
  );
  INV_X1 _49947_ (
    .A(_14893_),
    .ZN(_00881_)
  );
  AND2_X1 _49948_ (
    .A1(_12849_),
    .A2(_13078_),
    .ZN(_14894_)
  );
  INV_X1 _49949_ (
    .A(_14894_),
    .ZN(_14895_)
  );
  AND2_X1 _49950_ (
    .A1(\cpuregs[11] [14]),
    .A2(_12850_),
    .ZN(_14896_)
  );
  INV_X1 _49951_ (
    .A(_14896_),
    .ZN(_14897_)
  );
  AND2_X1 _49952_ (
    .A1(_14895_),
    .A2(_14897_),
    .ZN(_14898_)
  );
  INV_X1 _49953_ (
    .A(_14898_),
    .ZN(_00882_)
  );
  AND2_X1 _49954_ (
    .A1(_12849_),
    .A2(_13093_),
    .ZN(_14899_)
  );
  INV_X1 _49955_ (
    .A(_14899_),
    .ZN(_14900_)
  );
  AND2_X1 _49956_ (
    .A1(\cpuregs[11] [15]),
    .A2(_12850_),
    .ZN(_14901_)
  );
  INV_X1 _49957_ (
    .A(_14901_),
    .ZN(_14902_)
  );
  AND2_X1 _49958_ (
    .A1(_14900_),
    .A2(_14902_),
    .ZN(_14903_)
  );
  INV_X1 _49959_ (
    .A(_14903_),
    .ZN(_00883_)
  );
  AND2_X1 _49960_ (
    .A1(_12849_),
    .A2(_13108_),
    .ZN(_14904_)
  );
  INV_X1 _49961_ (
    .A(_14904_),
    .ZN(_14905_)
  );
  AND2_X1 _49962_ (
    .A1(\cpuregs[11] [16]),
    .A2(_12850_),
    .ZN(_14906_)
  );
  INV_X1 _49963_ (
    .A(_14906_),
    .ZN(_14907_)
  );
  AND2_X1 _49964_ (
    .A1(_14905_),
    .A2(_14907_),
    .ZN(_14908_)
  );
  INV_X1 _49965_ (
    .A(_14908_),
    .ZN(_00884_)
  );
  AND2_X1 _49966_ (
    .A1(_12849_),
    .A2(_13123_),
    .ZN(_14909_)
  );
  INV_X1 _49967_ (
    .A(_14909_),
    .ZN(_14910_)
  );
  AND2_X1 _49968_ (
    .A1(\cpuregs[11] [17]),
    .A2(_12850_),
    .ZN(_14911_)
  );
  INV_X1 _49969_ (
    .A(_14911_),
    .ZN(_14912_)
  );
  AND2_X1 _49970_ (
    .A1(_14910_),
    .A2(_14912_),
    .ZN(_14913_)
  );
  INV_X1 _49971_ (
    .A(_14913_),
    .ZN(_00885_)
  );
  AND2_X1 _49972_ (
    .A1(_12849_),
    .A2(_13139_),
    .ZN(_14914_)
  );
  INV_X1 _49973_ (
    .A(_14914_),
    .ZN(_14915_)
  );
  AND2_X1 _49974_ (
    .A1(\cpuregs[11] [18]),
    .A2(_12850_),
    .ZN(_14916_)
  );
  INV_X1 _49975_ (
    .A(_14916_),
    .ZN(_14917_)
  );
  AND2_X1 _49976_ (
    .A1(_14915_),
    .A2(_14917_),
    .ZN(_14918_)
  );
  INV_X1 _49977_ (
    .A(_14918_),
    .ZN(_00886_)
  );
  AND2_X1 _49978_ (
    .A1(_12849_),
    .A2(_13154_),
    .ZN(_14919_)
  );
  INV_X1 _49979_ (
    .A(_14919_),
    .ZN(_14920_)
  );
  AND2_X1 _49980_ (
    .A1(\cpuregs[11] [19]),
    .A2(_12850_),
    .ZN(_14921_)
  );
  INV_X1 _49981_ (
    .A(_14921_),
    .ZN(_14922_)
  );
  AND2_X1 _49982_ (
    .A1(_14920_),
    .A2(_14922_),
    .ZN(_14923_)
  );
  INV_X1 _49983_ (
    .A(_14923_),
    .ZN(_00887_)
  );
  AND2_X1 _49984_ (
    .A1(_12849_),
    .A2(_13169_),
    .ZN(_14924_)
  );
  INV_X1 _49985_ (
    .A(_14924_),
    .ZN(_14925_)
  );
  AND2_X1 _49986_ (
    .A1(\cpuregs[11] [20]),
    .A2(_12850_),
    .ZN(_14926_)
  );
  INV_X1 _49987_ (
    .A(_14926_),
    .ZN(_14927_)
  );
  AND2_X1 _49988_ (
    .A1(_14925_),
    .A2(_14927_),
    .ZN(_14928_)
  );
  INV_X1 _49989_ (
    .A(_14928_),
    .ZN(_00888_)
  );
  AND2_X1 _49990_ (
    .A1(_12849_),
    .A2(_13184_),
    .ZN(_14929_)
  );
  INV_X1 _49991_ (
    .A(_14929_),
    .ZN(_14930_)
  );
  AND2_X1 _49992_ (
    .A1(\cpuregs[11] [21]),
    .A2(_12850_),
    .ZN(_14931_)
  );
  INV_X1 _49993_ (
    .A(_14931_),
    .ZN(_14932_)
  );
  AND2_X1 _49994_ (
    .A1(_14930_),
    .A2(_14932_),
    .ZN(_14933_)
  );
  INV_X1 _49995_ (
    .A(_14933_),
    .ZN(_00889_)
  );
  AND2_X1 _49996_ (
    .A1(_12849_),
    .A2(_13199_),
    .ZN(_14934_)
  );
  INV_X1 _49997_ (
    .A(_14934_),
    .ZN(_14935_)
  );
  AND2_X1 _49998_ (
    .A1(\cpuregs[11] [22]),
    .A2(_12850_),
    .ZN(_14936_)
  );
  INV_X1 _49999_ (
    .A(_14936_),
    .ZN(_14937_)
  );
  AND2_X1 _50000_ (
    .A1(_14935_),
    .A2(_14937_),
    .ZN(_14938_)
  );
  INV_X1 _50001_ (
    .A(_14938_),
    .ZN(_00890_)
  );
  AND2_X1 _50002_ (
    .A1(_12849_),
    .A2(_13214_),
    .ZN(_14939_)
  );
  INV_X1 _50003_ (
    .A(_14939_),
    .ZN(_14940_)
  );
  AND2_X1 _50004_ (
    .A1(\cpuregs[11] [23]),
    .A2(_12850_),
    .ZN(_14941_)
  );
  INV_X1 _50005_ (
    .A(_14941_),
    .ZN(_14942_)
  );
  AND2_X1 _50006_ (
    .A1(_14940_),
    .A2(_14942_),
    .ZN(_14943_)
  );
  INV_X1 _50007_ (
    .A(_14943_),
    .ZN(_00891_)
  );
  AND2_X1 _50008_ (
    .A1(_12849_),
    .A2(_13229_),
    .ZN(_14944_)
  );
  INV_X1 _50009_ (
    .A(_14944_),
    .ZN(_14945_)
  );
  AND2_X1 _50010_ (
    .A1(\cpuregs[11] [24]),
    .A2(_12850_),
    .ZN(_14946_)
  );
  INV_X1 _50011_ (
    .A(_14946_),
    .ZN(_14947_)
  );
  AND2_X1 _50012_ (
    .A1(_14945_),
    .A2(_14947_),
    .ZN(_14948_)
  );
  INV_X1 _50013_ (
    .A(_14948_),
    .ZN(_00892_)
  );
  AND2_X1 _50014_ (
    .A1(_12849_),
    .A2(_13244_),
    .ZN(_14949_)
  );
  INV_X1 _50015_ (
    .A(_14949_),
    .ZN(_14950_)
  );
  AND2_X1 _50016_ (
    .A1(\cpuregs[11] [25]),
    .A2(_12850_),
    .ZN(_14951_)
  );
  INV_X1 _50017_ (
    .A(_14951_),
    .ZN(_14952_)
  );
  AND2_X1 _50018_ (
    .A1(_14950_),
    .A2(_14952_),
    .ZN(_14953_)
  );
  INV_X1 _50019_ (
    .A(_14953_),
    .ZN(_00893_)
  );
  AND2_X1 _50020_ (
    .A1(_12849_),
    .A2(_13259_),
    .ZN(_14954_)
  );
  INV_X1 _50021_ (
    .A(_14954_),
    .ZN(_14955_)
  );
  AND2_X1 _50022_ (
    .A1(\cpuregs[11] [26]),
    .A2(_12850_),
    .ZN(_14956_)
  );
  INV_X1 _50023_ (
    .A(_14956_),
    .ZN(_14957_)
  );
  AND2_X1 _50024_ (
    .A1(_14955_),
    .A2(_14957_),
    .ZN(_14958_)
  );
  INV_X1 _50025_ (
    .A(_14958_),
    .ZN(_00894_)
  );
  AND2_X1 _50026_ (
    .A1(_12849_),
    .A2(_13274_),
    .ZN(_14959_)
  );
  INV_X1 _50027_ (
    .A(_14959_),
    .ZN(_14960_)
  );
  AND2_X1 _50028_ (
    .A1(\cpuregs[11] [27]),
    .A2(_12850_),
    .ZN(_14961_)
  );
  INV_X1 _50029_ (
    .A(_14961_),
    .ZN(_14962_)
  );
  AND2_X1 _50030_ (
    .A1(_14960_),
    .A2(_14962_),
    .ZN(_14963_)
  );
  INV_X1 _50031_ (
    .A(_14963_),
    .ZN(_00895_)
  );
  AND2_X1 _50032_ (
    .A1(_12849_),
    .A2(_13289_),
    .ZN(_14964_)
  );
  INV_X1 _50033_ (
    .A(_14964_),
    .ZN(_14965_)
  );
  AND2_X1 _50034_ (
    .A1(\cpuregs[11] [28]),
    .A2(_12850_),
    .ZN(_14966_)
  );
  INV_X1 _50035_ (
    .A(_14966_),
    .ZN(_14967_)
  );
  AND2_X1 _50036_ (
    .A1(_14965_),
    .A2(_14967_),
    .ZN(_14968_)
  );
  INV_X1 _50037_ (
    .A(_14968_),
    .ZN(_00896_)
  );
  AND2_X1 _50038_ (
    .A1(_12849_),
    .A2(_13304_),
    .ZN(_14969_)
  );
  INV_X1 _50039_ (
    .A(_14969_),
    .ZN(_14970_)
  );
  AND2_X1 _50040_ (
    .A1(\cpuregs[11] [29]),
    .A2(_12850_),
    .ZN(_14971_)
  );
  INV_X1 _50041_ (
    .A(_14971_),
    .ZN(_14972_)
  );
  AND2_X1 _50042_ (
    .A1(_14970_),
    .A2(_14972_),
    .ZN(_14973_)
  );
  INV_X1 _50043_ (
    .A(_14973_),
    .ZN(_00897_)
  );
  AND2_X1 _50044_ (
    .A1(_12849_),
    .A2(_13319_),
    .ZN(_14974_)
  );
  INV_X1 _50045_ (
    .A(_14974_),
    .ZN(_14975_)
  );
  AND2_X1 _50046_ (
    .A1(\cpuregs[11] [30]),
    .A2(_12850_),
    .ZN(_14976_)
  );
  INV_X1 _50047_ (
    .A(_14976_),
    .ZN(_14977_)
  );
  AND2_X1 _50048_ (
    .A1(_14975_),
    .A2(_14977_),
    .ZN(_14978_)
  );
  INV_X1 _50049_ (
    .A(_14978_),
    .ZN(_00898_)
  );
  AND2_X1 _50050_ (
    .A1(_12798_),
    .A2(_12872_),
    .ZN(_14979_)
  );
  INV_X1 _50051_ (
    .A(_14979_),
    .ZN(_14980_)
  );
  AND2_X1 _50052_ (
    .A1(_21590_),
    .A2(_12799_),
    .ZN(_14981_)
  );
  INV_X1 _50053_ (
    .A(_14981_),
    .ZN(_14982_)
  );
  AND2_X1 _50054_ (
    .A1(_14980_),
    .A2(_14982_),
    .ZN(_00899_)
  );
  AND2_X1 _50055_ (
    .A1(_12798_),
    .A2(_12884_),
    .ZN(_14983_)
  );
  INV_X1 _50056_ (
    .A(_14983_),
    .ZN(_14984_)
  );
  AND2_X1 _50057_ (
    .A1(_21591_),
    .A2(_12799_),
    .ZN(_14985_)
  );
  INV_X1 _50058_ (
    .A(_14985_),
    .ZN(_14986_)
  );
  AND2_X1 _50059_ (
    .A1(_14984_),
    .A2(_14986_),
    .ZN(_00900_)
  );
  AND2_X1 _50060_ (
    .A1(_12798_),
    .A2(_12898_),
    .ZN(_14987_)
  );
  INV_X1 _50061_ (
    .A(_14987_),
    .ZN(_14988_)
  );
  AND2_X1 _50062_ (
    .A1(_21592_),
    .A2(_12799_),
    .ZN(_14989_)
  );
  INV_X1 _50063_ (
    .A(_14989_),
    .ZN(_14990_)
  );
  AND2_X1 _50064_ (
    .A1(_14988_),
    .A2(_14990_),
    .ZN(_00901_)
  );
  AND2_X1 _50065_ (
    .A1(\cpuregs[18] [3]),
    .A2(_12799_),
    .ZN(_14991_)
  );
  INV_X1 _50066_ (
    .A(_14991_),
    .ZN(_14992_)
  );
  AND2_X1 _50067_ (
    .A1(_12798_),
    .A2(_12913_),
    .ZN(_14993_)
  );
  INV_X1 _50068_ (
    .A(_14993_),
    .ZN(_14994_)
  );
  AND2_X1 _50069_ (
    .A1(_14992_),
    .A2(_14994_),
    .ZN(_14995_)
  );
  INV_X1 _50070_ (
    .A(_14995_),
    .ZN(_00902_)
  );
  AND2_X1 _50071_ (
    .A1(_12798_),
    .A2(_12928_),
    .ZN(_14996_)
  );
  INV_X1 _50072_ (
    .A(_14996_),
    .ZN(_14997_)
  );
  AND2_X1 _50073_ (
    .A1(\cpuregs[18] [4]),
    .A2(_12799_),
    .ZN(_14998_)
  );
  INV_X1 _50074_ (
    .A(_14998_),
    .ZN(_14999_)
  );
  AND2_X1 _50075_ (
    .A1(_14997_),
    .A2(_14999_),
    .ZN(_15000_)
  );
  INV_X1 _50076_ (
    .A(_15000_),
    .ZN(_00903_)
  );
  AND2_X1 _50077_ (
    .A1(_12798_),
    .A2(_12941_),
    .ZN(_15001_)
  );
  INV_X1 _50078_ (
    .A(_15001_),
    .ZN(_15002_)
  );
  AND2_X1 _50079_ (
    .A1(_21595_),
    .A2(_12799_),
    .ZN(_15003_)
  );
  INV_X1 _50080_ (
    .A(_15003_),
    .ZN(_15004_)
  );
  AND2_X1 _50081_ (
    .A1(_15002_),
    .A2(_15004_),
    .ZN(_00904_)
  );
  AND2_X1 _50082_ (
    .A1(_12798_),
    .A2(_12958_),
    .ZN(_15005_)
  );
  INV_X1 _50083_ (
    .A(_15005_),
    .ZN(_15006_)
  );
  AND2_X1 _50084_ (
    .A1(\cpuregs[18] [6]),
    .A2(_12799_),
    .ZN(_15007_)
  );
  INV_X1 _50085_ (
    .A(_15007_),
    .ZN(_15008_)
  );
  AND2_X1 _50086_ (
    .A1(_15006_),
    .A2(_15008_),
    .ZN(_15009_)
  );
  INV_X1 _50087_ (
    .A(_15009_),
    .ZN(_00905_)
  );
  AND2_X1 _50088_ (
    .A1(_12798_),
    .A2(_12971_),
    .ZN(_15010_)
  );
  INV_X1 _50089_ (
    .A(_15010_),
    .ZN(_15011_)
  );
  AND2_X1 _50090_ (
    .A1(_21596_),
    .A2(_12799_),
    .ZN(_15012_)
  );
  INV_X1 _50091_ (
    .A(_15012_),
    .ZN(_15013_)
  );
  AND2_X1 _50092_ (
    .A1(_15011_),
    .A2(_15013_),
    .ZN(_00906_)
  );
  AND2_X1 _50093_ (
    .A1(_12798_),
    .A2(_12988_),
    .ZN(_15014_)
  );
  INV_X1 _50094_ (
    .A(_15014_),
    .ZN(_15015_)
  );
  AND2_X1 _50095_ (
    .A1(\cpuregs[18] [8]),
    .A2(_12799_),
    .ZN(_15016_)
  );
  INV_X1 _50096_ (
    .A(_15016_),
    .ZN(_15017_)
  );
  AND2_X1 _50097_ (
    .A1(_15015_),
    .A2(_15017_),
    .ZN(_15018_)
  );
  INV_X1 _50098_ (
    .A(_15018_),
    .ZN(_00907_)
  );
  AND2_X1 _50099_ (
    .A1(_12798_),
    .A2(_13001_),
    .ZN(_15019_)
  );
  INV_X1 _50100_ (
    .A(_15019_),
    .ZN(_15020_)
  );
  AND2_X1 _50101_ (
    .A1(_21597_),
    .A2(_12799_),
    .ZN(_15021_)
  );
  INV_X1 _50102_ (
    .A(_15021_),
    .ZN(_15022_)
  );
  AND2_X1 _50103_ (
    .A1(_15020_),
    .A2(_15022_),
    .ZN(_00908_)
  );
  AND2_X1 _50104_ (
    .A1(_12798_),
    .A2(_13016_),
    .ZN(_15023_)
  );
  INV_X1 _50105_ (
    .A(_15023_),
    .ZN(_15024_)
  );
  AND2_X1 _50106_ (
    .A1(_21598_),
    .A2(_12799_),
    .ZN(_15025_)
  );
  INV_X1 _50107_ (
    .A(_15025_),
    .ZN(_15026_)
  );
  AND2_X1 _50108_ (
    .A1(_15024_),
    .A2(_15026_),
    .ZN(_00909_)
  );
  AND2_X1 _50109_ (
    .A1(_12798_),
    .A2(_13033_),
    .ZN(_15027_)
  );
  INV_X1 _50110_ (
    .A(_15027_),
    .ZN(_15028_)
  );
  AND2_X1 _50111_ (
    .A1(\cpuregs[18] [11]),
    .A2(_12799_),
    .ZN(_15029_)
  );
  INV_X1 _50112_ (
    .A(_15029_),
    .ZN(_15030_)
  );
  AND2_X1 _50113_ (
    .A1(_15028_),
    .A2(_15030_),
    .ZN(_15031_)
  );
  INV_X1 _50114_ (
    .A(_15031_),
    .ZN(_00910_)
  );
  AND2_X1 _50115_ (
    .A1(_12798_),
    .A2(_13046_),
    .ZN(_15032_)
  );
  INV_X1 _50116_ (
    .A(_15032_),
    .ZN(_15033_)
  );
  AND2_X1 _50117_ (
    .A1(_21599_),
    .A2(_12799_),
    .ZN(_15034_)
  );
  INV_X1 _50118_ (
    .A(_15034_),
    .ZN(_15035_)
  );
  AND2_X1 _50119_ (
    .A1(_15033_),
    .A2(_15035_),
    .ZN(_00911_)
  );
  AND2_X1 _50120_ (
    .A1(_12798_),
    .A2(_13061_),
    .ZN(_15036_)
  );
  INV_X1 _50121_ (
    .A(_15036_),
    .ZN(_15037_)
  );
  AND2_X1 _50122_ (
    .A1(_21600_),
    .A2(_12799_),
    .ZN(_15038_)
  );
  INV_X1 _50123_ (
    .A(_15038_),
    .ZN(_15039_)
  );
  AND2_X1 _50124_ (
    .A1(_15037_),
    .A2(_15039_),
    .ZN(_00912_)
  );
  AND2_X1 _50125_ (
    .A1(\cpuregs[18] [14]),
    .A2(_12799_),
    .ZN(_15040_)
  );
  INV_X1 _50126_ (
    .A(_15040_),
    .ZN(_15041_)
  );
  AND2_X1 _50127_ (
    .A1(_12798_),
    .A2(_13078_),
    .ZN(_15042_)
  );
  INV_X1 _50128_ (
    .A(_15042_),
    .ZN(_15043_)
  );
  AND2_X1 _50129_ (
    .A1(_15041_),
    .A2(_15043_),
    .ZN(_15044_)
  );
  INV_X1 _50130_ (
    .A(_15044_),
    .ZN(_00913_)
  );
  AND2_X1 _50131_ (
    .A1(_12798_),
    .A2(_13091_),
    .ZN(_15045_)
  );
  INV_X1 _50132_ (
    .A(_15045_),
    .ZN(_15046_)
  );
  AND2_X1 _50133_ (
    .A1(_21602_),
    .A2(_12799_),
    .ZN(_15047_)
  );
  INV_X1 _50134_ (
    .A(_15047_),
    .ZN(_15048_)
  );
  AND2_X1 _50135_ (
    .A1(_15046_),
    .A2(_15048_),
    .ZN(_00914_)
  );
  AND2_X1 _50136_ (
    .A1(\cpuregs[18] [16]),
    .A2(_12799_),
    .ZN(_15049_)
  );
  INV_X1 _50137_ (
    .A(_15049_),
    .ZN(_15050_)
  );
  AND2_X1 _50138_ (
    .A1(_12798_),
    .A2(_13108_),
    .ZN(_15051_)
  );
  INV_X1 _50139_ (
    .A(_15051_),
    .ZN(_15052_)
  );
  AND2_X1 _50140_ (
    .A1(_15050_),
    .A2(_15052_),
    .ZN(_15053_)
  );
  INV_X1 _50141_ (
    .A(_15053_),
    .ZN(_00915_)
  );
  AND2_X1 _50142_ (
    .A1(_12798_),
    .A2(_13123_),
    .ZN(_15054_)
  );
  INV_X1 _50143_ (
    .A(_15054_),
    .ZN(_15055_)
  );
  AND2_X1 _50144_ (
    .A1(\cpuregs[18] [17]),
    .A2(_12799_),
    .ZN(_15056_)
  );
  INV_X1 _50145_ (
    .A(_15056_),
    .ZN(_15057_)
  );
  AND2_X1 _50146_ (
    .A1(_15055_),
    .A2(_15057_),
    .ZN(_15058_)
  );
  INV_X1 _50147_ (
    .A(_15058_),
    .ZN(_00916_)
  );
  AND2_X1 _50148_ (
    .A1(_12798_),
    .A2(_13139_),
    .ZN(_15059_)
  );
  INV_X1 _50149_ (
    .A(_15059_),
    .ZN(_15060_)
  );
  AND2_X1 _50150_ (
    .A1(\cpuregs[18] [18]),
    .A2(_12799_),
    .ZN(_15061_)
  );
  INV_X1 _50151_ (
    .A(_15061_),
    .ZN(_15062_)
  );
  AND2_X1 _50152_ (
    .A1(_15060_),
    .A2(_15062_),
    .ZN(_15063_)
  );
  INV_X1 _50153_ (
    .A(_15063_),
    .ZN(_00917_)
  );
  AND2_X1 _50154_ (
    .A1(_12798_),
    .A2(_13152_),
    .ZN(_15064_)
  );
  INV_X1 _50155_ (
    .A(_15064_),
    .ZN(_15065_)
  );
  AND2_X1 _50156_ (
    .A1(_21605_),
    .A2(_12799_),
    .ZN(_15066_)
  );
  INV_X1 _50157_ (
    .A(_15066_),
    .ZN(_15067_)
  );
  AND2_X1 _50158_ (
    .A1(_15065_),
    .A2(_15067_),
    .ZN(_00918_)
  );
  AND2_X1 _50159_ (
    .A1(_12798_),
    .A2(_13169_),
    .ZN(_15068_)
  );
  INV_X1 _50160_ (
    .A(_15068_),
    .ZN(_15069_)
  );
  AND2_X1 _50161_ (
    .A1(\cpuregs[18] [20]),
    .A2(_12799_),
    .ZN(_15070_)
  );
  INV_X1 _50162_ (
    .A(_15070_),
    .ZN(_15071_)
  );
  AND2_X1 _50163_ (
    .A1(_15069_),
    .A2(_15071_),
    .ZN(_15072_)
  );
  INV_X1 _50164_ (
    .A(_15072_),
    .ZN(_00919_)
  );
  AND2_X1 _50165_ (
    .A1(_12798_),
    .A2(_13184_),
    .ZN(_15073_)
  );
  INV_X1 _50166_ (
    .A(_15073_),
    .ZN(_15074_)
  );
  AND2_X1 _50167_ (
    .A1(\cpuregs[18] [21]),
    .A2(_12799_),
    .ZN(_15075_)
  );
  INV_X1 _50168_ (
    .A(_15075_),
    .ZN(_15076_)
  );
  AND2_X1 _50169_ (
    .A1(_15074_),
    .A2(_15076_),
    .ZN(_15077_)
  );
  INV_X1 _50170_ (
    .A(_15077_),
    .ZN(_00920_)
  );
  AND2_X1 _50171_ (
    .A1(_12798_),
    .A2(_13199_),
    .ZN(_15078_)
  );
  INV_X1 _50172_ (
    .A(_15078_),
    .ZN(_15079_)
  );
  AND2_X1 _50173_ (
    .A1(\cpuregs[18] [22]),
    .A2(_12799_),
    .ZN(_15080_)
  );
  INV_X1 _50174_ (
    .A(_15080_),
    .ZN(_15081_)
  );
  AND2_X1 _50175_ (
    .A1(_15079_),
    .A2(_15081_),
    .ZN(_15082_)
  );
  INV_X1 _50176_ (
    .A(_15082_),
    .ZN(_00921_)
  );
  AND2_X1 _50177_ (
    .A1(_12798_),
    .A2(_13212_),
    .ZN(_15083_)
  );
  INV_X1 _50178_ (
    .A(_15083_),
    .ZN(_15084_)
  );
  AND2_X1 _50179_ (
    .A1(_21608_),
    .A2(_12799_),
    .ZN(_15085_)
  );
  INV_X1 _50180_ (
    .A(_15085_),
    .ZN(_15086_)
  );
  AND2_X1 _50181_ (
    .A1(_15084_),
    .A2(_15086_),
    .ZN(_00922_)
  );
  AND2_X1 _50182_ (
    .A1(_12798_),
    .A2(_13229_),
    .ZN(_15087_)
  );
  INV_X1 _50183_ (
    .A(_15087_),
    .ZN(_15088_)
  );
  AND2_X1 _50184_ (
    .A1(\cpuregs[18] [24]),
    .A2(_12799_),
    .ZN(_15089_)
  );
  INV_X1 _50185_ (
    .A(_15089_),
    .ZN(_15090_)
  );
  AND2_X1 _50186_ (
    .A1(_15088_),
    .A2(_15090_),
    .ZN(_15091_)
  );
  INV_X1 _50187_ (
    .A(_15091_),
    .ZN(_00923_)
  );
  AND2_X1 _50188_ (
    .A1(_12798_),
    .A2(_13242_),
    .ZN(_15092_)
  );
  INV_X1 _50189_ (
    .A(_15092_),
    .ZN(_15093_)
  );
  AND2_X1 _50190_ (
    .A1(_21610_),
    .A2(_12799_),
    .ZN(_15094_)
  );
  INV_X1 _50191_ (
    .A(_15094_),
    .ZN(_15095_)
  );
  AND2_X1 _50192_ (
    .A1(_15093_),
    .A2(_15095_),
    .ZN(_00924_)
  );
  AND2_X1 _50193_ (
    .A1(_12798_),
    .A2(_13259_),
    .ZN(_15096_)
  );
  INV_X1 _50194_ (
    .A(_15096_),
    .ZN(_15097_)
  );
  AND2_X1 _50195_ (
    .A1(\cpuregs[18] [26]),
    .A2(_12799_),
    .ZN(_15098_)
  );
  INV_X1 _50196_ (
    .A(_15098_),
    .ZN(_15099_)
  );
  AND2_X1 _50197_ (
    .A1(_15097_),
    .A2(_15099_),
    .ZN(_15100_)
  );
  INV_X1 _50198_ (
    .A(_15100_),
    .ZN(_00925_)
  );
  AND2_X1 _50199_ (
    .A1(_12798_),
    .A2(_13272_),
    .ZN(_15101_)
  );
  INV_X1 _50200_ (
    .A(_15101_),
    .ZN(_15102_)
  );
  AND2_X1 _50201_ (
    .A1(_21612_),
    .A2(_12799_),
    .ZN(_15103_)
  );
  INV_X1 _50202_ (
    .A(_15103_),
    .ZN(_15104_)
  );
  AND2_X1 _50203_ (
    .A1(_15102_),
    .A2(_15104_),
    .ZN(_00926_)
  );
  AND2_X1 _50204_ (
    .A1(_12798_),
    .A2(_13289_),
    .ZN(_15105_)
  );
  INV_X1 _50205_ (
    .A(_15105_),
    .ZN(_15106_)
  );
  AND2_X1 _50206_ (
    .A1(\cpuregs[18] [28]),
    .A2(_12799_),
    .ZN(_15107_)
  );
  INV_X1 _50207_ (
    .A(_15107_),
    .ZN(_15108_)
  );
  AND2_X1 _50208_ (
    .A1(_15106_),
    .A2(_15108_),
    .ZN(_15109_)
  );
  INV_X1 _50209_ (
    .A(_15109_),
    .ZN(_00927_)
  );
  AND2_X1 _50210_ (
    .A1(_12798_),
    .A2(_13302_),
    .ZN(_15110_)
  );
  INV_X1 _50211_ (
    .A(_15110_),
    .ZN(_15111_)
  );
  AND2_X1 _50212_ (
    .A1(_21614_),
    .A2(_12799_),
    .ZN(_15112_)
  );
  INV_X1 _50213_ (
    .A(_15112_),
    .ZN(_15113_)
  );
  AND2_X1 _50214_ (
    .A1(_15111_),
    .A2(_15113_),
    .ZN(_00928_)
  );
  AND2_X1 _50215_ (
    .A1(_12798_),
    .A2(_13317_),
    .ZN(_15114_)
  );
  INV_X1 _50216_ (
    .A(_15114_),
    .ZN(_15115_)
  );
  AND2_X1 _50217_ (
    .A1(_21615_),
    .A2(_12799_),
    .ZN(_15116_)
  );
  INV_X1 _50218_ (
    .A(_15116_),
    .ZN(_15117_)
  );
  AND2_X1 _50219_ (
    .A1(_15115_),
    .A2(_15117_),
    .ZN(_00929_)
  );
  AND2_X1 _50220_ (
    .A1(_12791_),
    .A2(_12874_),
    .ZN(_15118_)
  );
  INV_X1 _50221_ (
    .A(_15118_),
    .ZN(_15119_)
  );
  AND2_X1 _50222_ (
    .A1(\cpuregs[19] [0]),
    .A2(_12792_),
    .ZN(_15120_)
  );
  INV_X1 _50223_ (
    .A(_15120_),
    .ZN(_15121_)
  );
  AND2_X1 _50224_ (
    .A1(_15119_),
    .A2(_15121_),
    .ZN(_15122_)
  );
  INV_X1 _50225_ (
    .A(_15122_),
    .ZN(_00930_)
  );
  AND2_X1 _50226_ (
    .A1(\cpuregs[19] [1]),
    .A2(_12792_),
    .ZN(_15123_)
  );
  INV_X1 _50227_ (
    .A(_15123_),
    .ZN(_15124_)
  );
  AND2_X1 _50228_ (
    .A1(_12791_),
    .A2(_12886_),
    .ZN(_15125_)
  );
  INV_X1 _50229_ (
    .A(_15125_),
    .ZN(_15126_)
  );
  AND2_X1 _50230_ (
    .A1(_15124_),
    .A2(_15126_),
    .ZN(_15127_)
  );
  INV_X1 _50231_ (
    .A(_15127_),
    .ZN(_00931_)
  );
  AND2_X1 _50232_ (
    .A1(_12791_),
    .A2(_12900_),
    .ZN(_15128_)
  );
  INV_X1 _50233_ (
    .A(_15128_),
    .ZN(_15129_)
  );
  AND2_X1 _50234_ (
    .A1(\cpuregs[19] [2]),
    .A2(_12792_),
    .ZN(_15130_)
  );
  INV_X1 _50235_ (
    .A(_15130_),
    .ZN(_15131_)
  );
  AND2_X1 _50236_ (
    .A1(_15129_),
    .A2(_15131_),
    .ZN(_15132_)
  );
  INV_X1 _50237_ (
    .A(_15132_),
    .ZN(_00932_)
  );
  AND2_X1 _50238_ (
    .A1(_12791_),
    .A2(_12913_),
    .ZN(_15133_)
  );
  INV_X1 _50239_ (
    .A(_15133_),
    .ZN(_15134_)
  );
  AND2_X1 _50240_ (
    .A1(\cpuregs[19] [3]),
    .A2(_12792_),
    .ZN(_15135_)
  );
  INV_X1 _50241_ (
    .A(_15135_),
    .ZN(_15136_)
  );
  AND2_X1 _50242_ (
    .A1(_15134_),
    .A2(_15136_),
    .ZN(_15137_)
  );
  INV_X1 _50243_ (
    .A(_15137_),
    .ZN(_00933_)
  );
  AND2_X1 _50244_ (
    .A1(_12791_),
    .A2(_12928_),
    .ZN(_15138_)
  );
  INV_X1 _50245_ (
    .A(_15138_),
    .ZN(_15139_)
  );
  AND2_X1 _50246_ (
    .A1(\cpuregs[19] [4]),
    .A2(_12792_),
    .ZN(_15140_)
  );
  INV_X1 _50247_ (
    .A(_15140_),
    .ZN(_15141_)
  );
  AND2_X1 _50248_ (
    .A1(_15139_),
    .A2(_15141_),
    .ZN(_15142_)
  );
  INV_X1 _50249_ (
    .A(_15142_),
    .ZN(_00934_)
  );
  AND2_X1 _50250_ (
    .A1(_12791_),
    .A2(_12943_),
    .ZN(_15143_)
  );
  INV_X1 _50251_ (
    .A(_15143_),
    .ZN(_15144_)
  );
  AND2_X1 _50252_ (
    .A1(\cpuregs[19] [5]),
    .A2(_12792_),
    .ZN(_15145_)
  );
  INV_X1 _50253_ (
    .A(_15145_),
    .ZN(_15146_)
  );
  AND2_X1 _50254_ (
    .A1(_15144_),
    .A2(_15146_),
    .ZN(_15147_)
  );
  INV_X1 _50255_ (
    .A(_15147_),
    .ZN(_00935_)
  );
  AND2_X1 _50256_ (
    .A1(_12791_),
    .A2(_12958_),
    .ZN(_15148_)
  );
  INV_X1 _50257_ (
    .A(_15148_),
    .ZN(_15149_)
  );
  AND2_X1 _50258_ (
    .A1(\cpuregs[19] [6]),
    .A2(_12792_),
    .ZN(_15150_)
  );
  INV_X1 _50259_ (
    .A(_15150_),
    .ZN(_15151_)
  );
  AND2_X1 _50260_ (
    .A1(_15149_),
    .A2(_15151_),
    .ZN(_15152_)
  );
  INV_X1 _50261_ (
    .A(_15152_),
    .ZN(_00936_)
  );
  AND2_X1 _50262_ (
    .A1(_12791_),
    .A2(_12973_),
    .ZN(_15153_)
  );
  INV_X1 _50263_ (
    .A(_15153_),
    .ZN(_15154_)
  );
  AND2_X1 _50264_ (
    .A1(\cpuregs[19] [7]),
    .A2(_12792_),
    .ZN(_15155_)
  );
  INV_X1 _50265_ (
    .A(_15155_),
    .ZN(_15156_)
  );
  AND2_X1 _50266_ (
    .A1(_15154_),
    .A2(_15156_),
    .ZN(_15157_)
  );
  INV_X1 _50267_ (
    .A(_15157_),
    .ZN(_00937_)
  );
  AND2_X1 _50268_ (
    .A1(_12791_),
    .A2(_12988_),
    .ZN(_15158_)
  );
  INV_X1 _50269_ (
    .A(_15158_),
    .ZN(_15159_)
  );
  AND2_X1 _50270_ (
    .A1(\cpuregs[19] [8]),
    .A2(_12792_),
    .ZN(_15160_)
  );
  INV_X1 _50271_ (
    .A(_15160_),
    .ZN(_15161_)
  );
  AND2_X1 _50272_ (
    .A1(_15159_),
    .A2(_15161_),
    .ZN(_15162_)
  );
  INV_X1 _50273_ (
    .A(_15162_),
    .ZN(_00938_)
  );
  AND2_X1 _50274_ (
    .A1(_12791_),
    .A2(_13003_),
    .ZN(_15163_)
  );
  INV_X1 _50275_ (
    .A(_15163_),
    .ZN(_15164_)
  );
  AND2_X1 _50276_ (
    .A1(\cpuregs[19] [9]),
    .A2(_12792_),
    .ZN(_15165_)
  );
  INV_X1 _50277_ (
    .A(_15165_),
    .ZN(_15166_)
  );
  AND2_X1 _50278_ (
    .A1(_15164_),
    .A2(_15166_),
    .ZN(_15167_)
  );
  INV_X1 _50279_ (
    .A(_15167_),
    .ZN(_00939_)
  );
  AND2_X1 _50280_ (
    .A1(_12791_),
    .A2(_13018_),
    .ZN(_15168_)
  );
  INV_X1 _50281_ (
    .A(_15168_),
    .ZN(_15169_)
  );
  AND2_X1 _50282_ (
    .A1(\cpuregs[19] [10]),
    .A2(_12792_),
    .ZN(_15170_)
  );
  INV_X1 _50283_ (
    .A(_15170_),
    .ZN(_15171_)
  );
  AND2_X1 _50284_ (
    .A1(_15169_),
    .A2(_15171_),
    .ZN(_15172_)
  );
  INV_X1 _50285_ (
    .A(_15172_),
    .ZN(_00940_)
  );
  AND2_X1 _50286_ (
    .A1(_12791_),
    .A2(_13033_),
    .ZN(_15173_)
  );
  INV_X1 _50287_ (
    .A(_15173_),
    .ZN(_15174_)
  );
  AND2_X1 _50288_ (
    .A1(\cpuregs[19] [11]),
    .A2(_12792_),
    .ZN(_15175_)
  );
  INV_X1 _50289_ (
    .A(_15175_),
    .ZN(_15176_)
  );
  AND2_X1 _50290_ (
    .A1(_15174_),
    .A2(_15176_),
    .ZN(_15177_)
  );
  INV_X1 _50291_ (
    .A(_15177_),
    .ZN(_00941_)
  );
  AND2_X1 _50292_ (
    .A1(_12791_),
    .A2(_13048_),
    .ZN(_15178_)
  );
  INV_X1 _50293_ (
    .A(_15178_),
    .ZN(_15179_)
  );
  AND2_X1 _50294_ (
    .A1(\cpuregs[19] [12]),
    .A2(_12792_),
    .ZN(_15180_)
  );
  INV_X1 _50295_ (
    .A(_15180_),
    .ZN(_15181_)
  );
  AND2_X1 _50296_ (
    .A1(_15179_),
    .A2(_15181_),
    .ZN(_15182_)
  );
  INV_X1 _50297_ (
    .A(_15182_),
    .ZN(_00942_)
  );
  AND2_X1 _50298_ (
    .A1(_12791_),
    .A2(_13063_),
    .ZN(_15183_)
  );
  INV_X1 _50299_ (
    .A(_15183_),
    .ZN(_15184_)
  );
  AND2_X1 _50300_ (
    .A1(\cpuregs[19] [13]),
    .A2(_12792_),
    .ZN(_15185_)
  );
  INV_X1 _50301_ (
    .A(_15185_),
    .ZN(_15186_)
  );
  AND2_X1 _50302_ (
    .A1(_15184_),
    .A2(_15186_),
    .ZN(_15187_)
  );
  INV_X1 _50303_ (
    .A(_15187_),
    .ZN(_00943_)
  );
  AND2_X1 _50304_ (
    .A1(\cpuregs[19] [14]),
    .A2(_12792_),
    .ZN(_15188_)
  );
  INV_X1 _50305_ (
    .A(_15188_),
    .ZN(_15189_)
  );
  AND2_X1 _50306_ (
    .A1(_12791_),
    .A2(_13078_),
    .ZN(_15190_)
  );
  INV_X1 _50307_ (
    .A(_15190_),
    .ZN(_15191_)
  );
  AND2_X1 _50308_ (
    .A1(_15189_),
    .A2(_15191_),
    .ZN(_15192_)
  );
  INV_X1 _50309_ (
    .A(_15192_),
    .ZN(_00944_)
  );
  AND2_X1 _50310_ (
    .A1(_12791_),
    .A2(_13093_),
    .ZN(_15193_)
  );
  INV_X1 _50311_ (
    .A(_15193_),
    .ZN(_15194_)
  );
  AND2_X1 _50312_ (
    .A1(\cpuregs[19] [15]),
    .A2(_12792_),
    .ZN(_15195_)
  );
  INV_X1 _50313_ (
    .A(_15195_),
    .ZN(_15196_)
  );
  AND2_X1 _50314_ (
    .A1(_15194_),
    .A2(_15196_),
    .ZN(_15197_)
  );
  INV_X1 _50315_ (
    .A(_15197_),
    .ZN(_00945_)
  );
  AND2_X1 _50316_ (
    .A1(_12791_),
    .A2(_13108_),
    .ZN(_15198_)
  );
  INV_X1 _50317_ (
    .A(_15198_),
    .ZN(_15199_)
  );
  AND2_X1 _50318_ (
    .A1(\cpuregs[19] [16]),
    .A2(_12792_),
    .ZN(_15200_)
  );
  INV_X1 _50319_ (
    .A(_15200_),
    .ZN(_15201_)
  );
  AND2_X1 _50320_ (
    .A1(_15199_),
    .A2(_15201_),
    .ZN(_15202_)
  );
  INV_X1 _50321_ (
    .A(_15202_),
    .ZN(_00946_)
  );
  AND2_X1 _50322_ (
    .A1(_12791_),
    .A2(_13123_),
    .ZN(_15203_)
  );
  INV_X1 _50323_ (
    .A(_15203_),
    .ZN(_15204_)
  );
  AND2_X1 _50324_ (
    .A1(\cpuregs[19] [17]),
    .A2(_12792_),
    .ZN(_15205_)
  );
  INV_X1 _50325_ (
    .A(_15205_),
    .ZN(_15206_)
  );
  AND2_X1 _50326_ (
    .A1(_15204_),
    .A2(_15206_),
    .ZN(_15207_)
  );
  INV_X1 _50327_ (
    .A(_15207_),
    .ZN(_00947_)
  );
  AND2_X1 _50328_ (
    .A1(_12791_),
    .A2(_13139_),
    .ZN(_15208_)
  );
  INV_X1 _50329_ (
    .A(_15208_),
    .ZN(_15209_)
  );
  AND2_X1 _50330_ (
    .A1(\cpuregs[19] [18]),
    .A2(_12792_),
    .ZN(_15210_)
  );
  INV_X1 _50331_ (
    .A(_15210_),
    .ZN(_15211_)
  );
  AND2_X1 _50332_ (
    .A1(_15209_),
    .A2(_15211_),
    .ZN(_15212_)
  );
  INV_X1 _50333_ (
    .A(_15212_),
    .ZN(_00948_)
  );
  AND2_X1 _50334_ (
    .A1(_12791_),
    .A2(_13154_),
    .ZN(_15213_)
  );
  INV_X1 _50335_ (
    .A(_15213_),
    .ZN(_15214_)
  );
  AND2_X1 _50336_ (
    .A1(\cpuregs[19] [19]),
    .A2(_12792_),
    .ZN(_15215_)
  );
  INV_X1 _50337_ (
    .A(_15215_),
    .ZN(_15216_)
  );
  AND2_X1 _50338_ (
    .A1(_15214_),
    .A2(_15216_),
    .ZN(_15217_)
  );
  INV_X1 _50339_ (
    .A(_15217_),
    .ZN(_00949_)
  );
  AND2_X1 _50340_ (
    .A1(_12791_),
    .A2(_13169_),
    .ZN(_15218_)
  );
  INV_X1 _50341_ (
    .A(_15218_),
    .ZN(_15219_)
  );
  AND2_X1 _50342_ (
    .A1(\cpuregs[19] [20]),
    .A2(_12792_),
    .ZN(_15220_)
  );
  INV_X1 _50343_ (
    .A(_15220_),
    .ZN(_15221_)
  );
  AND2_X1 _50344_ (
    .A1(_15219_),
    .A2(_15221_),
    .ZN(_15222_)
  );
  INV_X1 _50345_ (
    .A(_15222_),
    .ZN(_00950_)
  );
  AND2_X1 _50346_ (
    .A1(_12791_),
    .A2(_13184_),
    .ZN(_15223_)
  );
  INV_X1 _50347_ (
    .A(_15223_),
    .ZN(_15224_)
  );
  AND2_X1 _50348_ (
    .A1(\cpuregs[19] [21]),
    .A2(_12792_),
    .ZN(_15225_)
  );
  INV_X1 _50349_ (
    .A(_15225_),
    .ZN(_15226_)
  );
  AND2_X1 _50350_ (
    .A1(_15224_),
    .A2(_15226_),
    .ZN(_15227_)
  );
  INV_X1 _50351_ (
    .A(_15227_),
    .ZN(_00951_)
  );
  AND2_X1 _50352_ (
    .A1(_12791_),
    .A2(_13199_),
    .ZN(_15228_)
  );
  INV_X1 _50353_ (
    .A(_15228_),
    .ZN(_15229_)
  );
  AND2_X1 _50354_ (
    .A1(\cpuregs[19] [22]),
    .A2(_12792_),
    .ZN(_15230_)
  );
  INV_X1 _50355_ (
    .A(_15230_),
    .ZN(_15231_)
  );
  AND2_X1 _50356_ (
    .A1(_15229_),
    .A2(_15231_),
    .ZN(_15232_)
  );
  INV_X1 _50357_ (
    .A(_15232_),
    .ZN(_00952_)
  );
  AND2_X1 _50358_ (
    .A1(_12791_),
    .A2(_13214_),
    .ZN(_15233_)
  );
  INV_X1 _50359_ (
    .A(_15233_),
    .ZN(_15234_)
  );
  AND2_X1 _50360_ (
    .A1(\cpuregs[19] [23]),
    .A2(_12792_),
    .ZN(_15235_)
  );
  INV_X1 _50361_ (
    .A(_15235_),
    .ZN(_15236_)
  );
  AND2_X1 _50362_ (
    .A1(_15234_),
    .A2(_15236_),
    .ZN(_15237_)
  );
  INV_X1 _50363_ (
    .A(_15237_),
    .ZN(_00953_)
  );
  AND2_X1 _50364_ (
    .A1(_12791_),
    .A2(_13229_),
    .ZN(_15238_)
  );
  INV_X1 _50365_ (
    .A(_15238_),
    .ZN(_15239_)
  );
  AND2_X1 _50366_ (
    .A1(\cpuregs[19] [24]),
    .A2(_12792_),
    .ZN(_15240_)
  );
  INV_X1 _50367_ (
    .A(_15240_),
    .ZN(_15241_)
  );
  AND2_X1 _50368_ (
    .A1(_15239_),
    .A2(_15241_),
    .ZN(_15242_)
  );
  INV_X1 _50369_ (
    .A(_15242_),
    .ZN(_00954_)
  );
  AND2_X1 _50370_ (
    .A1(_12791_),
    .A2(_13244_),
    .ZN(_15243_)
  );
  INV_X1 _50371_ (
    .A(_15243_),
    .ZN(_15244_)
  );
  AND2_X1 _50372_ (
    .A1(\cpuregs[19] [25]),
    .A2(_12792_),
    .ZN(_15245_)
  );
  INV_X1 _50373_ (
    .A(_15245_),
    .ZN(_15246_)
  );
  AND2_X1 _50374_ (
    .A1(_15244_),
    .A2(_15246_),
    .ZN(_15247_)
  );
  INV_X1 _50375_ (
    .A(_15247_),
    .ZN(_00955_)
  );
  AND2_X1 _50376_ (
    .A1(_12791_),
    .A2(_13259_),
    .ZN(_15248_)
  );
  INV_X1 _50377_ (
    .A(_15248_),
    .ZN(_15249_)
  );
  AND2_X1 _50378_ (
    .A1(\cpuregs[19] [26]),
    .A2(_12792_),
    .ZN(_15250_)
  );
  INV_X1 _50379_ (
    .A(_15250_),
    .ZN(_15251_)
  );
  AND2_X1 _50380_ (
    .A1(_15249_),
    .A2(_15251_),
    .ZN(_15252_)
  );
  INV_X1 _50381_ (
    .A(_15252_),
    .ZN(_00956_)
  );
  AND2_X1 _50382_ (
    .A1(_12791_),
    .A2(_13274_),
    .ZN(_15253_)
  );
  INV_X1 _50383_ (
    .A(_15253_),
    .ZN(_15254_)
  );
  AND2_X1 _50384_ (
    .A1(\cpuregs[19] [27]),
    .A2(_12792_),
    .ZN(_15255_)
  );
  INV_X1 _50385_ (
    .A(_15255_),
    .ZN(_15256_)
  );
  AND2_X1 _50386_ (
    .A1(_15254_),
    .A2(_15256_),
    .ZN(_15257_)
  );
  INV_X1 _50387_ (
    .A(_15257_),
    .ZN(_00957_)
  );
  AND2_X1 _50388_ (
    .A1(_12791_),
    .A2(_13289_),
    .ZN(_15258_)
  );
  INV_X1 _50389_ (
    .A(_15258_),
    .ZN(_15259_)
  );
  AND2_X1 _50390_ (
    .A1(\cpuregs[19] [28]),
    .A2(_12792_),
    .ZN(_15260_)
  );
  INV_X1 _50391_ (
    .A(_15260_),
    .ZN(_15261_)
  );
  AND2_X1 _50392_ (
    .A1(_15259_),
    .A2(_15261_),
    .ZN(_15262_)
  );
  INV_X1 _50393_ (
    .A(_15262_),
    .ZN(_00958_)
  );
  AND2_X1 _50394_ (
    .A1(_12791_),
    .A2(_13304_),
    .ZN(_15263_)
  );
  INV_X1 _50395_ (
    .A(_15263_),
    .ZN(_15264_)
  );
  AND2_X1 _50396_ (
    .A1(\cpuregs[19] [29]),
    .A2(_12792_),
    .ZN(_15265_)
  );
  INV_X1 _50397_ (
    .A(_15265_),
    .ZN(_15266_)
  );
  AND2_X1 _50398_ (
    .A1(_15264_),
    .A2(_15266_),
    .ZN(_15267_)
  );
  INV_X1 _50399_ (
    .A(_15267_),
    .ZN(_00959_)
  );
  AND2_X1 _50400_ (
    .A1(_12791_),
    .A2(_13319_),
    .ZN(_15268_)
  );
  INV_X1 _50401_ (
    .A(_15268_),
    .ZN(_15269_)
  );
  AND2_X1 _50402_ (
    .A1(\cpuregs[19] [30]),
    .A2(_12792_),
    .ZN(_15270_)
  );
  INV_X1 _50403_ (
    .A(_15270_),
    .ZN(_15271_)
  );
  AND2_X1 _50404_ (
    .A1(_15269_),
    .A2(_15271_),
    .ZN(_15272_)
  );
  INV_X1 _50405_ (
    .A(_15272_),
    .ZN(_00960_)
  );
  AND2_X1 _50406_ (
    .A1(_12835_),
    .A2(_12874_),
    .ZN(_15273_)
  );
  INV_X1 _50407_ (
    .A(_15273_),
    .ZN(_15274_)
  );
  AND2_X1 _50408_ (
    .A1(\cpuregs[13] [0]),
    .A2(_12836_),
    .ZN(_15275_)
  );
  INV_X1 _50409_ (
    .A(_15275_),
    .ZN(_15276_)
  );
  AND2_X1 _50410_ (
    .A1(_15274_),
    .A2(_15276_),
    .ZN(_15277_)
  );
  INV_X1 _50411_ (
    .A(_15277_),
    .ZN(_00961_)
  );
  AND2_X1 _50412_ (
    .A1(_12835_),
    .A2(_12886_),
    .ZN(_15278_)
  );
  INV_X1 _50413_ (
    .A(_15278_),
    .ZN(_15279_)
  );
  AND2_X1 _50414_ (
    .A1(\cpuregs[13] [1]),
    .A2(_12836_),
    .ZN(_15280_)
  );
  INV_X1 _50415_ (
    .A(_15280_),
    .ZN(_15281_)
  );
  AND2_X1 _50416_ (
    .A1(_15279_),
    .A2(_15281_),
    .ZN(_15282_)
  );
  INV_X1 _50417_ (
    .A(_15282_),
    .ZN(_00962_)
  );
  AND2_X1 _50418_ (
    .A1(\cpuregs[13] [2]),
    .A2(_12836_),
    .ZN(_15283_)
  );
  INV_X1 _50419_ (
    .A(_15283_),
    .ZN(_15284_)
  );
  AND2_X1 _50420_ (
    .A1(_12835_),
    .A2(_12900_),
    .ZN(_15285_)
  );
  INV_X1 _50421_ (
    .A(_15285_),
    .ZN(_15286_)
  );
  AND2_X1 _50422_ (
    .A1(_15284_),
    .A2(_15286_),
    .ZN(_15287_)
  );
  INV_X1 _50423_ (
    .A(_15287_),
    .ZN(_00963_)
  );
  AND2_X1 _50424_ (
    .A1(_12835_),
    .A2(_12913_),
    .ZN(_15288_)
  );
  INV_X1 _50425_ (
    .A(_15288_),
    .ZN(_15289_)
  );
  AND2_X1 _50426_ (
    .A1(\cpuregs[13] [3]),
    .A2(_12836_),
    .ZN(_15290_)
  );
  INV_X1 _50427_ (
    .A(_15290_),
    .ZN(_15291_)
  );
  AND2_X1 _50428_ (
    .A1(_15289_),
    .A2(_15291_),
    .ZN(_15292_)
  );
  INV_X1 _50429_ (
    .A(_15292_),
    .ZN(_00964_)
  );
  AND2_X1 _50430_ (
    .A1(\cpuregs[13] [4]),
    .A2(_12836_),
    .ZN(_15293_)
  );
  INV_X1 _50431_ (
    .A(_15293_),
    .ZN(_15294_)
  );
  AND2_X1 _50432_ (
    .A1(_12835_),
    .A2(_12928_),
    .ZN(_15295_)
  );
  INV_X1 _50433_ (
    .A(_15295_),
    .ZN(_15296_)
  );
  AND2_X1 _50434_ (
    .A1(_15294_),
    .A2(_15296_),
    .ZN(_15297_)
  );
  INV_X1 _50435_ (
    .A(_15297_),
    .ZN(_00965_)
  );
  AND2_X1 _50436_ (
    .A1(_12835_),
    .A2(_12943_),
    .ZN(_15298_)
  );
  INV_X1 _50437_ (
    .A(_15298_),
    .ZN(_15299_)
  );
  AND2_X1 _50438_ (
    .A1(\cpuregs[13] [5]),
    .A2(_12836_),
    .ZN(_15300_)
  );
  INV_X1 _50439_ (
    .A(_15300_),
    .ZN(_15301_)
  );
  AND2_X1 _50440_ (
    .A1(_15299_),
    .A2(_15301_),
    .ZN(_15302_)
  );
  INV_X1 _50441_ (
    .A(_15302_),
    .ZN(_00966_)
  );
  AND2_X1 _50442_ (
    .A1(_12835_),
    .A2(_12958_),
    .ZN(_15303_)
  );
  INV_X1 _50443_ (
    .A(_15303_),
    .ZN(_15304_)
  );
  AND2_X1 _50444_ (
    .A1(\cpuregs[13] [6]),
    .A2(_12836_),
    .ZN(_15305_)
  );
  INV_X1 _50445_ (
    .A(_15305_),
    .ZN(_15306_)
  );
  AND2_X1 _50446_ (
    .A1(_15304_),
    .A2(_15306_),
    .ZN(_15307_)
  );
  INV_X1 _50447_ (
    .A(_15307_),
    .ZN(_00967_)
  );
  AND2_X1 _50448_ (
    .A1(_12835_),
    .A2(_12973_),
    .ZN(_15308_)
  );
  INV_X1 _50449_ (
    .A(_15308_),
    .ZN(_15309_)
  );
  AND2_X1 _50450_ (
    .A1(\cpuregs[13] [7]),
    .A2(_12836_),
    .ZN(_15310_)
  );
  INV_X1 _50451_ (
    .A(_15310_),
    .ZN(_15311_)
  );
  AND2_X1 _50452_ (
    .A1(_15309_),
    .A2(_15311_),
    .ZN(_15312_)
  );
  INV_X1 _50453_ (
    .A(_15312_),
    .ZN(_00968_)
  );
  AND2_X1 _50454_ (
    .A1(_12835_),
    .A2(_12988_),
    .ZN(_15313_)
  );
  INV_X1 _50455_ (
    .A(_15313_),
    .ZN(_15314_)
  );
  AND2_X1 _50456_ (
    .A1(\cpuregs[13] [8]),
    .A2(_12836_),
    .ZN(_15315_)
  );
  INV_X1 _50457_ (
    .A(_15315_),
    .ZN(_15316_)
  );
  AND2_X1 _50458_ (
    .A1(_15314_),
    .A2(_15316_),
    .ZN(_15317_)
  );
  INV_X1 _50459_ (
    .A(_15317_),
    .ZN(_00969_)
  );
  AND2_X1 _50460_ (
    .A1(_12835_),
    .A2(_13003_),
    .ZN(_15318_)
  );
  INV_X1 _50461_ (
    .A(_15318_),
    .ZN(_15319_)
  );
  AND2_X1 _50462_ (
    .A1(\cpuregs[13] [9]),
    .A2(_12836_),
    .ZN(_15320_)
  );
  INV_X1 _50463_ (
    .A(_15320_),
    .ZN(_15321_)
  );
  AND2_X1 _50464_ (
    .A1(_15319_),
    .A2(_15321_),
    .ZN(_15322_)
  );
  INV_X1 _50465_ (
    .A(_15322_),
    .ZN(_00970_)
  );
  AND2_X1 _50466_ (
    .A1(_12835_),
    .A2(_13018_),
    .ZN(_15323_)
  );
  INV_X1 _50467_ (
    .A(_15323_),
    .ZN(_15324_)
  );
  AND2_X1 _50468_ (
    .A1(\cpuregs[13] [10]),
    .A2(_12836_),
    .ZN(_15325_)
  );
  INV_X1 _50469_ (
    .A(_15325_),
    .ZN(_15326_)
  );
  AND2_X1 _50470_ (
    .A1(_15324_),
    .A2(_15326_),
    .ZN(_15327_)
  );
  INV_X1 _50471_ (
    .A(_15327_),
    .ZN(_00971_)
  );
  AND2_X1 _50472_ (
    .A1(_12835_),
    .A2(_13033_),
    .ZN(_15328_)
  );
  INV_X1 _50473_ (
    .A(_15328_),
    .ZN(_15329_)
  );
  AND2_X1 _50474_ (
    .A1(\cpuregs[13] [11]),
    .A2(_12836_),
    .ZN(_15330_)
  );
  INV_X1 _50475_ (
    .A(_15330_),
    .ZN(_15331_)
  );
  AND2_X1 _50476_ (
    .A1(_15329_),
    .A2(_15331_),
    .ZN(_15332_)
  );
  INV_X1 _50477_ (
    .A(_15332_),
    .ZN(_00972_)
  );
  AND2_X1 _50478_ (
    .A1(_12835_),
    .A2(_13048_),
    .ZN(_15333_)
  );
  INV_X1 _50479_ (
    .A(_15333_),
    .ZN(_15334_)
  );
  AND2_X1 _50480_ (
    .A1(\cpuregs[13] [12]),
    .A2(_12836_),
    .ZN(_15335_)
  );
  INV_X1 _50481_ (
    .A(_15335_),
    .ZN(_15336_)
  );
  AND2_X1 _50482_ (
    .A1(_15334_),
    .A2(_15336_),
    .ZN(_15337_)
  );
  INV_X1 _50483_ (
    .A(_15337_),
    .ZN(_00973_)
  );
  AND2_X1 _50484_ (
    .A1(_12835_),
    .A2(_13063_),
    .ZN(_15338_)
  );
  INV_X1 _50485_ (
    .A(_15338_),
    .ZN(_15339_)
  );
  AND2_X1 _50486_ (
    .A1(\cpuregs[13] [13]),
    .A2(_12836_),
    .ZN(_15340_)
  );
  INV_X1 _50487_ (
    .A(_15340_),
    .ZN(_15341_)
  );
  AND2_X1 _50488_ (
    .A1(_15339_),
    .A2(_15341_),
    .ZN(_15342_)
  );
  INV_X1 _50489_ (
    .A(_15342_),
    .ZN(_00974_)
  );
  AND2_X1 _50490_ (
    .A1(_12835_),
    .A2(_13078_),
    .ZN(_15343_)
  );
  INV_X1 _50491_ (
    .A(_15343_),
    .ZN(_15344_)
  );
  AND2_X1 _50492_ (
    .A1(\cpuregs[13] [14]),
    .A2(_12836_),
    .ZN(_15345_)
  );
  INV_X1 _50493_ (
    .A(_15345_),
    .ZN(_15346_)
  );
  AND2_X1 _50494_ (
    .A1(_15344_),
    .A2(_15346_),
    .ZN(_15347_)
  );
  INV_X1 _50495_ (
    .A(_15347_),
    .ZN(_00975_)
  );
  AND2_X1 _50496_ (
    .A1(_12835_),
    .A2(_13093_),
    .ZN(_15348_)
  );
  INV_X1 _50497_ (
    .A(_15348_),
    .ZN(_15349_)
  );
  AND2_X1 _50498_ (
    .A1(\cpuregs[13] [15]),
    .A2(_12836_),
    .ZN(_15350_)
  );
  INV_X1 _50499_ (
    .A(_15350_),
    .ZN(_15351_)
  );
  AND2_X1 _50500_ (
    .A1(_15349_),
    .A2(_15351_),
    .ZN(_15352_)
  );
  INV_X1 _50501_ (
    .A(_15352_),
    .ZN(_00976_)
  );
  AND2_X1 _50502_ (
    .A1(_12835_),
    .A2(_13108_),
    .ZN(_15353_)
  );
  INV_X1 _50503_ (
    .A(_15353_),
    .ZN(_15354_)
  );
  AND2_X1 _50504_ (
    .A1(\cpuregs[13] [16]),
    .A2(_12836_),
    .ZN(_15355_)
  );
  INV_X1 _50505_ (
    .A(_15355_),
    .ZN(_15356_)
  );
  AND2_X1 _50506_ (
    .A1(_15354_),
    .A2(_15356_),
    .ZN(_15357_)
  );
  INV_X1 _50507_ (
    .A(_15357_),
    .ZN(_00977_)
  );
  AND2_X1 _50508_ (
    .A1(_21643_),
    .A2(_12836_),
    .ZN(_15358_)
  );
  INV_X1 _50509_ (
    .A(_15358_),
    .ZN(_15359_)
  );
  AND2_X1 _50510_ (
    .A1(_12835_),
    .A2(_13124_),
    .ZN(_15360_)
  );
  INV_X1 _50511_ (
    .A(_15360_),
    .ZN(_15361_)
  );
  AND2_X1 _50512_ (
    .A1(_15359_),
    .A2(_15361_),
    .ZN(_00978_)
  );
  AND2_X1 _50513_ (
    .A1(\cpuregs[13] [18]),
    .A2(_12836_),
    .ZN(_15362_)
  );
  INV_X1 _50514_ (
    .A(_15362_),
    .ZN(_15363_)
  );
  AND2_X1 _50515_ (
    .A1(_12835_),
    .A2(_13139_),
    .ZN(_15364_)
  );
  INV_X1 _50516_ (
    .A(_15364_),
    .ZN(_15365_)
  );
  AND2_X1 _50517_ (
    .A1(_15363_),
    .A2(_15365_),
    .ZN(_15366_)
  );
  INV_X1 _50518_ (
    .A(_15366_),
    .ZN(_00979_)
  );
  AND2_X1 _50519_ (
    .A1(\cpuregs[13] [19]),
    .A2(_12836_),
    .ZN(_15367_)
  );
  INV_X1 _50520_ (
    .A(_15367_),
    .ZN(_15368_)
  );
  AND2_X1 _50521_ (
    .A1(_12835_),
    .A2(_13154_),
    .ZN(_15369_)
  );
  INV_X1 _50522_ (
    .A(_15369_),
    .ZN(_15370_)
  );
  AND2_X1 _50523_ (
    .A1(_15368_),
    .A2(_15370_),
    .ZN(_15371_)
  );
  INV_X1 _50524_ (
    .A(_15371_),
    .ZN(_00980_)
  );
  AND2_X1 _50525_ (
    .A1(\cpuregs[13] [20]),
    .A2(_12836_),
    .ZN(_15372_)
  );
  INV_X1 _50526_ (
    .A(_15372_),
    .ZN(_15373_)
  );
  AND2_X1 _50527_ (
    .A1(_12835_),
    .A2(_13169_),
    .ZN(_15374_)
  );
  INV_X1 _50528_ (
    .A(_15374_),
    .ZN(_15375_)
  );
  AND2_X1 _50529_ (
    .A1(_15373_),
    .A2(_15375_),
    .ZN(_15376_)
  );
  INV_X1 _50530_ (
    .A(_15376_),
    .ZN(_00981_)
  );
  AND2_X1 _50531_ (
    .A1(\cpuregs[13] [21]),
    .A2(_12836_),
    .ZN(_15377_)
  );
  INV_X1 _50532_ (
    .A(_15377_),
    .ZN(_15378_)
  );
  AND2_X1 _50533_ (
    .A1(_12835_),
    .A2(_13184_),
    .ZN(_15379_)
  );
  INV_X1 _50534_ (
    .A(_15379_),
    .ZN(_15380_)
  );
  AND2_X1 _50535_ (
    .A1(_15378_),
    .A2(_15380_),
    .ZN(_15381_)
  );
  INV_X1 _50536_ (
    .A(_15381_),
    .ZN(_00982_)
  );
  AND2_X1 _50537_ (
    .A1(\cpuregs[13] [22]),
    .A2(_12836_),
    .ZN(_15382_)
  );
  INV_X1 _50538_ (
    .A(_15382_),
    .ZN(_15383_)
  );
  AND2_X1 _50539_ (
    .A1(_12835_),
    .A2(_13199_),
    .ZN(_15384_)
  );
  INV_X1 _50540_ (
    .A(_15384_),
    .ZN(_15385_)
  );
  AND2_X1 _50541_ (
    .A1(_15383_),
    .A2(_15385_),
    .ZN(_15386_)
  );
  INV_X1 _50542_ (
    .A(_15386_),
    .ZN(_00983_)
  );
  AND2_X1 _50543_ (
    .A1(\cpuregs[13] [23]),
    .A2(_12836_),
    .ZN(_15387_)
  );
  INV_X1 _50544_ (
    .A(_15387_),
    .ZN(_15388_)
  );
  AND2_X1 _50545_ (
    .A1(_12835_),
    .A2(_13214_),
    .ZN(_15389_)
  );
  INV_X1 _50546_ (
    .A(_15389_),
    .ZN(_15390_)
  );
  AND2_X1 _50547_ (
    .A1(_15388_),
    .A2(_15390_),
    .ZN(_15391_)
  );
  INV_X1 _50548_ (
    .A(_15391_),
    .ZN(_00984_)
  );
  AND2_X1 _50549_ (
    .A1(\cpuregs[13] [24]),
    .A2(_12836_),
    .ZN(_15392_)
  );
  INV_X1 _50550_ (
    .A(_15392_),
    .ZN(_15393_)
  );
  AND2_X1 _50551_ (
    .A1(_12835_),
    .A2(_13229_),
    .ZN(_15394_)
  );
  INV_X1 _50552_ (
    .A(_15394_),
    .ZN(_15395_)
  );
  AND2_X1 _50553_ (
    .A1(_15393_),
    .A2(_15395_),
    .ZN(_15396_)
  );
  INV_X1 _50554_ (
    .A(_15396_),
    .ZN(_00985_)
  );
  AND2_X1 _50555_ (
    .A1(\cpuregs[13] [25]),
    .A2(_12836_),
    .ZN(_15397_)
  );
  INV_X1 _50556_ (
    .A(_15397_),
    .ZN(_15398_)
  );
  AND2_X1 _50557_ (
    .A1(_12835_),
    .A2(_13244_),
    .ZN(_15399_)
  );
  INV_X1 _50558_ (
    .A(_15399_),
    .ZN(_15400_)
  );
  AND2_X1 _50559_ (
    .A1(_15398_),
    .A2(_15400_),
    .ZN(_15401_)
  );
  INV_X1 _50560_ (
    .A(_15401_),
    .ZN(_00986_)
  );
  AND2_X1 _50561_ (
    .A1(\cpuregs[13] [26]),
    .A2(_12836_),
    .ZN(_15402_)
  );
  INV_X1 _50562_ (
    .A(_15402_),
    .ZN(_15403_)
  );
  AND2_X1 _50563_ (
    .A1(_12835_),
    .A2(_13259_),
    .ZN(_15404_)
  );
  INV_X1 _50564_ (
    .A(_15404_),
    .ZN(_15405_)
  );
  AND2_X1 _50565_ (
    .A1(_15403_),
    .A2(_15405_),
    .ZN(_15406_)
  );
  INV_X1 _50566_ (
    .A(_15406_),
    .ZN(_00987_)
  );
  AND2_X1 _50567_ (
    .A1(\cpuregs[13] [27]),
    .A2(_12836_),
    .ZN(_15407_)
  );
  INV_X1 _50568_ (
    .A(_15407_),
    .ZN(_15408_)
  );
  AND2_X1 _50569_ (
    .A1(_12835_),
    .A2(_13274_),
    .ZN(_15409_)
  );
  INV_X1 _50570_ (
    .A(_15409_),
    .ZN(_15410_)
  );
  AND2_X1 _50571_ (
    .A1(_15408_),
    .A2(_15410_),
    .ZN(_15411_)
  );
  INV_X1 _50572_ (
    .A(_15411_),
    .ZN(_00988_)
  );
  AND2_X1 _50573_ (
    .A1(\cpuregs[13] [28]),
    .A2(_12836_),
    .ZN(_15412_)
  );
  INV_X1 _50574_ (
    .A(_15412_),
    .ZN(_15413_)
  );
  AND2_X1 _50575_ (
    .A1(_12835_),
    .A2(_13289_),
    .ZN(_15414_)
  );
  INV_X1 _50576_ (
    .A(_15414_),
    .ZN(_15415_)
  );
  AND2_X1 _50577_ (
    .A1(_15413_),
    .A2(_15415_),
    .ZN(_15416_)
  );
  INV_X1 _50578_ (
    .A(_15416_),
    .ZN(_00989_)
  );
  AND2_X1 _50579_ (
    .A1(\cpuregs[13] [29]),
    .A2(_12836_),
    .ZN(_15417_)
  );
  INV_X1 _50580_ (
    .A(_15417_),
    .ZN(_15418_)
  );
  AND2_X1 _50581_ (
    .A1(_12835_),
    .A2(_13304_),
    .ZN(_15419_)
  );
  INV_X1 _50582_ (
    .A(_15419_),
    .ZN(_15420_)
  );
  AND2_X1 _50583_ (
    .A1(_15418_),
    .A2(_15420_),
    .ZN(_15421_)
  );
  INV_X1 _50584_ (
    .A(_15421_),
    .ZN(_00990_)
  );
  AND2_X1 _50585_ (
    .A1(\cpuregs[13] [30]),
    .A2(_12836_),
    .ZN(_15422_)
  );
  INV_X1 _50586_ (
    .A(_15422_),
    .ZN(_15423_)
  );
  AND2_X1 _50587_ (
    .A1(_12835_),
    .A2(_13319_),
    .ZN(_15424_)
  );
  INV_X1 _50588_ (
    .A(_15424_),
    .ZN(_15425_)
  );
  AND2_X1 _50589_ (
    .A1(_15423_),
    .A2(_15425_),
    .ZN(_15426_)
  );
  INV_X1 _50590_ (
    .A(_15426_),
    .ZN(_00991_)
  );
  AND2_X1 _50591_ (
    .A1(_12776_),
    .A2(_12874_),
    .ZN(_15427_)
  );
  INV_X1 _50592_ (
    .A(_15427_),
    .ZN(_15428_)
  );
  AND2_X1 _50593_ (
    .A1(\cpuregs[20] [0]),
    .A2(_12777_),
    .ZN(_15429_)
  );
  INV_X1 _50594_ (
    .A(_15429_),
    .ZN(_15430_)
  );
  AND2_X1 _50595_ (
    .A1(_15428_),
    .A2(_15430_),
    .ZN(_15431_)
  );
  INV_X1 _50596_ (
    .A(_15431_),
    .ZN(_00992_)
  );
  AND2_X1 _50597_ (
    .A1(_12776_),
    .A2(_12886_),
    .ZN(_15432_)
  );
  INV_X1 _50598_ (
    .A(_15432_),
    .ZN(_15433_)
  );
  AND2_X1 _50599_ (
    .A1(\cpuregs[20] [1]),
    .A2(_12777_),
    .ZN(_15434_)
  );
  INV_X1 _50600_ (
    .A(_15434_),
    .ZN(_15435_)
  );
  AND2_X1 _50601_ (
    .A1(_15433_),
    .A2(_15435_),
    .ZN(_15436_)
  );
  INV_X1 _50602_ (
    .A(_15436_),
    .ZN(_00993_)
  );
  AND2_X1 _50603_ (
    .A1(_12776_),
    .A2(_12900_),
    .ZN(_15437_)
  );
  INV_X1 _50604_ (
    .A(_15437_),
    .ZN(_15438_)
  );
  AND2_X1 _50605_ (
    .A1(\cpuregs[20] [2]),
    .A2(_12777_),
    .ZN(_15439_)
  );
  INV_X1 _50606_ (
    .A(_15439_),
    .ZN(_15440_)
  );
  AND2_X1 _50607_ (
    .A1(_15438_),
    .A2(_15440_),
    .ZN(_15441_)
  );
  INV_X1 _50608_ (
    .A(_15441_),
    .ZN(_00994_)
  );
  AND2_X1 _50609_ (
    .A1(_12776_),
    .A2(_12913_),
    .ZN(_15442_)
  );
  INV_X1 _50610_ (
    .A(_15442_),
    .ZN(_15443_)
  );
  AND2_X1 _50611_ (
    .A1(\cpuregs[20] [3]),
    .A2(_12777_),
    .ZN(_15444_)
  );
  INV_X1 _50612_ (
    .A(_15444_),
    .ZN(_15445_)
  );
  AND2_X1 _50613_ (
    .A1(_15443_),
    .A2(_15445_),
    .ZN(_15446_)
  );
  INV_X1 _50614_ (
    .A(_15446_),
    .ZN(_00995_)
  );
  AND2_X1 _50615_ (
    .A1(_12776_),
    .A2(_12928_),
    .ZN(_15447_)
  );
  INV_X1 _50616_ (
    .A(_15447_),
    .ZN(_15448_)
  );
  AND2_X1 _50617_ (
    .A1(\cpuregs[20] [4]),
    .A2(_12777_),
    .ZN(_15449_)
  );
  INV_X1 _50618_ (
    .A(_15449_),
    .ZN(_15450_)
  );
  AND2_X1 _50619_ (
    .A1(_15448_),
    .A2(_15450_),
    .ZN(_15451_)
  );
  INV_X1 _50620_ (
    .A(_15451_),
    .ZN(_00996_)
  );
  AND2_X1 _50621_ (
    .A1(_12776_),
    .A2(_12943_),
    .ZN(_15452_)
  );
  INV_X1 _50622_ (
    .A(_15452_),
    .ZN(_15453_)
  );
  AND2_X1 _50623_ (
    .A1(\cpuregs[20] [5]),
    .A2(_12777_),
    .ZN(_15454_)
  );
  INV_X1 _50624_ (
    .A(_15454_),
    .ZN(_15455_)
  );
  AND2_X1 _50625_ (
    .A1(_15453_),
    .A2(_15455_),
    .ZN(_15456_)
  );
  INV_X1 _50626_ (
    .A(_15456_),
    .ZN(_00997_)
  );
  AND2_X1 _50627_ (
    .A1(_12776_),
    .A2(_12958_),
    .ZN(_15457_)
  );
  INV_X1 _50628_ (
    .A(_15457_),
    .ZN(_15458_)
  );
  AND2_X1 _50629_ (
    .A1(\cpuregs[20] [6]),
    .A2(_12777_),
    .ZN(_15459_)
  );
  INV_X1 _50630_ (
    .A(_15459_),
    .ZN(_15460_)
  );
  AND2_X1 _50631_ (
    .A1(_15458_),
    .A2(_15460_),
    .ZN(_15461_)
  );
  INV_X1 _50632_ (
    .A(_15461_),
    .ZN(_00998_)
  );
  AND2_X1 _50633_ (
    .A1(_12776_),
    .A2(_12973_),
    .ZN(_15462_)
  );
  INV_X1 _50634_ (
    .A(_15462_),
    .ZN(_15463_)
  );
  AND2_X1 _50635_ (
    .A1(\cpuregs[20] [7]),
    .A2(_12777_),
    .ZN(_15464_)
  );
  INV_X1 _50636_ (
    .A(_15464_),
    .ZN(_15465_)
  );
  AND2_X1 _50637_ (
    .A1(_15463_),
    .A2(_15465_),
    .ZN(_15466_)
  );
  INV_X1 _50638_ (
    .A(_15466_),
    .ZN(_00999_)
  );
  AND2_X1 _50639_ (
    .A1(_12776_),
    .A2(_12988_),
    .ZN(_15467_)
  );
  INV_X1 _50640_ (
    .A(_15467_),
    .ZN(_15468_)
  );
  AND2_X1 _50641_ (
    .A1(\cpuregs[20] [8]),
    .A2(_12777_),
    .ZN(_15469_)
  );
  INV_X1 _50642_ (
    .A(_15469_),
    .ZN(_15470_)
  );
  AND2_X1 _50643_ (
    .A1(_15468_),
    .A2(_15470_),
    .ZN(_15471_)
  );
  INV_X1 _50644_ (
    .A(_15471_),
    .ZN(_01000_)
  );
  AND2_X1 _50645_ (
    .A1(_12776_),
    .A2(_13003_),
    .ZN(_15472_)
  );
  INV_X1 _50646_ (
    .A(_15472_),
    .ZN(_15473_)
  );
  AND2_X1 _50647_ (
    .A1(\cpuregs[20] [9]),
    .A2(_12777_),
    .ZN(_15474_)
  );
  INV_X1 _50648_ (
    .A(_15474_),
    .ZN(_15475_)
  );
  AND2_X1 _50649_ (
    .A1(_15473_),
    .A2(_15475_),
    .ZN(_15476_)
  );
  INV_X1 _50650_ (
    .A(_15476_),
    .ZN(_01001_)
  );
  AND2_X1 _50651_ (
    .A1(_12776_),
    .A2(_13018_),
    .ZN(_15477_)
  );
  INV_X1 _50652_ (
    .A(_15477_),
    .ZN(_15478_)
  );
  AND2_X1 _50653_ (
    .A1(\cpuregs[20] [10]),
    .A2(_12777_),
    .ZN(_15479_)
  );
  INV_X1 _50654_ (
    .A(_15479_),
    .ZN(_15480_)
  );
  AND2_X1 _50655_ (
    .A1(_15478_),
    .A2(_15480_),
    .ZN(_15481_)
  );
  INV_X1 _50656_ (
    .A(_15481_),
    .ZN(_01002_)
  );
  AND2_X1 _50657_ (
    .A1(_12776_),
    .A2(_13033_),
    .ZN(_15482_)
  );
  INV_X1 _50658_ (
    .A(_15482_),
    .ZN(_15483_)
  );
  AND2_X1 _50659_ (
    .A1(\cpuregs[20] [11]),
    .A2(_12777_),
    .ZN(_15484_)
  );
  INV_X1 _50660_ (
    .A(_15484_),
    .ZN(_15485_)
  );
  AND2_X1 _50661_ (
    .A1(_15483_),
    .A2(_15485_),
    .ZN(_15486_)
  );
  INV_X1 _50662_ (
    .A(_15486_),
    .ZN(_01003_)
  );
  AND2_X1 _50663_ (
    .A1(_12776_),
    .A2(_13048_),
    .ZN(_15487_)
  );
  INV_X1 _50664_ (
    .A(_15487_),
    .ZN(_15488_)
  );
  AND2_X1 _50665_ (
    .A1(\cpuregs[20] [12]),
    .A2(_12777_),
    .ZN(_15489_)
  );
  INV_X1 _50666_ (
    .A(_15489_),
    .ZN(_15490_)
  );
  AND2_X1 _50667_ (
    .A1(_15488_),
    .A2(_15490_),
    .ZN(_15491_)
  );
  INV_X1 _50668_ (
    .A(_15491_),
    .ZN(_01004_)
  );
  AND2_X1 _50669_ (
    .A1(_12776_),
    .A2(_13063_),
    .ZN(_15492_)
  );
  INV_X1 _50670_ (
    .A(_15492_),
    .ZN(_15493_)
  );
  AND2_X1 _50671_ (
    .A1(\cpuregs[20] [13]),
    .A2(_12777_),
    .ZN(_15494_)
  );
  INV_X1 _50672_ (
    .A(_15494_),
    .ZN(_15495_)
  );
  AND2_X1 _50673_ (
    .A1(_15493_),
    .A2(_15495_),
    .ZN(_15496_)
  );
  INV_X1 _50674_ (
    .A(_15496_),
    .ZN(_01005_)
  );
  AND2_X1 _50675_ (
    .A1(\cpuregs[20] [14]),
    .A2(_12777_),
    .ZN(_15497_)
  );
  INV_X1 _50676_ (
    .A(_15497_),
    .ZN(_15498_)
  );
  AND2_X1 _50677_ (
    .A1(_12776_),
    .A2(_13078_),
    .ZN(_15499_)
  );
  INV_X1 _50678_ (
    .A(_15499_),
    .ZN(_15500_)
  );
  AND2_X1 _50679_ (
    .A1(_15498_),
    .A2(_15500_),
    .ZN(_15501_)
  );
  INV_X1 _50680_ (
    .A(_15501_),
    .ZN(_01006_)
  );
  AND2_X1 _50681_ (
    .A1(_12776_),
    .A2(_13093_),
    .ZN(_15502_)
  );
  INV_X1 _50682_ (
    .A(_15502_),
    .ZN(_15503_)
  );
  AND2_X1 _50683_ (
    .A1(\cpuregs[20] [15]),
    .A2(_12777_),
    .ZN(_15504_)
  );
  INV_X1 _50684_ (
    .A(_15504_),
    .ZN(_15505_)
  );
  AND2_X1 _50685_ (
    .A1(_15503_),
    .A2(_15505_),
    .ZN(_15506_)
  );
  INV_X1 _50686_ (
    .A(_15506_),
    .ZN(_01007_)
  );
  AND2_X1 _50687_ (
    .A1(\cpuregs[20] [16]),
    .A2(_12777_),
    .ZN(_15507_)
  );
  INV_X1 _50688_ (
    .A(_15507_),
    .ZN(_15508_)
  );
  AND2_X1 _50689_ (
    .A1(_12776_),
    .A2(_13108_),
    .ZN(_15509_)
  );
  INV_X1 _50690_ (
    .A(_15509_),
    .ZN(_15510_)
  );
  AND2_X1 _50691_ (
    .A1(_15508_),
    .A2(_15510_),
    .ZN(_15511_)
  );
  INV_X1 _50692_ (
    .A(_15511_),
    .ZN(_01008_)
  );
  AND2_X1 _50693_ (
    .A1(_12776_),
    .A2(_13123_),
    .ZN(_15512_)
  );
  INV_X1 _50694_ (
    .A(_15512_),
    .ZN(_15513_)
  );
  AND2_X1 _50695_ (
    .A1(\cpuregs[20] [17]),
    .A2(_12777_),
    .ZN(_15514_)
  );
  INV_X1 _50696_ (
    .A(_15514_),
    .ZN(_15515_)
  );
  AND2_X1 _50697_ (
    .A1(_15513_),
    .A2(_15515_),
    .ZN(_15516_)
  );
  INV_X1 _50698_ (
    .A(_15516_),
    .ZN(_01009_)
  );
  AND2_X1 _50699_ (
    .A1(_12776_),
    .A2(_13139_),
    .ZN(_15517_)
  );
  INV_X1 _50700_ (
    .A(_15517_),
    .ZN(_15518_)
  );
  AND2_X1 _50701_ (
    .A1(\cpuregs[20] [18]),
    .A2(_12777_),
    .ZN(_15519_)
  );
  INV_X1 _50702_ (
    .A(_15519_),
    .ZN(_15520_)
  );
  AND2_X1 _50703_ (
    .A1(_15518_),
    .A2(_15520_),
    .ZN(_15521_)
  );
  INV_X1 _50704_ (
    .A(_15521_),
    .ZN(_01010_)
  );
  AND2_X1 _50705_ (
    .A1(_12776_),
    .A2(_13154_),
    .ZN(_15522_)
  );
  INV_X1 _50706_ (
    .A(_15522_),
    .ZN(_15523_)
  );
  AND2_X1 _50707_ (
    .A1(\cpuregs[20] [19]),
    .A2(_12777_),
    .ZN(_15524_)
  );
  INV_X1 _50708_ (
    .A(_15524_),
    .ZN(_15525_)
  );
  AND2_X1 _50709_ (
    .A1(_15523_),
    .A2(_15525_),
    .ZN(_15526_)
  );
  INV_X1 _50710_ (
    .A(_15526_),
    .ZN(_01011_)
  );
  AND2_X1 _50711_ (
    .A1(_12776_),
    .A2(_13169_),
    .ZN(_15527_)
  );
  INV_X1 _50712_ (
    .A(_15527_),
    .ZN(_15528_)
  );
  AND2_X1 _50713_ (
    .A1(\cpuregs[20] [20]),
    .A2(_12777_),
    .ZN(_15529_)
  );
  INV_X1 _50714_ (
    .A(_15529_),
    .ZN(_15530_)
  );
  AND2_X1 _50715_ (
    .A1(_15528_),
    .A2(_15530_),
    .ZN(_15531_)
  );
  INV_X1 _50716_ (
    .A(_15531_),
    .ZN(_01012_)
  );
  AND2_X1 _50717_ (
    .A1(_12776_),
    .A2(_13184_),
    .ZN(_15532_)
  );
  INV_X1 _50718_ (
    .A(_15532_),
    .ZN(_15533_)
  );
  AND2_X1 _50719_ (
    .A1(\cpuregs[20] [21]),
    .A2(_12777_),
    .ZN(_15534_)
  );
  INV_X1 _50720_ (
    .A(_15534_),
    .ZN(_15535_)
  );
  AND2_X1 _50721_ (
    .A1(_15533_),
    .A2(_15535_),
    .ZN(_15536_)
  );
  INV_X1 _50722_ (
    .A(_15536_),
    .ZN(_01013_)
  );
  AND2_X1 _50723_ (
    .A1(_12776_),
    .A2(_13199_),
    .ZN(_15537_)
  );
  INV_X1 _50724_ (
    .A(_15537_),
    .ZN(_15538_)
  );
  AND2_X1 _50725_ (
    .A1(\cpuregs[20] [22]),
    .A2(_12777_),
    .ZN(_15539_)
  );
  INV_X1 _50726_ (
    .A(_15539_),
    .ZN(_15540_)
  );
  AND2_X1 _50727_ (
    .A1(_15538_),
    .A2(_15540_),
    .ZN(_15541_)
  );
  INV_X1 _50728_ (
    .A(_15541_),
    .ZN(_01014_)
  );
  AND2_X1 _50729_ (
    .A1(_12776_),
    .A2(_13214_),
    .ZN(_15542_)
  );
  INV_X1 _50730_ (
    .A(_15542_),
    .ZN(_15543_)
  );
  AND2_X1 _50731_ (
    .A1(\cpuregs[20] [23]),
    .A2(_12777_),
    .ZN(_15544_)
  );
  INV_X1 _50732_ (
    .A(_15544_),
    .ZN(_15545_)
  );
  AND2_X1 _50733_ (
    .A1(_15543_),
    .A2(_15545_),
    .ZN(_15546_)
  );
  INV_X1 _50734_ (
    .A(_15546_),
    .ZN(_01015_)
  );
  AND2_X1 _50735_ (
    .A1(_12776_),
    .A2(_13229_),
    .ZN(_15547_)
  );
  INV_X1 _50736_ (
    .A(_15547_),
    .ZN(_15548_)
  );
  AND2_X1 _50737_ (
    .A1(\cpuregs[20] [24]),
    .A2(_12777_),
    .ZN(_15549_)
  );
  INV_X1 _50738_ (
    .A(_15549_),
    .ZN(_15550_)
  );
  AND2_X1 _50739_ (
    .A1(_15548_),
    .A2(_15550_),
    .ZN(_15551_)
  );
  INV_X1 _50740_ (
    .A(_15551_),
    .ZN(_01016_)
  );
  AND2_X1 _50741_ (
    .A1(_12776_),
    .A2(_13244_),
    .ZN(_15552_)
  );
  INV_X1 _50742_ (
    .A(_15552_),
    .ZN(_15553_)
  );
  AND2_X1 _50743_ (
    .A1(\cpuregs[20] [25]),
    .A2(_12777_),
    .ZN(_15554_)
  );
  INV_X1 _50744_ (
    .A(_15554_),
    .ZN(_15555_)
  );
  AND2_X1 _50745_ (
    .A1(_15553_),
    .A2(_15555_),
    .ZN(_15556_)
  );
  INV_X1 _50746_ (
    .A(_15556_),
    .ZN(_01017_)
  );
  AND2_X1 _50747_ (
    .A1(_12776_),
    .A2(_13259_),
    .ZN(_15557_)
  );
  INV_X1 _50748_ (
    .A(_15557_),
    .ZN(_15558_)
  );
  AND2_X1 _50749_ (
    .A1(\cpuregs[20] [26]),
    .A2(_12777_),
    .ZN(_15559_)
  );
  INV_X1 _50750_ (
    .A(_15559_),
    .ZN(_15560_)
  );
  AND2_X1 _50751_ (
    .A1(_15558_),
    .A2(_15560_),
    .ZN(_15561_)
  );
  INV_X1 _50752_ (
    .A(_15561_),
    .ZN(_01018_)
  );
  AND2_X1 _50753_ (
    .A1(_12776_),
    .A2(_13274_),
    .ZN(_15562_)
  );
  INV_X1 _50754_ (
    .A(_15562_),
    .ZN(_15563_)
  );
  AND2_X1 _50755_ (
    .A1(\cpuregs[20] [27]),
    .A2(_12777_),
    .ZN(_15564_)
  );
  INV_X1 _50756_ (
    .A(_15564_),
    .ZN(_15565_)
  );
  AND2_X1 _50757_ (
    .A1(_15563_),
    .A2(_15565_),
    .ZN(_15566_)
  );
  INV_X1 _50758_ (
    .A(_15566_),
    .ZN(_01019_)
  );
  AND2_X1 _50759_ (
    .A1(_12776_),
    .A2(_13289_),
    .ZN(_15567_)
  );
  INV_X1 _50760_ (
    .A(_15567_),
    .ZN(_15568_)
  );
  AND2_X1 _50761_ (
    .A1(\cpuregs[20] [28]),
    .A2(_12777_),
    .ZN(_15569_)
  );
  INV_X1 _50762_ (
    .A(_15569_),
    .ZN(_15570_)
  );
  AND2_X1 _50763_ (
    .A1(_15568_),
    .A2(_15570_),
    .ZN(_15571_)
  );
  INV_X1 _50764_ (
    .A(_15571_),
    .ZN(_01020_)
  );
  AND2_X1 _50765_ (
    .A1(_12776_),
    .A2(_13304_),
    .ZN(_15572_)
  );
  INV_X1 _50766_ (
    .A(_15572_),
    .ZN(_15573_)
  );
  AND2_X1 _50767_ (
    .A1(\cpuregs[20] [29]),
    .A2(_12777_),
    .ZN(_15574_)
  );
  INV_X1 _50768_ (
    .A(_15574_),
    .ZN(_15575_)
  );
  AND2_X1 _50769_ (
    .A1(_15573_),
    .A2(_15575_),
    .ZN(_15576_)
  );
  INV_X1 _50770_ (
    .A(_15576_),
    .ZN(_01021_)
  );
  AND2_X1 _50771_ (
    .A1(_12776_),
    .A2(_13319_),
    .ZN(_15577_)
  );
  INV_X1 _50772_ (
    .A(_15577_),
    .ZN(_15578_)
  );
  AND2_X1 _50773_ (
    .A1(\cpuregs[20] [30]),
    .A2(_12777_),
    .ZN(_15579_)
  );
  INV_X1 _50774_ (
    .A(_15579_),
    .ZN(_15580_)
  );
  AND2_X1 _50775_ (
    .A1(_15578_),
    .A2(_15580_),
    .ZN(_15581_)
  );
  INV_X1 _50776_ (
    .A(_15581_),
    .ZN(_01022_)
  );
  AND2_X1 _50777_ (
    .A1(_12672_),
    .A2(_12874_),
    .ZN(_15582_)
  );
  INV_X1 _50778_ (
    .A(_15582_),
    .ZN(_15583_)
  );
  AND2_X1 _50779_ (
    .A1(\cpuregs[4] [0]),
    .A2(_12673_),
    .ZN(_15584_)
  );
  INV_X1 _50780_ (
    .A(_15584_),
    .ZN(_15585_)
  );
  AND2_X1 _50781_ (
    .A1(_15583_),
    .A2(_15585_),
    .ZN(_15586_)
  );
  INV_X1 _50782_ (
    .A(_15586_),
    .ZN(_01023_)
  );
  AND2_X1 _50783_ (
    .A1(\cpuregs[4] [1]),
    .A2(_12673_),
    .ZN(_15587_)
  );
  INV_X1 _50784_ (
    .A(_15587_),
    .ZN(_15588_)
  );
  AND2_X1 _50785_ (
    .A1(_12672_),
    .A2(_12886_),
    .ZN(_15589_)
  );
  INV_X1 _50786_ (
    .A(_15589_),
    .ZN(_15590_)
  );
  AND2_X1 _50787_ (
    .A1(_15588_),
    .A2(_15590_),
    .ZN(_15591_)
  );
  INV_X1 _50788_ (
    .A(_15591_),
    .ZN(_01024_)
  );
  AND2_X1 _50789_ (
    .A1(_12672_),
    .A2(_12900_),
    .ZN(_15592_)
  );
  INV_X1 _50790_ (
    .A(_15592_),
    .ZN(_15593_)
  );
  AND2_X1 _50791_ (
    .A1(\cpuregs[4] [2]),
    .A2(_12673_),
    .ZN(_15594_)
  );
  INV_X1 _50792_ (
    .A(_15594_),
    .ZN(_15595_)
  );
  AND2_X1 _50793_ (
    .A1(_15593_),
    .A2(_15595_),
    .ZN(_15596_)
  );
  INV_X1 _50794_ (
    .A(_15596_),
    .ZN(_01025_)
  );
  AND2_X1 _50795_ (
    .A1(_12672_),
    .A2(_12913_),
    .ZN(_15597_)
  );
  INV_X1 _50796_ (
    .A(_15597_),
    .ZN(_15598_)
  );
  AND2_X1 _50797_ (
    .A1(\cpuregs[4] [3]),
    .A2(_12673_),
    .ZN(_15599_)
  );
  INV_X1 _50798_ (
    .A(_15599_),
    .ZN(_15600_)
  );
  AND2_X1 _50799_ (
    .A1(_15598_),
    .A2(_15600_),
    .ZN(_15601_)
  );
  INV_X1 _50800_ (
    .A(_15601_),
    .ZN(_01026_)
  );
  AND2_X1 _50801_ (
    .A1(_12672_),
    .A2(_12928_),
    .ZN(_15602_)
  );
  INV_X1 _50802_ (
    .A(_15602_),
    .ZN(_15603_)
  );
  AND2_X1 _50803_ (
    .A1(\cpuregs[4] [4]),
    .A2(_12673_),
    .ZN(_15604_)
  );
  INV_X1 _50804_ (
    .A(_15604_),
    .ZN(_15605_)
  );
  AND2_X1 _50805_ (
    .A1(_15603_),
    .A2(_15605_),
    .ZN(_15606_)
  );
  INV_X1 _50806_ (
    .A(_15606_),
    .ZN(_01027_)
  );
  AND2_X1 _50807_ (
    .A1(_12672_),
    .A2(_12943_),
    .ZN(_15607_)
  );
  INV_X1 _50808_ (
    .A(_15607_),
    .ZN(_15608_)
  );
  AND2_X1 _50809_ (
    .A1(\cpuregs[4] [5]),
    .A2(_12673_),
    .ZN(_15609_)
  );
  INV_X1 _50810_ (
    .A(_15609_),
    .ZN(_15610_)
  );
  AND2_X1 _50811_ (
    .A1(_15608_),
    .A2(_15610_),
    .ZN(_15611_)
  );
  INV_X1 _50812_ (
    .A(_15611_),
    .ZN(_01028_)
  );
  AND2_X1 _50813_ (
    .A1(_12672_),
    .A2(_12958_),
    .ZN(_15612_)
  );
  INV_X1 _50814_ (
    .A(_15612_),
    .ZN(_15613_)
  );
  AND2_X1 _50815_ (
    .A1(\cpuregs[4] [6]),
    .A2(_12673_),
    .ZN(_15614_)
  );
  INV_X1 _50816_ (
    .A(_15614_),
    .ZN(_15615_)
  );
  AND2_X1 _50817_ (
    .A1(_15613_),
    .A2(_15615_),
    .ZN(_15616_)
  );
  INV_X1 _50818_ (
    .A(_15616_),
    .ZN(_01029_)
  );
  AND2_X1 _50819_ (
    .A1(_12672_),
    .A2(_12973_),
    .ZN(_15617_)
  );
  INV_X1 _50820_ (
    .A(_15617_),
    .ZN(_15618_)
  );
  AND2_X1 _50821_ (
    .A1(\cpuregs[4] [7]),
    .A2(_12673_),
    .ZN(_15619_)
  );
  INV_X1 _50822_ (
    .A(_15619_),
    .ZN(_15620_)
  );
  AND2_X1 _50823_ (
    .A1(_15618_),
    .A2(_15620_),
    .ZN(_15621_)
  );
  INV_X1 _50824_ (
    .A(_15621_),
    .ZN(_01030_)
  );
  AND2_X1 _50825_ (
    .A1(_12672_),
    .A2(_12988_),
    .ZN(_15622_)
  );
  INV_X1 _50826_ (
    .A(_15622_),
    .ZN(_15623_)
  );
  AND2_X1 _50827_ (
    .A1(\cpuregs[4] [8]),
    .A2(_12673_),
    .ZN(_15624_)
  );
  INV_X1 _50828_ (
    .A(_15624_),
    .ZN(_15625_)
  );
  AND2_X1 _50829_ (
    .A1(_15623_),
    .A2(_15625_),
    .ZN(_15626_)
  );
  INV_X1 _50830_ (
    .A(_15626_),
    .ZN(_01031_)
  );
  AND2_X1 _50831_ (
    .A1(_12672_),
    .A2(_13003_),
    .ZN(_15627_)
  );
  INV_X1 _50832_ (
    .A(_15627_),
    .ZN(_15628_)
  );
  AND2_X1 _50833_ (
    .A1(\cpuregs[4] [9]),
    .A2(_12673_),
    .ZN(_15629_)
  );
  INV_X1 _50834_ (
    .A(_15629_),
    .ZN(_15630_)
  );
  AND2_X1 _50835_ (
    .A1(_15628_),
    .A2(_15630_),
    .ZN(_15631_)
  );
  INV_X1 _50836_ (
    .A(_15631_),
    .ZN(_01032_)
  );
  AND2_X1 _50837_ (
    .A1(_12672_),
    .A2(_13018_),
    .ZN(_15632_)
  );
  INV_X1 _50838_ (
    .A(_15632_),
    .ZN(_15633_)
  );
  AND2_X1 _50839_ (
    .A1(\cpuregs[4] [10]),
    .A2(_12673_),
    .ZN(_15634_)
  );
  INV_X1 _50840_ (
    .A(_15634_),
    .ZN(_15635_)
  );
  AND2_X1 _50841_ (
    .A1(_15633_),
    .A2(_15635_),
    .ZN(_15636_)
  );
  INV_X1 _50842_ (
    .A(_15636_),
    .ZN(_01033_)
  );
  AND2_X1 _50843_ (
    .A1(_12672_),
    .A2(_13033_),
    .ZN(_15637_)
  );
  INV_X1 _50844_ (
    .A(_15637_),
    .ZN(_15638_)
  );
  AND2_X1 _50845_ (
    .A1(\cpuregs[4] [11]),
    .A2(_12673_),
    .ZN(_15639_)
  );
  INV_X1 _50846_ (
    .A(_15639_),
    .ZN(_15640_)
  );
  AND2_X1 _50847_ (
    .A1(_15638_),
    .A2(_15640_),
    .ZN(_15641_)
  );
  INV_X1 _50848_ (
    .A(_15641_),
    .ZN(_01034_)
  );
  AND2_X1 _50849_ (
    .A1(_12672_),
    .A2(_13048_),
    .ZN(_15642_)
  );
  INV_X1 _50850_ (
    .A(_15642_),
    .ZN(_15643_)
  );
  AND2_X1 _50851_ (
    .A1(\cpuregs[4] [12]),
    .A2(_12673_),
    .ZN(_15644_)
  );
  INV_X1 _50852_ (
    .A(_15644_),
    .ZN(_15645_)
  );
  AND2_X1 _50853_ (
    .A1(_15643_),
    .A2(_15645_),
    .ZN(_15646_)
  );
  INV_X1 _50854_ (
    .A(_15646_),
    .ZN(_01035_)
  );
  AND2_X1 _50855_ (
    .A1(_12672_),
    .A2(_13063_),
    .ZN(_15647_)
  );
  INV_X1 _50856_ (
    .A(_15647_),
    .ZN(_15648_)
  );
  AND2_X1 _50857_ (
    .A1(\cpuregs[4] [13]),
    .A2(_12673_),
    .ZN(_15649_)
  );
  INV_X1 _50858_ (
    .A(_15649_),
    .ZN(_15650_)
  );
  AND2_X1 _50859_ (
    .A1(_15648_),
    .A2(_15650_),
    .ZN(_15651_)
  );
  INV_X1 _50860_ (
    .A(_15651_),
    .ZN(_01036_)
  );
  AND2_X1 _50861_ (
    .A1(\cpuregs[4] [14]),
    .A2(_12673_),
    .ZN(_15652_)
  );
  INV_X1 _50862_ (
    .A(_15652_),
    .ZN(_15653_)
  );
  AND2_X1 _50863_ (
    .A1(_12672_),
    .A2(_13078_),
    .ZN(_15654_)
  );
  INV_X1 _50864_ (
    .A(_15654_),
    .ZN(_15655_)
  );
  AND2_X1 _50865_ (
    .A1(_15653_),
    .A2(_15655_),
    .ZN(_15656_)
  );
  INV_X1 _50866_ (
    .A(_15656_),
    .ZN(_01037_)
  );
  AND2_X1 _50867_ (
    .A1(_12672_),
    .A2(_13093_),
    .ZN(_15657_)
  );
  INV_X1 _50868_ (
    .A(_15657_),
    .ZN(_15658_)
  );
  AND2_X1 _50869_ (
    .A1(\cpuregs[4] [15]),
    .A2(_12673_),
    .ZN(_15659_)
  );
  INV_X1 _50870_ (
    .A(_15659_),
    .ZN(_15660_)
  );
  AND2_X1 _50871_ (
    .A1(_15658_),
    .A2(_15660_),
    .ZN(_15661_)
  );
  INV_X1 _50872_ (
    .A(_15661_),
    .ZN(_01038_)
  );
  AND2_X1 _50873_ (
    .A1(_12672_),
    .A2(_13108_),
    .ZN(_15662_)
  );
  INV_X1 _50874_ (
    .A(_15662_),
    .ZN(_15663_)
  );
  AND2_X1 _50875_ (
    .A1(\cpuregs[4] [16]),
    .A2(_12673_),
    .ZN(_15664_)
  );
  INV_X1 _50876_ (
    .A(_15664_),
    .ZN(_15665_)
  );
  AND2_X1 _50877_ (
    .A1(_15663_),
    .A2(_15665_),
    .ZN(_15666_)
  );
  INV_X1 _50878_ (
    .A(_15666_),
    .ZN(_01039_)
  );
  AND2_X1 _50879_ (
    .A1(_12672_),
    .A2(_13123_),
    .ZN(_15667_)
  );
  INV_X1 _50880_ (
    .A(_15667_),
    .ZN(_15668_)
  );
  AND2_X1 _50881_ (
    .A1(\cpuregs[4] [17]),
    .A2(_12673_),
    .ZN(_15669_)
  );
  INV_X1 _50882_ (
    .A(_15669_),
    .ZN(_15670_)
  );
  AND2_X1 _50883_ (
    .A1(_15668_),
    .A2(_15670_),
    .ZN(_15671_)
  );
  INV_X1 _50884_ (
    .A(_15671_),
    .ZN(_01040_)
  );
  AND2_X1 _50885_ (
    .A1(_12672_),
    .A2(_13139_),
    .ZN(_15672_)
  );
  INV_X1 _50886_ (
    .A(_15672_),
    .ZN(_15673_)
  );
  AND2_X1 _50887_ (
    .A1(\cpuregs[4] [18]),
    .A2(_12673_),
    .ZN(_15674_)
  );
  INV_X1 _50888_ (
    .A(_15674_),
    .ZN(_15675_)
  );
  AND2_X1 _50889_ (
    .A1(_15673_),
    .A2(_15675_),
    .ZN(_15676_)
  );
  INV_X1 _50890_ (
    .A(_15676_),
    .ZN(_01041_)
  );
  AND2_X1 _50891_ (
    .A1(_12672_),
    .A2(_13154_),
    .ZN(_15677_)
  );
  INV_X1 _50892_ (
    .A(_15677_),
    .ZN(_15678_)
  );
  AND2_X1 _50893_ (
    .A1(\cpuregs[4] [19]),
    .A2(_12673_),
    .ZN(_15679_)
  );
  INV_X1 _50894_ (
    .A(_15679_),
    .ZN(_15680_)
  );
  AND2_X1 _50895_ (
    .A1(_15678_),
    .A2(_15680_),
    .ZN(_15681_)
  );
  INV_X1 _50896_ (
    .A(_15681_),
    .ZN(_01042_)
  );
  AND2_X1 _50897_ (
    .A1(_12672_),
    .A2(_13169_),
    .ZN(_15682_)
  );
  INV_X1 _50898_ (
    .A(_15682_),
    .ZN(_15683_)
  );
  AND2_X1 _50899_ (
    .A1(\cpuregs[4] [20]),
    .A2(_12673_),
    .ZN(_15684_)
  );
  INV_X1 _50900_ (
    .A(_15684_),
    .ZN(_15685_)
  );
  AND2_X1 _50901_ (
    .A1(_15683_),
    .A2(_15685_),
    .ZN(_15686_)
  );
  INV_X1 _50902_ (
    .A(_15686_),
    .ZN(_01043_)
  );
  AND2_X1 _50903_ (
    .A1(_12672_),
    .A2(_13184_),
    .ZN(_15687_)
  );
  INV_X1 _50904_ (
    .A(_15687_),
    .ZN(_15688_)
  );
  AND2_X1 _50905_ (
    .A1(\cpuregs[4] [21]),
    .A2(_12673_),
    .ZN(_15689_)
  );
  INV_X1 _50906_ (
    .A(_15689_),
    .ZN(_15690_)
  );
  AND2_X1 _50907_ (
    .A1(_15688_),
    .A2(_15690_),
    .ZN(_15691_)
  );
  INV_X1 _50908_ (
    .A(_15691_),
    .ZN(_01044_)
  );
  AND2_X1 _50909_ (
    .A1(_12672_),
    .A2(_13199_),
    .ZN(_15692_)
  );
  INV_X1 _50910_ (
    .A(_15692_),
    .ZN(_15693_)
  );
  AND2_X1 _50911_ (
    .A1(\cpuregs[4] [22]),
    .A2(_12673_),
    .ZN(_15694_)
  );
  INV_X1 _50912_ (
    .A(_15694_),
    .ZN(_15695_)
  );
  AND2_X1 _50913_ (
    .A1(_15693_),
    .A2(_15695_),
    .ZN(_15696_)
  );
  INV_X1 _50914_ (
    .A(_15696_),
    .ZN(_01045_)
  );
  AND2_X1 _50915_ (
    .A1(_12672_),
    .A2(_13214_),
    .ZN(_15697_)
  );
  INV_X1 _50916_ (
    .A(_15697_),
    .ZN(_15698_)
  );
  AND2_X1 _50917_ (
    .A1(\cpuregs[4] [23]),
    .A2(_12673_),
    .ZN(_15699_)
  );
  INV_X1 _50918_ (
    .A(_15699_),
    .ZN(_15700_)
  );
  AND2_X1 _50919_ (
    .A1(_15698_),
    .A2(_15700_),
    .ZN(_15701_)
  );
  INV_X1 _50920_ (
    .A(_15701_),
    .ZN(_01046_)
  );
  AND2_X1 _50921_ (
    .A1(_12672_),
    .A2(_13229_),
    .ZN(_15702_)
  );
  INV_X1 _50922_ (
    .A(_15702_),
    .ZN(_15703_)
  );
  AND2_X1 _50923_ (
    .A1(\cpuregs[4] [24]),
    .A2(_12673_),
    .ZN(_15704_)
  );
  INV_X1 _50924_ (
    .A(_15704_),
    .ZN(_15705_)
  );
  AND2_X1 _50925_ (
    .A1(_15703_),
    .A2(_15705_),
    .ZN(_15706_)
  );
  INV_X1 _50926_ (
    .A(_15706_),
    .ZN(_01047_)
  );
  AND2_X1 _50927_ (
    .A1(_12672_),
    .A2(_13244_),
    .ZN(_15707_)
  );
  INV_X1 _50928_ (
    .A(_15707_),
    .ZN(_15708_)
  );
  AND2_X1 _50929_ (
    .A1(\cpuregs[4] [25]),
    .A2(_12673_),
    .ZN(_15709_)
  );
  INV_X1 _50930_ (
    .A(_15709_),
    .ZN(_15710_)
  );
  AND2_X1 _50931_ (
    .A1(_15708_),
    .A2(_15710_),
    .ZN(_15711_)
  );
  INV_X1 _50932_ (
    .A(_15711_),
    .ZN(_01048_)
  );
  AND2_X1 _50933_ (
    .A1(_12672_),
    .A2(_13259_),
    .ZN(_15712_)
  );
  INV_X1 _50934_ (
    .A(_15712_),
    .ZN(_15713_)
  );
  AND2_X1 _50935_ (
    .A1(\cpuregs[4] [26]),
    .A2(_12673_),
    .ZN(_15714_)
  );
  INV_X1 _50936_ (
    .A(_15714_),
    .ZN(_15715_)
  );
  AND2_X1 _50937_ (
    .A1(_15713_),
    .A2(_15715_),
    .ZN(_15716_)
  );
  INV_X1 _50938_ (
    .A(_15716_),
    .ZN(_01049_)
  );
  AND2_X1 _50939_ (
    .A1(_12672_),
    .A2(_13274_),
    .ZN(_15717_)
  );
  INV_X1 _50940_ (
    .A(_15717_),
    .ZN(_15718_)
  );
  AND2_X1 _50941_ (
    .A1(\cpuregs[4] [27]),
    .A2(_12673_),
    .ZN(_15719_)
  );
  INV_X1 _50942_ (
    .A(_15719_),
    .ZN(_15720_)
  );
  AND2_X1 _50943_ (
    .A1(_15718_),
    .A2(_15720_),
    .ZN(_15721_)
  );
  INV_X1 _50944_ (
    .A(_15721_),
    .ZN(_01050_)
  );
  AND2_X1 _50945_ (
    .A1(_12672_),
    .A2(_13289_),
    .ZN(_15722_)
  );
  INV_X1 _50946_ (
    .A(_15722_),
    .ZN(_15723_)
  );
  AND2_X1 _50947_ (
    .A1(\cpuregs[4] [28]),
    .A2(_12673_),
    .ZN(_15724_)
  );
  INV_X1 _50948_ (
    .A(_15724_),
    .ZN(_15725_)
  );
  AND2_X1 _50949_ (
    .A1(_15723_),
    .A2(_15725_),
    .ZN(_15726_)
  );
  INV_X1 _50950_ (
    .A(_15726_),
    .ZN(_01051_)
  );
  AND2_X1 _50951_ (
    .A1(_12672_),
    .A2(_13304_),
    .ZN(_15727_)
  );
  INV_X1 _50952_ (
    .A(_15727_),
    .ZN(_15728_)
  );
  AND2_X1 _50953_ (
    .A1(\cpuregs[4] [29]),
    .A2(_12673_),
    .ZN(_15729_)
  );
  INV_X1 _50954_ (
    .A(_15729_),
    .ZN(_15730_)
  );
  AND2_X1 _50955_ (
    .A1(_15728_),
    .A2(_15730_),
    .ZN(_15731_)
  );
  INV_X1 _50956_ (
    .A(_15731_),
    .ZN(_01052_)
  );
  AND2_X1 _50957_ (
    .A1(_12672_),
    .A2(_13319_),
    .ZN(_15732_)
  );
  INV_X1 _50958_ (
    .A(_15732_),
    .ZN(_15733_)
  );
  AND2_X1 _50959_ (
    .A1(\cpuregs[4] [30]),
    .A2(_12673_),
    .ZN(_15734_)
  );
  INV_X1 _50960_ (
    .A(_15734_),
    .ZN(_15735_)
  );
  AND2_X1 _50961_ (
    .A1(_15733_),
    .A2(_15735_),
    .ZN(_15736_)
  );
  INV_X1 _50962_ (
    .A(_15736_),
    .ZN(_01053_)
  );
  AND2_X1 _50963_ (
    .A1(_12856_),
    .A2(_12872_),
    .ZN(_15737_)
  );
  INV_X1 _50964_ (
    .A(_15737_),
    .ZN(_15738_)
  );
  AND2_X1 _50965_ (
    .A1(_21694_),
    .A2(_12857_),
    .ZN(_15739_)
  );
  INV_X1 _50966_ (
    .A(_15739_),
    .ZN(_15740_)
  );
  AND2_X1 _50967_ (
    .A1(_15738_),
    .A2(_15740_),
    .ZN(_01054_)
  );
  AND2_X1 _50968_ (
    .A1(_12856_),
    .A2(_12884_),
    .ZN(_15741_)
  );
  INV_X1 _50969_ (
    .A(_15741_),
    .ZN(_15742_)
  );
  AND2_X1 _50970_ (
    .A1(_21695_),
    .A2(_12857_),
    .ZN(_15743_)
  );
  INV_X1 _50971_ (
    .A(_15743_),
    .ZN(_15744_)
  );
  AND2_X1 _50972_ (
    .A1(_15742_),
    .A2(_15744_),
    .ZN(_01055_)
  );
  AND2_X1 _50973_ (
    .A1(_12856_),
    .A2(_12898_),
    .ZN(_15745_)
  );
  INV_X1 _50974_ (
    .A(_15745_),
    .ZN(_15746_)
  );
  AND2_X1 _50975_ (
    .A1(_21696_),
    .A2(_12857_),
    .ZN(_15747_)
  );
  INV_X1 _50976_ (
    .A(_15747_),
    .ZN(_15748_)
  );
  AND2_X1 _50977_ (
    .A1(_15746_),
    .A2(_15748_),
    .ZN(_01056_)
  );
  AND2_X1 _50978_ (
    .A1(_12856_),
    .A2(_12911_),
    .ZN(_15749_)
  );
  INV_X1 _50979_ (
    .A(_15749_),
    .ZN(_15750_)
  );
  AND2_X1 _50980_ (
    .A1(_21697_),
    .A2(_12857_),
    .ZN(_15751_)
  );
  INV_X1 _50981_ (
    .A(_15751_),
    .ZN(_15752_)
  );
  AND2_X1 _50982_ (
    .A1(_15750_),
    .A2(_15752_),
    .ZN(_01057_)
  );
  AND2_X1 _50983_ (
    .A1(_12856_),
    .A2(_12928_),
    .ZN(_15753_)
  );
  INV_X1 _50984_ (
    .A(_15753_),
    .ZN(_15754_)
  );
  AND2_X1 _50985_ (
    .A1(\cpuregs[10] [4]),
    .A2(_12857_),
    .ZN(_15755_)
  );
  INV_X1 _50986_ (
    .A(_15755_),
    .ZN(_15756_)
  );
  AND2_X1 _50987_ (
    .A1(_15754_),
    .A2(_15756_),
    .ZN(_15757_)
  );
  INV_X1 _50988_ (
    .A(_15757_),
    .ZN(_01058_)
  );
  AND2_X1 _50989_ (
    .A1(_12856_),
    .A2(_12941_),
    .ZN(_15758_)
  );
  INV_X1 _50990_ (
    .A(_15758_),
    .ZN(_15759_)
  );
  AND2_X1 _50991_ (
    .A1(_21698_),
    .A2(_12857_),
    .ZN(_15760_)
  );
  INV_X1 _50992_ (
    .A(_15760_),
    .ZN(_15761_)
  );
  AND2_X1 _50993_ (
    .A1(_15759_),
    .A2(_15761_),
    .ZN(_01059_)
  );
  AND2_X1 _50994_ (
    .A1(_12856_),
    .A2(_12956_),
    .ZN(_15762_)
  );
  INV_X1 _50995_ (
    .A(_15762_),
    .ZN(_15763_)
  );
  AND2_X1 _50996_ (
    .A1(_21699_),
    .A2(_12857_),
    .ZN(_15764_)
  );
  INV_X1 _50997_ (
    .A(_15764_),
    .ZN(_15765_)
  );
  AND2_X1 _50998_ (
    .A1(_15763_),
    .A2(_15765_),
    .ZN(_01060_)
  );
  AND2_X1 _50999_ (
    .A1(_12856_),
    .A2(_12971_),
    .ZN(_15766_)
  );
  INV_X1 _51000_ (
    .A(_15766_),
    .ZN(_15767_)
  );
  AND2_X1 _51001_ (
    .A1(_21700_),
    .A2(_12857_),
    .ZN(_15768_)
  );
  INV_X1 _51002_ (
    .A(_15768_),
    .ZN(_15769_)
  );
  AND2_X1 _51003_ (
    .A1(_15767_),
    .A2(_15769_),
    .ZN(_01061_)
  );
  AND2_X1 _51004_ (
    .A1(_12856_),
    .A2(_12988_),
    .ZN(_15770_)
  );
  INV_X1 _51005_ (
    .A(_15770_),
    .ZN(_15771_)
  );
  AND2_X1 _51006_ (
    .A1(\cpuregs[10] [8]),
    .A2(_12857_),
    .ZN(_15772_)
  );
  INV_X1 _51007_ (
    .A(_15772_),
    .ZN(_15773_)
  );
  AND2_X1 _51008_ (
    .A1(_15771_),
    .A2(_15773_),
    .ZN(_15774_)
  );
  INV_X1 _51009_ (
    .A(_15774_),
    .ZN(_01062_)
  );
  AND2_X1 _51010_ (
    .A1(_12856_),
    .A2(_13001_),
    .ZN(_15775_)
  );
  INV_X1 _51011_ (
    .A(_15775_),
    .ZN(_15776_)
  );
  AND2_X1 _51012_ (
    .A1(_21701_),
    .A2(_12857_),
    .ZN(_15777_)
  );
  INV_X1 _51013_ (
    .A(_15777_),
    .ZN(_15778_)
  );
  AND2_X1 _51014_ (
    .A1(_15776_),
    .A2(_15778_),
    .ZN(_01063_)
  );
  AND2_X1 _51015_ (
    .A1(_12856_),
    .A2(_13016_),
    .ZN(_15779_)
  );
  INV_X1 _51016_ (
    .A(_15779_),
    .ZN(_15780_)
  );
  AND2_X1 _51017_ (
    .A1(_21702_),
    .A2(_12857_),
    .ZN(_15781_)
  );
  INV_X1 _51018_ (
    .A(_15781_),
    .ZN(_15782_)
  );
  AND2_X1 _51019_ (
    .A1(_15780_),
    .A2(_15782_),
    .ZN(_01064_)
  );
  AND2_X1 _51020_ (
    .A1(_12856_),
    .A2(_13031_),
    .ZN(_15783_)
  );
  INV_X1 _51021_ (
    .A(_15783_),
    .ZN(_15784_)
  );
  AND2_X1 _51022_ (
    .A1(_21703_),
    .A2(_12857_),
    .ZN(_15785_)
  );
  INV_X1 _51023_ (
    .A(_15785_),
    .ZN(_15786_)
  );
  AND2_X1 _51024_ (
    .A1(_15784_),
    .A2(_15786_),
    .ZN(_01065_)
  );
  AND2_X1 _51025_ (
    .A1(_12856_),
    .A2(_13046_),
    .ZN(_15787_)
  );
  INV_X1 _51026_ (
    .A(_15787_),
    .ZN(_15788_)
  );
  AND2_X1 _51027_ (
    .A1(_21704_),
    .A2(_12857_),
    .ZN(_15789_)
  );
  INV_X1 _51028_ (
    .A(_15789_),
    .ZN(_15790_)
  );
  AND2_X1 _51029_ (
    .A1(_15788_),
    .A2(_15790_),
    .ZN(_01066_)
  );
  AND2_X1 _51030_ (
    .A1(_12856_),
    .A2(_13061_),
    .ZN(_15791_)
  );
  INV_X1 _51031_ (
    .A(_15791_),
    .ZN(_15792_)
  );
  AND2_X1 _51032_ (
    .A1(_21705_),
    .A2(_12857_),
    .ZN(_15793_)
  );
  INV_X1 _51033_ (
    .A(_15793_),
    .ZN(_15794_)
  );
  AND2_X1 _51034_ (
    .A1(_15792_),
    .A2(_15794_),
    .ZN(_01067_)
  );
  AND2_X1 _51035_ (
    .A1(_12856_),
    .A2(_13078_),
    .ZN(_15795_)
  );
  INV_X1 _51036_ (
    .A(_15795_),
    .ZN(_15796_)
  );
  AND2_X1 _51037_ (
    .A1(\cpuregs[10] [14]),
    .A2(_12857_),
    .ZN(_15797_)
  );
  INV_X1 _51038_ (
    .A(_15797_),
    .ZN(_15798_)
  );
  AND2_X1 _51039_ (
    .A1(_15796_),
    .A2(_15798_),
    .ZN(_15799_)
  );
  INV_X1 _51040_ (
    .A(_15799_),
    .ZN(_01068_)
  );
  AND2_X1 _51041_ (
    .A1(_12856_),
    .A2(_13091_),
    .ZN(_15800_)
  );
  INV_X1 _51042_ (
    .A(_15800_),
    .ZN(_15801_)
  );
  AND2_X1 _51043_ (
    .A1(_21706_),
    .A2(_12857_),
    .ZN(_15802_)
  );
  INV_X1 _51044_ (
    .A(_15802_),
    .ZN(_15803_)
  );
  AND2_X1 _51045_ (
    .A1(_15801_),
    .A2(_15803_),
    .ZN(_01069_)
  );
  AND2_X1 _51046_ (
    .A1(_12856_),
    .A2(_13108_),
    .ZN(_15804_)
  );
  INV_X1 _51047_ (
    .A(_15804_),
    .ZN(_15805_)
  );
  AND2_X1 _51048_ (
    .A1(\cpuregs[10] [16]),
    .A2(_12857_),
    .ZN(_15806_)
  );
  INV_X1 _51049_ (
    .A(_15806_),
    .ZN(_15807_)
  );
  AND2_X1 _51050_ (
    .A1(_15805_),
    .A2(_15807_),
    .ZN(_15808_)
  );
  INV_X1 _51051_ (
    .A(_15808_),
    .ZN(_01070_)
  );
  AND2_X1 _51052_ (
    .A1(_12856_),
    .A2(_13121_),
    .ZN(_15809_)
  );
  INV_X1 _51053_ (
    .A(_15809_),
    .ZN(_15810_)
  );
  AND2_X1 _51054_ (
    .A1(_21707_),
    .A2(_12857_),
    .ZN(_15811_)
  );
  INV_X1 _51055_ (
    .A(_15811_),
    .ZN(_15812_)
  );
  AND2_X1 _51056_ (
    .A1(_15810_),
    .A2(_15812_),
    .ZN(_01071_)
  );
  AND2_X1 _51057_ (
    .A1(_12856_),
    .A2(_13139_),
    .ZN(_15813_)
  );
  INV_X1 _51058_ (
    .A(_15813_),
    .ZN(_15814_)
  );
  AND2_X1 _51059_ (
    .A1(\cpuregs[10] [18]),
    .A2(_12857_),
    .ZN(_15815_)
  );
  INV_X1 _51060_ (
    .A(_15815_),
    .ZN(_15816_)
  );
  AND2_X1 _51061_ (
    .A1(_15814_),
    .A2(_15816_),
    .ZN(_15817_)
  );
  INV_X1 _51062_ (
    .A(_15817_),
    .ZN(_01072_)
  );
  AND2_X1 _51063_ (
    .A1(_12856_),
    .A2(_13152_),
    .ZN(_15818_)
  );
  INV_X1 _51064_ (
    .A(_15818_),
    .ZN(_15819_)
  );
  AND2_X1 _51065_ (
    .A1(_21708_),
    .A2(_12857_),
    .ZN(_15820_)
  );
  INV_X1 _51066_ (
    .A(_15820_),
    .ZN(_15821_)
  );
  AND2_X1 _51067_ (
    .A1(_15819_),
    .A2(_15821_),
    .ZN(_01073_)
  );
  AND2_X1 _51068_ (
    .A1(_12856_),
    .A2(_13169_),
    .ZN(_15822_)
  );
  INV_X1 _51069_ (
    .A(_15822_),
    .ZN(_15823_)
  );
  AND2_X1 _51070_ (
    .A1(\cpuregs[10] [20]),
    .A2(_12857_),
    .ZN(_15824_)
  );
  INV_X1 _51071_ (
    .A(_15824_),
    .ZN(_15825_)
  );
  AND2_X1 _51072_ (
    .A1(_15823_),
    .A2(_15825_),
    .ZN(_15826_)
  );
  INV_X1 _51073_ (
    .A(_15826_),
    .ZN(_01074_)
  );
  AND2_X1 _51074_ (
    .A1(_12856_),
    .A2(_13184_),
    .ZN(_15827_)
  );
  INV_X1 _51075_ (
    .A(_15827_),
    .ZN(_15828_)
  );
  AND2_X1 _51076_ (
    .A1(\cpuregs[10] [21]),
    .A2(_12857_),
    .ZN(_15829_)
  );
  INV_X1 _51077_ (
    .A(_15829_),
    .ZN(_15830_)
  );
  AND2_X1 _51078_ (
    .A1(_15828_),
    .A2(_15830_),
    .ZN(_15831_)
  );
  INV_X1 _51079_ (
    .A(_15831_),
    .ZN(_01075_)
  );
  AND2_X1 _51080_ (
    .A1(_12856_),
    .A2(_13197_),
    .ZN(_15832_)
  );
  INV_X1 _51081_ (
    .A(_15832_),
    .ZN(_15833_)
  );
  AND2_X1 _51082_ (
    .A1(_21709_),
    .A2(_12857_),
    .ZN(_15834_)
  );
  INV_X1 _51083_ (
    .A(_15834_),
    .ZN(_15835_)
  );
  AND2_X1 _51084_ (
    .A1(_15833_),
    .A2(_15835_),
    .ZN(_01076_)
  );
  AND2_X1 _51085_ (
    .A1(_12856_),
    .A2(_13212_),
    .ZN(_15836_)
  );
  INV_X1 _51086_ (
    .A(_15836_),
    .ZN(_15837_)
  );
  AND2_X1 _51087_ (
    .A1(_21710_),
    .A2(_12857_),
    .ZN(_15838_)
  );
  INV_X1 _51088_ (
    .A(_15838_),
    .ZN(_15839_)
  );
  AND2_X1 _51089_ (
    .A1(_15837_),
    .A2(_15839_),
    .ZN(_01077_)
  );
  AND2_X1 _51090_ (
    .A1(_12856_),
    .A2(_13229_),
    .ZN(_15840_)
  );
  INV_X1 _51091_ (
    .A(_15840_),
    .ZN(_15841_)
  );
  AND2_X1 _51092_ (
    .A1(\cpuregs[10] [24]),
    .A2(_12857_),
    .ZN(_15842_)
  );
  INV_X1 _51093_ (
    .A(_15842_),
    .ZN(_15843_)
  );
  AND2_X1 _51094_ (
    .A1(_15841_),
    .A2(_15843_),
    .ZN(_15844_)
  );
  INV_X1 _51095_ (
    .A(_15844_),
    .ZN(_01078_)
  );
  AND2_X1 _51096_ (
    .A1(_12856_),
    .A2(_13242_),
    .ZN(_15845_)
  );
  INV_X1 _51097_ (
    .A(_15845_),
    .ZN(_15846_)
  );
  AND2_X1 _51098_ (
    .A1(_21711_),
    .A2(_12857_),
    .ZN(_15847_)
  );
  INV_X1 _51099_ (
    .A(_15847_),
    .ZN(_15848_)
  );
  AND2_X1 _51100_ (
    .A1(_15846_),
    .A2(_15848_),
    .ZN(_01079_)
  );
  AND2_X1 _51101_ (
    .A1(_12856_),
    .A2(_13257_),
    .ZN(_15849_)
  );
  INV_X1 _51102_ (
    .A(_15849_),
    .ZN(_15850_)
  );
  AND2_X1 _51103_ (
    .A1(_21712_),
    .A2(_12857_),
    .ZN(_15851_)
  );
  INV_X1 _51104_ (
    .A(_15851_),
    .ZN(_15852_)
  );
  AND2_X1 _51105_ (
    .A1(_15850_),
    .A2(_15852_),
    .ZN(_01080_)
  );
  AND2_X1 _51106_ (
    .A1(_12856_),
    .A2(_13272_),
    .ZN(_15853_)
  );
  INV_X1 _51107_ (
    .A(_15853_),
    .ZN(_15854_)
  );
  AND2_X1 _51108_ (
    .A1(_21713_),
    .A2(_12857_),
    .ZN(_15855_)
  );
  INV_X1 _51109_ (
    .A(_15855_),
    .ZN(_15856_)
  );
  AND2_X1 _51110_ (
    .A1(_15854_),
    .A2(_15856_),
    .ZN(_01081_)
  );
  AND2_X1 _51111_ (
    .A1(_12856_),
    .A2(_13287_),
    .ZN(_15857_)
  );
  INV_X1 _51112_ (
    .A(_15857_),
    .ZN(_15858_)
  );
  AND2_X1 _51113_ (
    .A1(_21714_),
    .A2(_12857_),
    .ZN(_15859_)
  );
  INV_X1 _51114_ (
    .A(_15859_),
    .ZN(_15860_)
  );
  AND2_X1 _51115_ (
    .A1(_15858_),
    .A2(_15860_),
    .ZN(_01082_)
  );
  AND2_X1 _51116_ (
    .A1(_12856_),
    .A2(_13302_),
    .ZN(_15861_)
  );
  INV_X1 _51117_ (
    .A(_15861_),
    .ZN(_15862_)
  );
  AND2_X1 _51118_ (
    .A1(_21715_),
    .A2(_12857_),
    .ZN(_15863_)
  );
  INV_X1 _51119_ (
    .A(_15863_),
    .ZN(_15864_)
  );
  AND2_X1 _51120_ (
    .A1(_15862_),
    .A2(_15864_),
    .ZN(_01083_)
  );
  AND2_X1 _51121_ (
    .A1(_12856_),
    .A2(_13317_),
    .ZN(_15865_)
  );
  INV_X1 _51122_ (
    .A(_15865_),
    .ZN(_15866_)
  );
  AND2_X1 _51123_ (
    .A1(_21716_),
    .A2(_12857_),
    .ZN(_15867_)
  );
  INV_X1 _51124_ (
    .A(_15867_),
    .ZN(_15868_)
  );
  AND2_X1 _51125_ (
    .A1(_15866_),
    .A2(_15868_),
    .ZN(_01084_)
  );
  AND2_X1 _51126_ (
    .A1(_12559_),
    .A2(_12874_),
    .ZN(_15869_)
  );
  INV_X1 _51127_ (
    .A(_15869_),
    .ZN(_15870_)
  );
  AND2_X1 _51128_ (
    .A1(\cpuregs[9] [0]),
    .A2(_12560_),
    .ZN(_15871_)
  );
  INV_X1 _51129_ (
    .A(_15871_),
    .ZN(_15872_)
  );
  AND2_X1 _51130_ (
    .A1(_15870_),
    .A2(_15872_),
    .ZN(_15873_)
  );
  INV_X1 _51131_ (
    .A(_15873_),
    .ZN(_01085_)
  );
  AND2_X1 _51132_ (
    .A1(_12559_),
    .A2(_12886_),
    .ZN(_15874_)
  );
  INV_X1 _51133_ (
    .A(_15874_),
    .ZN(_15875_)
  );
  AND2_X1 _51134_ (
    .A1(\cpuregs[9] [1]),
    .A2(_12560_),
    .ZN(_15876_)
  );
  INV_X1 _51135_ (
    .A(_15876_),
    .ZN(_15877_)
  );
  AND2_X1 _51136_ (
    .A1(_15875_),
    .A2(_15877_),
    .ZN(_15878_)
  );
  INV_X1 _51137_ (
    .A(_15878_),
    .ZN(_01086_)
  );
  AND2_X1 _51138_ (
    .A1(\cpuregs[9] [2]),
    .A2(_12560_),
    .ZN(_15879_)
  );
  INV_X1 _51139_ (
    .A(_15879_),
    .ZN(_15880_)
  );
  AND2_X1 _51140_ (
    .A1(_12559_),
    .A2(_12900_),
    .ZN(_15881_)
  );
  INV_X1 _51141_ (
    .A(_15881_),
    .ZN(_15882_)
  );
  AND2_X1 _51142_ (
    .A1(_15880_),
    .A2(_15882_),
    .ZN(_15883_)
  );
  INV_X1 _51143_ (
    .A(_15883_),
    .ZN(_01087_)
  );
  AND2_X1 _51144_ (
    .A1(_12559_),
    .A2(_12913_),
    .ZN(_15884_)
  );
  INV_X1 _51145_ (
    .A(_15884_),
    .ZN(_15885_)
  );
  AND2_X1 _51146_ (
    .A1(\cpuregs[9] [3]),
    .A2(_12560_),
    .ZN(_15886_)
  );
  INV_X1 _51147_ (
    .A(_15886_),
    .ZN(_15887_)
  );
  AND2_X1 _51148_ (
    .A1(_15885_),
    .A2(_15887_),
    .ZN(_15888_)
  );
  INV_X1 _51149_ (
    .A(_15888_),
    .ZN(_01088_)
  );
  AND2_X1 _51150_ (
    .A1(\cpuregs[9] [4]),
    .A2(_12560_),
    .ZN(_15889_)
  );
  INV_X1 _51151_ (
    .A(_15889_),
    .ZN(_15890_)
  );
  AND2_X1 _51152_ (
    .A1(_12559_),
    .A2(_12928_),
    .ZN(_15891_)
  );
  INV_X1 _51153_ (
    .A(_15891_),
    .ZN(_15892_)
  );
  AND2_X1 _51154_ (
    .A1(_15890_),
    .A2(_15892_),
    .ZN(_15893_)
  );
  INV_X1 _51155_ (
    .A(_15893_),
    .ZN(_01089_)
  );
  AND2_X1 _51156_ (
    .A1(_12559_),
    .A2(_12943_),
    .ZN(_15894_)
  );
  INV_X1 _51157_ (
    .A(_15894_),
    .ZN(_15895_)
  );
  AND2_X1 _51158_ (
    .A1(\cpuregs[9] [5]),
    .A2(_12560_),
    .ZN(_15896_)
  );
  INV_X1 _51159_ (
    .A(_15896_),
    .ZN(_15897_)
  );
  AND2_X1 _51160_ (
    .A1(_15895_),
    .A2(_15897_),
    .ZN(_15898_)
  );
  INV_X1 _51161_ (
    .A(_15898_),
    .ZN(_01090_)
  );
  AND2_X1 _51162_ (
    .A1(_12559_),
    .A2(_12958_),
    .ZN(_15899_)
  );
  INV_X1 _51163_ (
    .A(_15899_),
    .ZN(_15900_)
  );
  AND2_X1 _51164_ (
    .A1(\cpuregs[9] [6]),
    .A2(_12560_),
    .ZN(_15901_)
  );
  INV_X1 _51165_ (
    .A(_15901_),
    .ZN(_15902_)
  );
  AND2_X1 _51166_ (
    .A1(_15900_),
    .A2(_15902_),
    .ZN(_15903_)
  );
  INV_X1 _51167_ (
    .A(_15903_),
    .ZN(_01091_)
  );
  AND2_X1 _51168_ (
    .A1(_12559_),
    .A2(_12973_),
    .ZN(_15904_)
  );
  INV_X1 _51169_ (
    .A(_15904_),
    .ZN(_15905_)
  );
  AND2_X1 _51170_ (
    .A1(\cpuregs[9] [7]),
    .A2(_12560_),
    .ZN(_15906_)
  );
  INV_X1 _51171_ (
    .A(_15906_),
    .ZN(_15907_)
  );
  AND2_X1 _51172_ (
    .A1(_15905_),
    .A2(_15907_),
    .ZN(_15908_)
  );
  INV_X1 _51173_ (
    .A(_15908_),
    .ZN(_01092_)
  );
  AND2_X1 _51174_ (
    .A1(_12559_),
    .A2(_12988_),
    .ZN(_15909_)
  );
  INV_X1 _51175_ (
    .A(_15909_),
    .ZN(_15910_)
  );
  AND2_X1 _51176_ (
    .A1(\cpuregs[9] [8]),
    .A2(_12560_),
    .ZN(_15911_)
  );
  INV_X1 _51177_ (
    .A(_15911_),
    .ZN(_15912_)
  );
  AND2_X1 _51178_ (
    .A1(_15910_),
    .A2(_15912_),
    .ZN(_15913_)
  );
  INV_X1 _51179_ (
    .A(_15913_),
    .ZN(_01093_)
  );
  AND2_X1 _51180_ (
    .A1(_12559_),
    .A2(_13003_),
    .ZN(_15914_)
  );
  INV_X1 _51181_ (
    .A(_15914_),
    .ZN(_15915_)
  );
  AND2_X1 _51182_ (
    .A1(\cpuregs[9] [9]),
    .A2(_12560_),
    .ZN(_15916_)
  );
  INV_X1 _51183_ (
    .A(_15916_),
    .ZN(_15917_)
  );
  AND2_X1 _51184_ (
    .A1(_15915_),
    .A2(_15917_),
    .ZN(_15918_)
  );
  INV_X1 _51185_ (
    .A(_15918_),
    .ZN(_01094_)
  );
  AND2_X1 _51186_ (
    .A1(_12559_),
    .A2(_13018_),
    .ZN(_15919_)
  );
  INV_X1 _51187_ (
    .A(_15919_),
    .ZN(_15920_)
  );
  AND2_X1 _51188_ (
    .A1(\cpuregs[9] [10]),
    .A2(_12560_),
    .ZN(_15921_)
  );
  INV_X1 _51189_ (
    .A(_15921_),
    .ZN(_15922_)
  );
  AND2_X1 _51190_ (
    .A1(_15920_),
    .A2(_15922_),
    .ZN(_15923_)
  );
  INV_X1 _51191_ (
    .A(_15923_),
    .ZN(_01095_)
  );
  AND2_X1 _51192_ (
    .A1(_12559_),
    .A2(_13033_),
    .ZN(_15924_)
  );
  INV_X1 _51193_ (
    .A(_15924_),
    .ZN(_15925_)
  );
  AND2_X1 _51194_ (
    .A1(\cpuregs[9] [11]),
    .A2(_12560_),
    .ZN(_15926_)
  );
  INV_X1 _51195_ (
    .A(_15926_),
    .ZN(_15927_)
  );
  AND2_X1 _51196_ (
    .A1(_15925_),
    .A2(_15927_),
    .ZN(_15928_)
  );
  INV_X1 _51197_ (
    .A(_15928_),
    .ZN(_01096_)
  );
  AND2_X1 _51198_ (
    .A1(_12559_),
    .A2(_13048_),
    .ZN(_15929_)
  );
  INV_X1 _51199_ (
    .A(_15929_),
    .ZN(_15930_)
  );
  AND2_X1 _51200_ (
    .A1(\cpuregs[9] [12]),
    .A2(_12560_),
    .ZN(_15931_)
  );
  INV_X1 _51201_ (
    .A(_15931_),
    .ZN(_15932_)
  );
  AND2_X1 _51202_ (
    .A1(_15930_),
    .A2(_15932_),
    .ZN(_15933_)
  );
  INV_X1 _51203_ (
    .A(_15933_),
    .ZN(_01097_)
  );
  AND2_X1 _51204_ (
    .A1(_12559_),
    .A2(_13063_),
    .ZN(_15934_)
  );
  INV_X1 _51205_ (
    .A(_15934_),
    .ZN(_15935_)
  );
  AND2_X1 _51206_ (
    .A1(\cpuregs[9] [13]),
    .A2(_12560_),
    .ZN(_15936_)
  );
  INV_X1 _51207_ (
    .A(_15936_),
    .ZN(_15937_)
  );
  AND2_X1 _51208_ (
    .A1(_15935_),
    .A2(_15937_),
    .ZN(_15938_)
  );
  INV_X1 _51209_ (
    .A(_15938_),
    .ZN(_01098_)
  );
  AND2_X1 _51210_ (
    .A1(_12559_),
    .A2(_13078_),
    .ZN(_15939_)
  );
  INV_X1 _51211_ (
    .A(_15939_),
    .ZN(_15940_)
  );
  AND2_X1 _51212_ (
    .A1(\cpuregs[9] [14]),
    .A2(_12560_),
    .ZN(_15941_)
  );
  INV_X1 _51213_ (
    .A(_15941_),
    .ZN(_15942_)
  );
  AND2_X1 _51214_ (
    .A1(_15940_),
    .A2(_15942_),
    .ZN(_15943_)
  );
  INV_X1 _51215_ (
    .A(_15943_),
    .ZN(_01099_)
  );
  AND2_X1 _51216_ (
    .A1(_12559_),
    .A2(_13093_),
    .ZN(_15944_)
  );
  INV_X1 _51217_ (
    .A(_15944_),
    .ZN(_15945_)
  );
  AND2_X1 _51218_ (
    .A1(\cpuregs[9] [15]),
    .A2(_12560_),
    .ZN(_15946_)
  );
  INV_X1 _51219_ (
    .A(_15946_),
    .ZN(_15947_)
  );
  AND2_X1 _51220_ (
    .A1(_15945_),
    .A2(_15947_),
    .ZN(_15948_)
  );
  INV_X1 _51221_ (
    .A(_15948_),
    .ZN(_01100_)
  );
  AND2_X1 _51222_ (
    .A1(\cpuregs[9] [16]),
    .A2(_12560_),
    .ZN(_15949_)
  );
  INV_X1 _51223_ (
    .A(_15949_),
    .ZN(_15950_)
  );
  AND2_X1 _51224_ (
    .A1(_12559_),
    .A2(_13108_),
    .ZN(_15951_)
  );
  INV_X1 _51225_ (
    .A(_15951_),
    .ZN(_15952_)
  );
  AND2_X1 _51226_ (
    .A1(_15950_),
    .A2(_15952_),
    .ZN(_15953_)
  );
  INV_X1 _51227_ (
    .A(_15953_),
    .ZN(_01101_)
  );
  AND2_X1 _51228_ (
    .A1(_12559_),
    .A2(_13123_),
    .ZN(_15954_)
  );
  INV_X1 _51229_ (
    .A(_15954_),
    .ZN(_15955_)
  );
  AND2_X1 _51230_ (
    .A1(\cpuregs[9] [17]),
    .A2(_12560_),
    .ZN(_15956_)
  );
  INV_X1 _51231_ (
    .A(_15956_),
    .ZN(_15957_)
  );
  AND2_X1 _51232_ (
    .A1(_15955_),
    .A2(_15957_),
    .ZN(_15958_)
  );
  INV_X1 _51233_ (
    .A(_15958_),
    .ZN(_01102_)
  );
  AND2_X1 _51234_ (
    .A1(_12559_),
    .A2(_13139_),
    .ZN(_15959_)
  );
  INV_X1 _51235_ (
    .A(_15959_),
    .ZN(_15960_)
  );
  AND2_X1 _51236_ (
    .A1(\cpuregs[9] [18]),
    .A2(_12560_),
    .ZN(_15961_)
  );
  INV_X1 _51237_ (
    .A(_15961_),
    .ZN(_15962_)
  );
  AND2_X1 _51238_ (
    .A1(_15960_),
    .A2(_15962_),
    .ZN(_15963_)
  );
  INV_X1 _51239_ (
    .A(_15963_),
    .ZN(_01103_)
  );
  AND2_X1 _51240_ (
    .A1(_12559_),
    .A2(_13154_),
    .ZN(_15964_)
  );
  INV_X1 _51241_ (
    .A(_15964_),
    .ZN(_15965_)
  );
  AND2_X1 _51242_ (
    .A1(\cpuregs[9] [19]),
    .A2(_12560_),
    .ZN(_15966_)
  );
  INV_X1 _51243_ (
    .A(_15966_),
    .ZN(_15967_)
  );
  AND2_X1 _51244_ (
    .A1(_15965_),
    .A2(_15967_),
    .ZN(_15968_)
  );
  INV_X1 _51245_ (
    .A(_15968_),
    .ZN(_01104_)
  );
  AND2_X1 _51246_ (
    .A1(_12559_),
    .A2(_13169_),
    .ZN(_15969_)
  );
  INV_X1 _51247_ (
    .A(_15969_),
    .ZN(_15970_)
  );
  AND2_X1 _51248_ (
    .A1(\cpuregs[9] [20]),
    .A2(_12560_),
    .ZN(_15971_)
  );
  INV_X1 _51249_ (
    .A(_15971_),
    .ZN(_15972_)
  );
  AND2_X1 _51250_ (
    .A1(_15970_),
    .A2(_15972_),
    .ZN(_15973_)
  );
  INV_X1 _51251_ (
    .A(_15973_),
    .ZN(_01105_)
  );
  AND2_X1 _51252_ (
    .A1(_12559_),
    .A2(_13184_),
    .ZN(_15974_)
  );
  INV_X1 _51253_ (
    .A(_15974_),
    .ZN(_15975_)
  );
  AND2_X1 _51254_ (
    .A1(\cpuregs[9] [21]),
    .A2(_12560_),
    .ZN(_15976_)
  );
  INV_X1 _51255_ (
    .A(_15976_),
    .ZN(_15977_)
  );
  AND2_X1 _51256_ (
    .A1(_15975_),
    .A2(_15977_),
    .ZN(_15978_)
  );
  INV_X1 _51257_ (
    .A(_15978_),
    .ZN(_01106_)
  );
  AND2_X1 _51258_ (
    .A1(_12559_),
    .A2(_13199_),
    .ZN(_15979_)
  );
  INV_X1 _51259_ (
    .A(_15979_),
    .ZN(_15980_)
  );
  AND2_X1 _51260_ (
    .A1(\cpuregs[9] [22]),
    .A2(_12560_),
    .ZN(_15981_)
  );
  INV_X1 _51261_ (
    .A(_15981_),
    .ZN(_15982_)
  );
  AND2_X1 _51262_ (
    .A1(_15980_),
    .A2(_15982_),
    .ZN(_15983_)
  );
  INV_X1 _51263_ (
    .A(_15983_),
    .ZN(_01107_)
  );
  AND2_X1 _51264_ (
    .A1(_12559_),
    .A2(_13214_),
    .ZN(_15984_)
  );
  INV_X1 _51265_ (
    .A(_15984_),
    .ZN(_15985_)
  );
  AND2_X1 _51266_ (
    .A1(\cpuregs[9] [23]),
    .A2(_12560_),
    .ZN(_15986_)
  );
  INV_X1 _51267_ (
    .A(_15986_),
    .ZN(_15987_)
  );
  AND2_X1 _51268_ (
    .A1(_15985_),
    .A2(_15987_),
    .ZN(_15988_)
  );
  INV_X1 _51269_ (
    .A(_15988_),
    .ZN(_01108_)
  );
  AND2_X1 _51270_ (
    .A1(_12559_),
    .A2(_13229_),
    .ZN(_15989_)
  );
  INV_X1 _51271_ (
    .A(_15989_),
    .ZN(_15990_)
  );
  AND2_X1 _51272_ (
    .A1(\cpuregs[9] [24]),
    .A2(_12560_),
    .ZN(_15991_)
  );
  INV_X1 _51273_ (
    .A(_15991_),
    .ZN(_15992_)
  );
  AND2_X1 _51274_ (
    .A1(_15990_),
    .A2(_15992_),
    .ZN(_15993_)
  );
  INV_X1 _51275_ (
    .A(_15993_),
    .ZN(_01109_)
  );
  AND2_X1 _51276_ (
    .A1(_12559_),
    .A2(_13244_),
    .ZN(_15994_)
  );
  INV_X1 _51277_ (
    .A(_15994_),
    .ZN(_15995_)
  );
  AND2_X1 _51278_ (
    .A1(\cpuregs[9] [25]),
    .A2(_12560_),
    .ZN(_15996_)
  );
  INV_X1 _51279_ (
    .A(_15996_),
    .ZN(_15997_)
  );
  AND2_X1 _51280_ (
    .A1(_15995_),
    .A2(_15997_),
    .ZN(_15998_)
  );
  INV_X1 _51281_ (
    .A(_15998_),
    .ZN(_01110_)
  );
  AND2_X1 _51282_ (
    .A1(_12559_),
    .A2(_13259_),
    .ZN(_15999_)
  );
  INV_X1 _51283_ (
    .A(_15999_),
    .ZN(_16000_)
  );
  AND2_X1 _51284_ (
    .A1(\cpuregs[9] [26]),
    .A2(_12560_),
    .ZN(_16001_)
  );
  INV_X1 _51285_ (
    .A(_16001_),
    .ZN(_16002_)
  );
  AND2_X1 _51286_ (
    .A1(_16000_),
    .A2(_16002_),
    .ZN(_16003_)
  );
  INV_X1 _51287_ (
    .A(_16003_),
    .ZN(_01111_)
  );
  AND2_X1 _51288_ (
    .A1(_12559_),
    .A2(_13274_),
    .ZN(_16004_)
  );
  INV_X1 _51289_ (
    .A(_16004_),
    .ZN(_16005_)
  );
  AND2_X1 _51290_ (
    .A1(\cpuregs[9] [27]),
    .A2(_12560_),
    .ZN(_16006_)
  );
  INV_X1 _51291_ (
    .A(_16006_),
    .ZN(_16007_)
  );
  AND2_X1 _51292_ (
    .A1(_16005_),
    .A2(_16007_),
    .ZN(_16008_)
  );
  INV_X1 _51293_ (
    .A(_16008_),
    .ZN(_01112_)
  );
  AND2_X1 _51294_ (
    .A1(_12559_),
    .A2(_13289_),
    .ZN(_16009_)
  );
  INV_X1 _51295_ (
    .A(_16009_),
    .ZN(_16010_)
  );
  AND2_X1 _51296_ (
    .A1(\cpuregs[9] [28]),
    .A2(_12560_),
    .ZN(_16011_)
  );
  INV_X1 _51297_ (
    .A(_16011_),
    .ZN(_16012_)
  );
  AND2_X1 _51298_ (
    .A1(_16010_),
    .A2(_16012_),
    .ZN(_16013_)
  );
  INV_X1 _51299_ (
    .A(_16013_),
    .ZN(_01113_)
  );
  AND2_X1 _51300_ (
    .A1(_12559_),
    .A2(_13304_),
    .ZN(_16014_)
  );
  INV_X1 _51301_ (
    .A(_16014_),
    .ZN(_16015_)
  );
  AND2_X1 _51302_ (
    .A1(\cpuregs[9] [29]),
    .A2(_12560_),
    .ZN(_16016_)
  );
  INV_X1 _51303_ (
    .A(_16016_),
    .ZN(_16017_)
  );
  AND2_X1 _51304_ (
    .A1(_16015_),
    .A2(_16017_),
    .ZN(_16018_)
  );
  INV_X1 _51305_ (
    .A(_16018_),
    .ZN(_01114_)
  );
  AND2_X1 _51306_ (
    .A1(_12559_),
    .A2(_13319_),
    .ZN(_16019_)
  );
  INV_X1 _51307_ (
    .A(_16019_),
    .ZN(_16020_)
  );
  AND2_X1 _51308_ (
    .A1(\cpuregs[9] [30]),
    .A2(_12560_),
    .ZN(_16021_)
  );
  INV_X1 _51309_ (
    .A(_16021_),
    .ZN(_16022_)
  );
  AND2_X1 _51310_ (
    .A1(_16020_),
    .A2(_16022_),
    .ZN(_16023_)
  );
  INV_X1 _51311_ (
    .A(_16023_),
    .ZN(_01115_)
  );
  AND2_X1 _51312_ (
    .A1(_12634_),
    .A2(_12874_),
    .ZN(_16024_)
  );
  INV_X1 _51313_ (
    .A(_16024_),
    .ZN(_16025_)
  );
  AND2_X1 _51314_ (
    .A1(\cpuregs[8] [0]),
    .A2(_12635_),
    .ZN(_16026_)
  );
  INV_X1 _51315_ (
    .A(_16026_),
    .ZN(_16027_)
  );
  AND2_X1 _51316_ (
    .A1(_16025_),
    .A2(_16027_),
    .ZN(_16028_)
  );
  INV_X1 _51317_ (
    .A(_16028_),
    .ZN(_01116_)
  );
  AND2_X1 _51318_ (
    .A1(_12634_),
    .A2(_12886_),
    .ZN(_16029_)
  );
  INV_X1 _51319_ (
    .A(_16029_),
    .ZN(_16030_)
  );
  AND2_X1 _51320_ (
    .A1(\cpuregs[8] [1]),
    .A2(_12635_),
    .ZN(_16031_)
  );
  INV_X1 _51321_ (
    .A(_16031_),
    .ZN(_16032_)
  );
  AND2_X1 _51322_ (
    .A1(_16030_),
    .A2(_16032_),
    .ZN(_16033_)
  );
  INV_X1 _51323_ (
    .A(_16033_),
    .ZN(_01117_)
  );
  AND2_X1 _51324_ (
    .A1(_12634_),
    .A2(_12900_),
    .ZN(_16034_)
  );
  INV_X1 _51325_ (
    .A(_16034_),
    .ZN(_16035_)
  );
  AND2_X1 _51326_ (
    .A1(\cpuregs[8] [2]),
    .A2(_12635_),
    .ZN(_16036_)
  );
  INV_X1 _51327_ (
    .A(_16036_),
    .ZN(_16037_)
  );
  AND2_X1 _51328_ (
    .A1(_16035_),
    .A2(_16037_),
    .ZN(_16038_)
  );
  INV_X1 _51329_ (
    .A(_16038_),
    .ZN(_01118_)
  );
  AND2_X1 _51330_ (
    .A1(_12634_),
    .A2(_12913_),
    .ZN(_16039_)
  );
  INV_X1 _51331_ (
    .A(_16039_),
    .ZN(_16040_)
  );
  AND2_X1 _51332_ (
    .A1(\cpuregs[8] [3]),
    .A2(_12635_),
    .ZN(_16041_)
  );
  INV_X1 _51333_ (
    .A(_16041_),
    .ZN(_16042_)
  );
  AND2_X1 _51334_ (
    .A1(_16040_),
    .A2(_16042_),
    .ZN(_16043_)
  );
  INV_X1 _51335_ (
    .A(_16043_),
    .ZN(_01119_)
  );
  AND2_X1 _51336_ (
    .A1(\cpuregs[8] [4]),
    .A2(_12635_),
    .ZN(_16044_)
  );
  INV_X1 _51337_ (
    .A(_16044_),
    .ZN(_16045_)
  );
  AND2_X1 _51338_ (
    .A1(_12634_),
    .A2(_12928_),
    .ZN(_16046_)
  );
  INV_X1 _51339_ (
    .A(_16046_),
    .ZN(_16047_)
  );
  AND2_X1 _51340_ (
    .A1(_16045_),
    .A2(_16047_),
    .ZN(_16048_)
  );
  INV_X1 _51341_ (
    .A(_16048_),
    .ZN(_01120_)
  );
  AND2_X1 _51342_ (
    .A1(_12634_),
    .A2(_12943_),
    .ZN(_16049_)
  );
  INV_X1 _51343_ (
    .A(_16049_),
    .ZN(_16050_)
  );
  AND2_X1 _51344_ (
    .A1(\cpuregs[8] [5]),
    .A2(_12635_),
    .ZN(_16051_)
  );
  INV_X1 _51345_ (
    .A(_16051_),
    .ZN(_16052_)
  );
  AND2_X1 _51346_ (
    .A1(_16050_),
    .A2(_16052_),
    .ZN(_16053_)
  );
  INV_X1 _51347_ (
    .A(_16053_),
    .ZN(_01121_)
  );
  AND2_X1 _51348_ (
    .A1(_12634_),
    .A2(_12958_),
    .ZN(_16054_)
  );
  INV_X1 _51349_ (
    .A(_16054_),
    .ZN(_16055_)
  );
  AND2_X1 _51350_ (
    .A1(\cpuregs[8] [6]),
    .A2(_12635_),
    .ZN(_16056_)
  );
  INV_X1 _51351_ (
    .A(_16056_),
    .ZN(_16057_)
  );
  AND2_X1 _51352_ (
    .A1(_16055_),
    .A2(_16057_),
    .ZN(_16058_)
  );
  INV_X1 _51353_ (
    .A(_16058_),
    .ZN(_01122_)
  );
  AND2_X1 _51354_ (
    .A1(_12634_),
    .A2(_12973_),
    .ZN(_16059_)
  );
  INV_X1 _51355_ (
    .A(_16059_),
    .ZN(_16060_)
  );
  AND2_X1 _51356_ (
    .A1(\cpuregs[8] [7]),
    .A2(_12635_),
    .ZN(_16061_)
  );
  INV_X1 _51357_ (
    .A(_16061_),
    .ZN(_16062_)
  );
  AND2_X1 _51358_ (
    .A1(_16060_),
    .A2(_16062_),
    .ZN(_16063_)
  );
  INV_X1 _51359_ (
    .A(_16063_),
    .ZN(_01123_)
  );
  AND2_X1 _51360_ (
    .A1(_12634_),
    .A2(_12988_),
    .ZN(_16064_)
  );
  INV_X1 _51361_ (
    .A(_16064_),
    .ZN(_16065_)
  );
  AND2_X1 _51362_ (
    .A1(\cpuregs[8] [8]),
    .A2(_12635_),
    .ZN(_16066_)
  );
  INV_X1 _51363_ (
    .A(_16066_),
    .ZN(_16067_)
  );
  AND2_X1 _51364_ (
    .A1(_16065_),
    .A2(_16067_),
    .ZN(_16068_)
  );
  INV_X1 _51365_ (
    .A(_16068_),
    .ZN(_01124_)
  );
  AND2_X1 _51366_ (
    .A1(_12634_),
    .A2(_13003_),
    .ZN(_16069_)
  );
  INV_X1 _51367_ (
    .A(_16069_),
    .ZN(_16070_)
  );
  AND2_X1 _51368_ (
    .A1(\cpuregs[8] [9]),
    .A2(_12635_),
    .ZN(_16071_)
  );
  INV_X1 _51369_ (
    .A(_16071_),
    .ZN(_16072_)
  );
  AND2_X1 _51370_ (
    .A1(_16070_),
    .A2(_16072_),
    .ZN(_16073_)
  );
  INV_X1 _51371_ (
    .A(_16073_),
    .ZN(_01125_)
  );
  AND2_X1 _51372_ (
    .A1(_12634_),
    .A2(_13018_),
    .ZN(_16074_)
  );
  INV_X1 _51373_ (
    .A(_16074_),
    .ZN(_16075_)
  );
  AND2_X1 _51374_ (
    .A1(\cpuregs[8] [10]),
    .A2(_12635_),
    .ZN(_16076_)
  );
  INV_X1 _51375_ (
    .A(_16076_),
    .ZN(_16077_)
  );
  AND2_X1 _51376_ (
    .A1(_16075_),
    .A2(_16077_),
    .ZN(_16078_)
  );
  INV_X1 _51377_ (
    .A(_16078_),
    .ZN(_01126_)
  );
  AND2_X1 _51378_ (
    .A1(_12634_),
    .A2(_13033_),
    .ZN(_16079_)
  );
  INV_X1 _51379_ (
    .A(_16079_),
    .ZN(_16080_)
  );
  AND2_X1 _51380_ (
    .A1(\cpuregs[8] [11]),
    .A2(_12635_),
    .ZN(_16081_)
  );
  INV_X1 _51381_ (
    .A(_16081_),
    .ZN(_16082_)
  );
  AND2_X1 _51382_ (
    .A1(_16080_),
    .A2(_16082_),
    .ZN(_16083_)
  );
  INV_X1 _51383_ (
    .A(_16083_),
    .ZN(_01127_)
  );
  AND2_X1 _51384_ (
    .A1(_12634_),
    .A2(_13048_),
    .ZN(_16084_)
  );
  INV_X1 _51385_ (
    .A(_16084_),
    .ZN(_16085_)
  );
  AND2_X1 _51386_ (
    .A1(\cpuregs[8] [12]),
    .A2(_12635_),
    .ZN(_16086_)
  );
  INV_X1 _51387_ (
    .A(_16086_),
    .ZN(_16087_)
  );
  AND2_X1 _51388_ (
    .A1(_16085_),
    .A2(_16087_),
    .ZN(_16088_)
  );
  INV_X1 _51389_ (
    .A(_16088_),
    .ZN(_01128_)
  );
  AND2_X1 _51390_ (
    .A1(_12634_),
    .A2(_13063_),
    .ZN(_16089_)
  );
  INV_X1 _51391_ (
    .A(_16089_),
    .ZN(_16090_)
  );
  AND2_X1 _51392_ (
    .A1(\cpuregs[8] [13]),
    .A2(_12635_),
    .ZN(_16091_)
  );
  INV_X1 _51393_ (
    .A(_16091_),
    .ZN(_16092_)
  );
  AND2_X1 _51394_ (
    .A1(_16090_),
    .A2(_16092_),
    .ZN(_16093_)
  );
  INV_X1 _51395_ (
    .A(_16093_),
    .ZN(_01129_)
  );
  AND2_X1 _51396_ (
    .A1(_12634_),
    .A2(_13078_),
    .ZN(_16094_)
  );
  INV_X1 _51397_ (
    .A(_16094_),
    .ZN(_16095_)
  );
  AND2_X1 _51398_ (
    .A1(\cpuregs[8] [14]),
    .A2(_12635_),
    .ZN(_16096_)
  );
  INV_X1 _51399_ (
    .A(_16096_),
    .ZN(_16097_)
  );
  AND2_X1 _51400_ (
    .A1(_16095_),
    .A2(_16097_),
    .ZN(_16098_)
  );
  INV_X1 _51401_ (
    .A(_16098_),
    .ZN(_01130_)
  );
  AND2_X1 _51402_ (
    .A1(_12634_),
    .A2(_13093_),
    .ZN(_16099_)
  );
  INV_X1 _51403_ (
    .A(_16099_),
    .ZN(_16100_)
  );
  AND2_X1 _51404_ (
    .A1(\cpuregs[8] [15]),
    .A2(_12635_),
    .ZN(_16101_)
  );
  INV_X1 _51405_ (
    .A(_16101_),
    .ZN(_16102_)
  );
  AND2_X1 _51406_ (
    .A1(_16100_),
    .A2(_16102_),
    .ZN(_16103_)
  );
  INV_X1 _51407_ (
    .A(_16103_),
    .ZN(_01131_)
  );
  AND2_X1 _51408_ (
    .A1(_12634_),
    .A2(_13108_),
    .ZN(_16104_)
  );
  INV_X1 _51409_ (
    .A(_16104_),
    .ZN(_16105_)
  );
  AND2_X1 _51410_ (
    .A1(\cpuregs[8] [16]),
    .A2(_12635_),
    .ZN(_16106_)
  );
  INV_X1 _51411_ (
    .A(_16106_),
    .ZN(_16107_)
  );
  AND2_X1 _51412_ (
    .A1(_16105_),
    .A2(_16107_),
    .ZN(_16108_)
  );
  INV_X1 _51413_ (
    .A(_16108_),
    .ZN(_01132_)
  );
  AND2_X1 _51414_ (
    .A1(\cpuregs[8] [17]),
    .A2(_12635_),
    .ZN(_16109_)
  );
  INV_X1 _51415_ (
    .A(_16109_),
    .ZN(_16110_)
  );
  AND2_X1 _51416_ (
    .A1(_12634_),
    .A2(_13123_),
    .ZN(_16111_)
  );
  INV_X1 _51417_ (
    .A(_16111_),
    .ZN(_16112_)
  );
  AND2_X1 _51418_ (
    .A1(_16110_),
    .A2(_16112_),
    .ZN(_16113_)
  );
  INV_X1 _51419_ (
    .A(_16113_),
    .ZN(_01133_)
  );
  AND2_X1 _51420_ (
    .A1(\cpuregs[8] [18]),
    .A2(_12635_),
    .ZN(_16114_)
  );
  INV_X1 _51421_ (
    .A(_16114_),
    .ZN(_16115_)
  );
  AND2_X1 _51422_ (
    .A1(_12634_),
    .A2(_13139_),
    .ZN(_16116_)
  );
  INV_X1 _51423_ (
    .A(_16116_),
    .ZN(_16117_)
  );
  AND2_X1 _51424_ (
    .A1(_16115_),
    .A2(_16117_),
    .ZN(_16118_)
  );
  INV_X1 _51425_ (
    .A(_16118_),
    .ZN(_01134_)
  );
  AND2_X1 _51426_ (
    .A1(\cpuregs[8] [19]),
    .A2(_12635_),
    .ZN(_16119_)
  );
  INV_X1 _51427_ (
    .A(_16119_),
    .ZN(_16120_)
  );
  AND2_X1 _51428_ (
    .A1(_12634_),
    .A2(_13154_),
    .ZN(_16121_)
  );
  INV_X1 _51429_ (
    .A(_16121_),
    .ZN(_16122_)
  );
  AND2_X1 _51430_ (
    .A1(_16120_),
    .A2(_16122_),
    .ZN(_16123_)
  );
  INV_X1 _51431_ (
    .A(_16123_),
    .ZN(_01135_)
  );
  AND2_X1 _51432_ (
    .A1(\cpuregs[8] [20]),
    .A2(_12635_),
    .ZN(_16124_)
  );
  INV_X1 _51433_ (
    .A(_16124_),
    .ZN(_16125_)
  );
  AND2_X1 _51434_ (
    .A1(_12634_),
    .A2(_13169_),
    .ZN(_16126_)
  );
  INV_X1 _51435_ (
    .A(_16126_),
    .ZN(_16127_)
  );
  AND2_X1 _51436_ (
    .A1(_16125_),
    .A2(_16127_),
    .ZN(_16128_)
  );
  INV_X1 _51437_ (
    .A(_16128_),
    .ZN(_01136_)
  );
  AND2_X1 _51438_ (
    .A1(\cpuregs[8] [21]),
    .A2(_12635_),
    .ZN(_16129_)
  );
  INV_X1 _51439_ (
    .A(_16129_),
    .ZN(_16130_)
  );
  AND2_X1 _51440_ (
    .A1(_12634_),
    .A2(_13184_),
    .ZN(_16131_)
  );
  INV_X1 _51441_ (
    .A(_16131_),
    .ZN(_16132_)
  );
  AND2_X1 _51442_ (
    .A1(_16130_),
    .A2(_16132_),
    .ZN(_16133_)
  );
  INV_X1 _51443_ (
    .A(_16133_),
    .ZN(_01137_)
  );
  AND2_X1 _51444_ (
    .A1(\cpuregs[8] [22]),
    .A2(_12635_),
    .ZN(_16134_)
  );
  INV_X1 _51445_ (
    .A(_16134_),
    .ZN(_16135_)
  );
  AND2_X1 _51446_ (
    .A1(_12634_),
    .A2(_13199_),
    .ZN(_16136_)
  );
  INV_X1 _51447_ (
    .A(_16136_),
    .ZN(_16137_)
  );
  AND2_X1 _51448_ (
    .A1(_16135_),
    .A2(_16137_),
    .ZN(_16138_)
  );
  INV_X1 _51449_ (
    .A(_16138_),
    .ZN(_01138_)
  );
  AND2_X1 _51450_ (
    .A1(\cpuregs[8] [23]),
    .A2(_12635_),
    .ZN(_16139_)
  );
  INV_X1 _51451_ (
    .A(_16139_),
    .ZN(_16140_)
  );
  AND2_X1 _51452_ (
    .A1(_12634_),
    .A2(_13214_),
    .ZN(_16141_)
  );
  INV_X1 _51453_ (
    .A(_16141_),
    .ZN(_16142_)
  );
  AND2_X1 _51454_ (
    .A1(_16140_),
    .A2(_16142_),
    .ZN(_16143_)
  );
  INV_X1 _51455_ (
    .A(_16143_),
    .ZN(_01139_)
  );
  AND2_X1 _51456_ (
    .A1(\cpuregs[8] [24]),
    .A2(_12635_),
    .ZN(_16144_)
  );
  INV_X1 _51457_ (
    .A(_16144_),
    .ZN(_16145_)
  );
  AND2_X1 _51458_ (
    .A1(_12634_),
    .A2(_13229_),
    .ZN(_16146_)
  );
  INV_X1 _51459_ (
    .A(_16146_),
    .ZN(_16147_)
  );
  AND2_X1 _51460_ (
    .A1(_16145_),
    .A2(_16147_),
    .ZN(_16148_)
  );
  INV_X1 _51461_ (
    .A(_16148_),
    .ZN(_01140_)
  );
  AND2_X1 _51462_ (
    .A1(\cpuregs[8] [25]),
    .A2(_12635_),
    .ZN(_16149_)
  );
  INV_X1 _51463_ (
    .A(_16149_),
    .ZN(_16150_)
  );
  AND2_X1 _51464_ (
    .A1(_12634_),
    .A2(_13244_),
    .ZN(_16151_)
  );
  INV_X1 _51465_ (
    .A(_16151_),
    .ZN(_16152_)
  );
  AND2_X1 _51466_ (
    .A1(_16150_),
    .A2(_16152_),
    .ZN(_16153_)
  );
  INV_X1 _51467_ (
    .A(_16153_),
    .ZN(_01141_)
  );
  AND2_X1 _51468_ (
    .A1(\cpuregs[8] [26]),
    .A2(_12635_),
    .ZN(_16154_)
  );
  INV_X1 _51469_ (
    .A(_16154_),
    .ZN(_16155_)
  );
  AND2_X1 _51470_ (
    .A1(_12634_),
    .A2(_13259_),
    .ZN(_16156_)
  );
  INV_X1 _51471_ (
    .A(_16156_),
    .ZN(_16157_)
  );
  AND2_X1 _51472_ (
    .A1(_16155_),
    .A2(_16157_),
    .ZN(_16158_)
  );
  INV_X1 _51473_ (
    .A(_16158_),
    .ZN(_01142_)
  );
  AND2_X1 _51474_ (
    .A1(\cpuregs[8] [27]),
    .A2(_12635_),
    .ZN(_16159_)
  );
  INV_X1 _51475_ (
    .A(_16159_),
    .ZN(_16160_)
  );
  AND2_X1 _51476_ (
    .A1(_12634_),
    .A2(_13274_),
    .ZN(_16161_)
  );
  INV_X1 _51477_ (
    .A(_16161_),
    .ZN(_16162_)
  );
  AND2_X1 _51478_ (
    .A1(_16160_),
    .A2(_16162_),
    .ZN(_16163_)
  );
  INV_X1 _51479_ (
    .A(_16163_),
    .ZN(_01143_)
  );
  AND2_X1 _51480_ (
    .A1(\cpuregs[8] [28]),
    .A2(_12635_),
    .ZN(_16164_)
  );
  INV_X1 _51481_ (
    .A(_16164_),
    .ZN(_16165_)
  );
  AND2_X1 _51482_ (
    .A1(_12634_),
    .A2(_13289_),
    .ZN(_16166_)
  );
  INV_X1 _51483_ (
    .A(_16166_),
    .ZN(_16167_)
  );
  AND2_X1 _51484_ (
    .A1(_16165_),
    .A2(_16167_),
    .ZN(_16168_)
  );
  INV_X1 _51485_ (
    .A(_16168_),
    .ZN(_01144_)
  );
  AND2_X1 _51486_ (
    .A1(\cpuregs[8] [29]),
    .A2(_12635_),
    .ZN(_16169_)
  );
  INV_X1 _51487_ (
    .A(_16169_),
    .ZN(_16170_)
  );
  AND2_X1 _51488_ (
    .A1(_12634_),
    .A2(_13304_),
    .ZN(_16171_)
  );
  INV_X1 _51489_ (
    .A(_16171_),
    .ZN(_16172_)
  );
  AND2_X1 _51490_ (
    .A1(_16170_),
    .A2(_16172_),
    .ZN(_16173_)
  );
  INV_X1 _51491_ (
    .A(_16173_),
    .ZN(_01145_)
  );
  AND2_X1 _51492_ (
    .A1(\cpuregs[8] [30]),
    .A2(_12635_),
    .ZN(_16174_)
  );
  INV_X1 _51493_ (
    .A(_16174_),
    .ZN(_16175_)
  );
  AND2_X1 _51494_ (
    .A1(_12634_),
    .A2(_13319_),
    .ZN(_16176_)
  );
  INV_X1 _51495_ (
    .A(_16176_),
    .ZN(_16177_)
  );
  AND2_X1 _51496_ (
    .A1(_16175_),
    .A2(_16177_),
    .ZN(_16178_)
  );
  INV_X1 _51497_ (
    .A(_16178_),
    .ZN(_01146_)
  );
  AND2_X1 _51498_ (
    .A1(_12665_),
    .A2(_12874_),
    .ZN(_16179_)
  );
  INV_X1 _51499_ (
    .A(_16179_),
    .ZN(_16180_)
  );
  AND2_X1 _51500_ (
    .A1(\cpuregs[5] [0]),
    .A2(_12666_),
    .ZN(_16181_)
  );
  INV_X1 _51501_ (
    .A(_16181_),
    .ZN(_16182_)
  );
  AND2_X1 _51502_ (
    .A1(_16180_),
    .A2(_16182_),
    .ZN(_16183_)
  );
  INV_X1 _51503_ (
    .A(_16183_),
    .ZN(_01147_)
  );
  AND2_X1 _51504_ (
    .A1(_12665_),
    .A2(_12886_),
    .ZN(_16184_)
  );
  INV_X1 _51505_ (
    .A(_16184_),
    .ZN(_16185_)
  );
  AND2_X1 _51506_ (
    .A1(\cpuregs[5] [1]),
    .A2(_12666_),
    .ZN(_16186_)
  );
  INV_X1 _51507_ (
    .A(_16186_),
    .ZN(_16187_)
  );
  AND2_X1 _51508_ (
    .A1(_16185_),
    .A2(_16187_),
    .ZN(_16188_)
  );
  INV_X1 _51509_ (
    .A(_16188_),
    .ZN(_01148_)
  );
  AND2_X1 _51510_ (
    .A1(\cpuregs[5] [2]),
    .A2(_12666_),
    .ZN(_16189_)
  );
  INV_X1 _51511_ (
    .A(_16189_),
    .ZN(_16190_)
  );
  AND2_X1 _51512_ (
    .A1(_12665_),
    .A2(_12900_),
    .ZN(_16191_)
  );
  INV_X1 _51513_ (
    .A(_16191_),
    .ZN(_16192_)
  );
  AND2_X1 _51514_ (
    .A1(_16190_),
    .A2(_16192_),
    .ZN(_16193_)
  );
  INV_X1 _51515_ (
    .A(_16193_),
    .ZN(_01149_)
  );
  AND2_X1 _51516_ (
    .A1(_12665_),
    .A2(_12913_),
    .ZN(_16194_)
  );
  INV_X1 _51517_ (
    .A(_16194_),
    .ZN(_16195_)
  );
  AND2_X1 _51518_ (
    .A1(\cpuregs[5] [3]),
    .A2(_12666_),
    .ZN(_16196_)
  );
  INV_X1 _51519_ (
    .A(_16196_),
    .ZN(_16197_)
  );
  AND2_X1 _51520_ (
    .A1(_16195_),
    .A2(_16197_),
    .ZN(_16198_)
  );
  INV_X1 _51521_ (
    .A(_16198_),
    .ZN(_01150_)
  );
  AND2_X1 _51522_ (
    .A1(\cpuregs[5] [4]),
    .A2(_12666_),
    .ZN(_16199_)
  );
  INV_X1 _51523_ (
    .A(_16199_),
    .ZN(_16200_)
  );
  AND2_X1 _51524_ (
    .A1(_12665_),
    .A2(_12928_),
    .ZN(_16201_)
  );
  INV_X1 _51525_ (
    .A(_16201_),
    .ZN(_16202_)
  );
  AND2_X1 _51526_ (
    .A1(_16200_),
    .A2(_16202_),
    .ZN(_16203_)
  );
  INV_X1 _51527_ (
    .A(_16203_),
    .ZN(_01151_)
  );
  AND2_X1 _51528_ (
    .A1(_12665_),
    .A2(_12943_),
    .ZN(_16204_)
  );
  INV_X1 _51529_ (
    .A(_16204_),
    .ZN(_16205_)
  );
  AND2_X1 _51530_ (
    .A1(\cpuregs[5] [5]),
    .A2(_12666_),
    .ZN(_16206_)
  );
  INV_X1 _51531_ (
    .A(_16206_),
    .ZN(_16207_)
  );
  AND2_X1 _51532_ (
    .A1(_16205_),
    .A2(_16207_),
    .ZN(_16208_)
  );
  INV_X1 _51533_ (
    .A(_16208_),
    .ZN(_01152_)
  );
  AND2_X1 _51534_ (
    .A1(_12665_),
    .A2(_12958_),
    .ZN(_16209_)
  );
  INV_X1 _51535_ (
    .A(_16209_),
    .ZN(_16210_)
  );
  AND2_X1 _51536_ (
    .A1(\cpuregs[5] [6]),
    .A2(_12666_),
    .ZN(_16211_)
  );
  INV_X1 _51537_ (
    .A(_16211_),
    .ZN(_16212_)
  );
  AND2_X1 _51538_ (
    .A1(_16210_),
    .A2(_16212_),
    .ZN(_16213_)
  );
  INV_X1 _51539_ (
    .A(_16213_),
    .ZN(_01153_)
  );
  AND2_X1 _51540_ (
    .A1(_12665_),
    .A2(_12973_),
    .ZN(_16214_)
  );
  INV_X1 _51541_ (
    .A(_16214_),
    .ZN(_16215_)
  );
  AND2_X1 _51542_ (
    .A1(\cpuregs[5] [7]),
    .A2(_12666_),
    .ZN(_16216_)
  );
  INV_X1 _51543_ (
    .A(_16216_),
    .ZN(_16217_)
  );
  AND2_X1 _51544_ (
    .A1(_16215_),
    .A2(_16217_),
    .ZN(_16218_)
  );
  INV_X1 _51545_ (
    .A(_16218_),
    .ZN(_01154_)
  );
  AND2_X1 _51546_ (
    .A1(_12665_),
    .A2(_12988_),
    .ZN(_16219_)
  );
  INV_X1 _51547_ (
    .A(_16219_),
    .ZN(_16220_)
  );
  AND2_X1 _51548_ (
    .A1(\cpuregs[5] [8]),
    .A2(_12666_),
    .ZN(_16221_)
  );
  INV_X1 _51549_ (
    .A(_16221_),
    .ZN(_16222_)
  );
  AND2_X1 _51550_ (
    .A1(_16220_),
    .A2(_16222_),
    .ZN(_16223_)
  );
  INV_X1 _51551_ (
    .A(_16223_),
    .ZN(_01155_)
  );
  AND2_X1 _51552_ (
    .A1(_12665_),
    .A2(_13003_),
    .ZN(_16224_)
  );
  INV_X1 _51553_ (
    .A(_16224_),
    .ZN(_16225_)
  );
  AND2_X1 _51554_ (
    .A1(\cpuregs[5] [9]),
    .A2(_12666_),
    .ZN(_16226_)
  );
  INV_X1 _51555_ (
    .A(_16226_),
    .ZN(_16227_)
  );
  AND2_X1 _51556_ (
    .A1(_16225_),
    .A2(_16227_),
    .ZN(_16228_)
  );
  INV_X1 _51557_ (
    .A(_16228_),
    .ZN(_01156_)
  );
  AND2_X1 _51558_ (
    .A1(_12665_),
    .A2(_13018_),
    .ZN(_16229_)
  );
  INV_X1 _51559_ (
    .A(_16229_),
    .ZN(_16230_)
  );
  AND2_X1 _51560_ (
    .A1(\cpuregs[5] [10]),
    .A2(_12666_),
    .ZN(_16231_)
  );
  INV_X1 _51561_ (
    .A(_16231_),
    .ZN(_16232_)
  );
  AND2_X1 _51562_ (
    .A1(_16230_),
    .A2(_16232_),
    .ZN(_16233_)
  );
  INV_X1 _51563_ (
    .A(_16233_),
    .ZN(_01157_)
  );
  AND2_X1 _51564_ (
    .A1(_12665_),
    .A2(_13033_),
    .ZN(_16234_)
  );
  INV_X1 _51565_ (
    .A(_16234_),
    .ZN(_16235_)
  );
  AND2_X1 _51566_ (
    .A1(\cpuregs[5] [11]),
    .A2(_12666_),
    .ZN(_16236_)
  );
  INV_X1 _51567_ (
    .A(_16236_),
    .ZN(_16237_)
  );
  AND2_X1 _51568_ (
    .A1(_16235_),
    .A2(_16237_),
    .ZN(_16238_)
  );
  INV_X1 _51569_ (
    .A(_16238_),
    .ZN(_01158_)
  );
  AND2_X1 _51570_ (
    .A1(_12665_),
    .A2(_13048_),
    .ZN(_16239_)
  );
  INV_X1 _51571_ (
    .A(_16239_),
    .ZN(_16240_)
  );
  AND2_X1 _51572_ (
    .A1(\cpuregs[5] [12]),
    .A2(_12666_),
    .ZN(_16241_)
  );
  INV_X1 _51573_ (
    .A(_16241_),
    .ZN(_16242_)
  );
  AND2_X1 _51574_ (
    .A1(_16240_),
    .A2(_16242_),
    .ZN(_16243_)
  );
  INV_X1 _51575_ (
    .A(_16243_),
    .ZN(_01159_)
  );
  AND2_X1 _51576_ (
    .A1(_12665_),
    .A2(_13063_),
    .ZN(_16244_)
  );
  INV_X1 _51577_ (
    .A(_16244_),
    .ZN(_16245_)
  );
  AND2_X1 _51578_ (
    .A1(\cpuregs[5] [13]),
    .A2(_12666_),
    .ZN(_16246_)
  );
  INV_X1 _51579_ (
    .A(_16246_),
    .ZN(_16247_)
  );
  AND2_X1 _51580_ (
    .A1(_16245_),
    .A2(_16247_),
    .ZN(_16248_)
  );
  INV_X1 _51581_ (
    .A(_16248_),
    .ZN(_01160_)
  );
  AND2_X1 _51582_ (
    .A1(_12665_),
    .A2(_13078_),
    .ZN(_16249_)
  );
  INV_X1 _51583_ (
    .A(_16249_),
    .ZN(_16250_)
  );
  AND2_X1 _51584_ (
    .A1(\cpuregs[5] [14]),
    .A2(_12666_),
    .ZN(_16251_)
  );
  INV_X1 _51585_ (
    .A(_16251_),
    .ZN(_16252_)
  );
  AND2_X1 _51586_ (
    .A1(_16250_),
    .A2(_16252_),
    .ZN(_16253_)
  );
  INV_X1 _51587_ (
    .A(_16253_),
    .ZN(_01161_)
  );
  AND2_X1 _51588_ (
    .A1(_12665_),
    .A2(_13093_),
    .ZN(_16254_)
  );
  INV_X1 _51589_ (
    .A(_16254_),
    .ZN(_16255_)
  );
  AND2_X1 _51590_ (
    .A1(\cpuregs[5] [15]),
    .A2(_12666_),
    .ZN(_16256_)
  );
  INV_X1 _51591_ (
    .A(_16256_),
    .ZN(_16257_)
  );
  AND2_X1 _51592_ (
    .A1(_16255_),
    .A2(_16257_),
    .ZN(_16258_)
  );
  INV_X1 _51593_ (
    .A(_16258_),
    .ZN(_01162_)
  );
  AND2_X1 _51594_ (
    .A1(_12665_),
    .A2(_13108_),
    .ZN(_16259_)
  );
  INV_X1 _51595_ (
    .A(_16259_),
    .ZN(_16260_)
  );
  AND2_X1 _51596_ (
    .A1(\cpuregs[5] [16]),
    .A2(_12666_),
    .ZN(_16261_)
  );
  INV_X1 _51597_ (
    .A(_16261_),
    .ZN(_16262_)
  );
  AND2_X1 _51598_ (
    .A1(_16260_),
    .A2(_16262_),
    .ZN(_16263_)
  );
  INV_X1 _51599_ (
    .A(_16263_),
    .ZN(_01163_)
  );
  AND2_X1 _51600_ (
    .A1(_12665_),
    .A2(_13123_),
    .ZN(_16264_)
  );
  INV_X1 _51601_ (
    .A(_16264_),
    .ZN(_16265_)
  );
  AND2_X1 _51602_ (
    .A1(\cpuregs[5] [17]),
    .A2(_12666_),
    .ZN(_16266_)
  );
  INV_X1 _51603_ (
    .A(_16266_),
    .ZN(_16267_)
  );
  AND2_X1 _51604_ (
    .A1(_16265_),
    .A2(_16267_),
    .ZN(_16268_)
  );
  INV_X1 _51605_ (
    .A(_16268_),
    .ZN(_01164_)
  );
  AND2_X1 _51606_ (
    .A1(_12665_),
    .A2(_13139_),
    .ZN(_16269_)
  );
  INV_X1 _51607_ (
    .A(_16269_),
    .ZN(_16270_)
  );
  AND2_X1 _51608_ (
    .A1(\cpuregs[5] [18]),
    .A2(_12666_),
    .ZN(_16271_)
  );
  INV_X1 _51609_ (
    .A(_16271_),
    .ZN(_16272_)
  );
  AND2_X1 _51610_ (
    .A1(_16270_),
    .A2(_16272_),
    .ZN(_16273_)
  );
  INV_X1 _51611_ (
    .A(_16273_),
    .ZN(_01165_)
  );
  AND2_X1 _51612_ (
    .A1(_12665_),
    .A2(_13154_),
    .ZN(_16274_)
  );
  INV_X1 _51613_ (
    .A(_16274_),
    .ZN(_16275_)
  );
  AND2_X1 _51614_ (
    .A1(\cpuregs[5] [19]),
    .A2(_12666_),
    .ZN(_16276_)
  );
  INV_X1 _51615_ (
    .A(_16276_),
    .ZN(_16277_)
  );
  AND2_X1 _51616_ (
    .A1(_16275_),
    .A2(_16277_),
    .ZN(_16278_)
  );
  INV_X1 _51617_ (
    .A(_16278_),
    .ZN(_01166_)
  );
  AND2_X1 _51618_ (
    .A1(_12665_),
    .A2(_13169_),
    .ZN(_16279_)
  );
  INV_X1 _51619_ (
    .A(_16279_),
    .ZN(_16280_)
  );
  AND2_X1 _51620_ (
    .A1(\cpuregs[5] [20]),
    .A2(_12666_),
    .ZN(_16281_)
  );
  INV_X1 _51621_ (
    .A(_16281_),
    .ZN(_16282_)
  );
  AND2_X1 _51622_ (
    .A1(_16280_),
    .A2(_16282_),
    .ZN(_16283_)
  );
  INV_X1 _51623_ (
    .A(_16283_),
    .ZN(_01167_)
  );
  AND2_X1 _51624_ (
    .A1(_12665_),
    .A2(_13184_),
    .ZN(_16284_)
  );
  INV_X1 _51625_ (
    .A(_16284_),
    .ZN(_16285_)
  );
  AND2_X1 _51626_ (
    .A1(\cpuregs[5] [21]),
    .A2(_12666_),
    .ZN(_16286_)
  );
  INV_X1 _51627_ (
    .A(_16286_),
    .ZN(_16287_)
  );
  AND2_X1 _51628_ (
    .A1(_16285_),
    .A2(_16287_),
    .ZN(_16288_)
  );
  INV_X1 _51629_ (
    .A(_16288_),
    .ZN(_01168_)
  );
  AND2_X1 _51630_ (
    .A1(_12665_),
    .A2(_13199_),
    .ZN(_16289_)
  );
  INV_X1 _51631_ (
    .A(_16289_),
    .ZN(_16290_)
  );
  AND2_X1 _51632_ (
    .A1(\cpuregs[5] [22]),
    .A2(_12666_),
    .ZN(_16291_)
  );
  INV_X1 _51633_ (
    .A(_16291_),
    .ZN(_16292_)
  );
  AND2_X1 _51634_ (
    .A1(_16290_),
    .A2(_16292_),
    .ZN(_16293_)
  );
  INV_X1 _51635_ (
    .A(_16293_),
    .ZN(_01169_)
  );
  AND2_X1 _51636_ (
    .A1(_12665_),
    .A2(_13214_),
    .ZN(_16294_)
  );
  INV_X1 _51637_ (
    .A(_16294_),
    .ZN(_16295_)
  );
  AND2_X1 _51638_ (
    .A1(\cpuregs[5] [23]),
    .A2(_12666_),
    .ZN(_16296_)
  );
  INV_X1 _51639_ (
    .A(_16296_),
    .ZN(_16297_)
  );
  AND2_X1 _51640_ (
    .A1(_16295_),
    .A2(_16297_),
    .ZN(_16298_)
  );
  INV_X1 _51641_ (
    .A(_16298_),
    .ZN(_01170_)
  );
  AND2_X1 _51642_ (
    .A1(_12665_),
    .A2(_13229_),
    .ZN(_16299_)
  );
  INV_X1 _51643_ (
    .A(_16299_),
    .ZN(_16300_)
  );
  AND2_X1 _51644_ (
    .A1(\cpuregs[5] [24]),
    .A2(_12666_),
    .ZN(_16301_)
  );
  INV_X1 _51645_ (
    .A(_16301_),
    .ZN(_16302_)
  );
  AND2_X1 _51646_ (
    .A1(_16300_),
    .A2(_16302_),
    .ZN(_16303_)
  );
  INV_X1 _51647_ (
    .A(_16303_),
    .ZN(_01171_)
  );
  AND2_X1 _51648_ (
    .A1(_12665_),
    .A2(_13244_),
    .ZN(_16304_)
  );
  INV_X1 _51649_ (
    .A(_16304_),
    .ZN(_16305_)
  );
  AND2_X1 _51650_ (
    .A1(\cpuregs[5] [25]),
    .A2(_12666_),
    .ZN(_16306_)
  );
  INV_X1 _51651_ (
    .A(_16306_),
    .ZN(_16307_)
  );
  AND2_X1 _51652_ (
    .A1(_16305_),
    .A2(_16307_),
    .ZN(_16308_)
  );
  INV_X1 _51653_ (
    .A(_16308_),
    .ZN(_01172_)
  );
  AND2_X1 _51654_ (
    .A1(_12665_),
    .A2(_13259_),
    .ZN(_16309_)
  );
  INV_X1 _51655_ (
    .A(_16309_),
    .ZN(_16310_)
  );
  AND2_X1 _51656_ (
    .A1(\cpuregs[5] [26]),
    .A2(_12666_),
    .ZN(_16311_)
  );
  INV_X1 _51657_ (
    .A(_16311_),
    .ZN(_16312_)
  );
  AND2_X1 _51658_ (
    .A1(_16310_),
    .A2(_16312_),
    .ZN(_16313_)
  );
  INV_X1 _51659_ (
    .A(_16313_),
    .ZN(_01173_)
  );
  AND2_X1 _51660_ (
    .A1(_12665_),
    .A2(_13274_),
    .ZN(_16314_)
  );
  INV_X1 _51661_ (
    .A(_16314_),
    .ZN(_16315_)
  );
  AND2_X1 _51662_ (
    .A1(\cpuregs[5] [27]),
    .A2(_12666_),
    .ZN(_16316_)
  );
  INV_X1 _51663_ (
    .A(_16316_),
    .ZN(_16317_)
  );
  AND2_X1 _51664_ (
    .A1(_16315_),
    .A2(_16317_),
    .ZN(_16318_)
  );
  INV_X1 _51665_ (
    .A(_16318_),
    .ZN(_01174_)
  );
  AND2_X1 _51666_ (
    .A1(_12665_),
    .A2(_13289_),
    .ZN(_16319_)
  );
  INV_X1 _51667_ (
    .A(_16319_),
    .ZN(_16320_)
  );
  AND2_X1 _51668_ (
    .A1(\cpuregs[5] [28]),
    .A2(_12666_),
    .ZN(_16321_)
  );
  INV_X1 _51669_ (
    .A(_16321_),
    .ZN(_16322_)
  );
  AND2_X1 _51670_ (
    .A1(_16320_),
    .A2(_16322_),
    .ZN(_16323_)
  );
  INV_X1 _51671_ (
    .A(_16323_),
    .ZN(_01175_)
  );
  AND2_X1 _51672_ (
    .A1(_12665_),
    .A2(_13304_),
    .ZN(_16324_)
  );
  INV_X1 _51673_ (
    .A(_16324_),
    .ZN(_16325_)
  );
  AND2_X1 _51674_ (
    .A1(\cpuregs[5] [29]),
    .A2(_12666_),
    .ZN(_16326_)
  );
  INV_X1 _51675_ (
    .A(_16326_),
    .ZN(_16327_)
  );
  AND2_X1 _51676_ (
    .A1(_16325_),
    .A2(_16327_),
    .ZN(_16328_)
  );
  INV_X1 _51677_ (
    .A(_16328_),
    .ZN(_01176_)
  );
  AND2_X1 _51678_ (
    .A1(_12665_),
    .A2(_13319_),
    .ZN(_16329_)
  );
  INV_X1 _51679_ (
    .A(_16329_),
    .ZN(_16330_)
  );
  AND2_X1 _51680_ (
    .A1(\cpuregs[5] [30]),
    .A2(_12666_),
    .ZN(_16331_)
  );
  INV_X1 _51681_ (
    .A(_16331_),
    .ZN(_16332_)
  );
  AND2_X1 _51682_ (
    .A1(_16330_),
    .A2(_16332_),
    .ZN(_16333_)
  );
  INV_X1 _51683_ (
    .A(_16333_),
    .ZN(_01177_)
  );
  AND2_X1 _51684_ (
    .A1(_12769_),
    .A2(_12874_),
    .ZN(_16334_)
  );
  INV_X1 _51685_ (
    .A(_16334_),
    .ZN(_16335_)
  );
  AND2_X1 _51686_ (
    .A1(\cpuregs[21] [0]),
    .A2(_12770_),
    .ZN(_16336_)
  );
  INV_X1 _51687_ (
    .A(_16336_),
    .ZN(_16337_)
  );
  AND2_X1 _51688_ (
    .A1(_16335_),
    .A2(_16337_),
    .ZN(_16338_)
  );
  INV_X1 _51689_ (
    .A(_16338_),
    .ZN(_01178_)
  );
  AND2_X1 _51690_ (
    .A1(_12769_),
    .A2(_12886_),
    .ZN(_16339_)
  );
  INV_X1 _51691_ (
    .A(_16339_),
    .ZN(_16340_)
  );
  AND2_X1 _51692_ (
    .A1(\cpuregs[21] [1]),
    .A2(_12770_),
    .ZN(_16341_)
  );
  INV_X1 _51693_ (
    .A(_16341_),
    .ZN(_16342_)
  );
  AND2_X1 _51694_ (
    .A1(_16340_),
    .A2(_16342_),
    .ZN(_16343_)
  );
  INV_X1 _51695_ (
    .A(_16343_),
    .ZN(_01179_)
  );
  AND2_X1 _51696_ (
    .A1(_12769_),
    .A2(_12900_),
    .ZN(_16344_)
  );
  INV_X1 _51697_ (
    .A(_16344_),
    .ZN(_16345_)
  );
  AND2_X1 _51698_ (
    .A1(\cpuregs[21] [2]),
    .A2(_12770_),
    .ZN(_16346_)
  );
  INV_X1 _51699_ (
    .A(_16346_),
    .ZN(_16347_)
  );
  AND2_X1 _51700_ (
    .A1(_16345_),
    .A2(_16347_),
    .ZN(_16348_)
  );
  INV_X1 _51701_ (
    .A(_16348_),
    .ZN(_01180_)
  );
  AND2_X1 _51702_ (
    .A1(_12769_),
    .A2(_12913_),
    .ZN(_16349_)
  );
  INV_X1 _51703_ (
    .A(_16349_),
    .ZN(_16350_)
  );
  AND2_X1 _51704_ (
    .A1(\cpuregs[21] [3]),
    .A2(_12770_),
    .ZN(_16351_)
  );
  INV_X1 _51705_ (
    .A(_16351_),
    .ZN(_16352_)
  );
  AND2_X1 _51706_ (
    .A1(_16350_),
    .A2(_16352_),
    .ZN(_16353_)
  );
  INV_X1 _51707_ (
    .A(_16353_),
    .ZN(_01181_)
  );
  AND2_X1 _51708_ (
    .A1(_12769_),
    .A2(_12928_),
    .ZN(_16354_)
  );
  INV_X1 _51709_ (
    .A(_16354_),
    .ZN(_16355_)
  );
  AND2_X1 _51710_ (
    .A1(\cpuregs[21] [4]),
    .A2(_12770_),
    .ZN(_16356_)
  );
  INV_X1 _51711_ (
    .A(_16356_),
    .ZN(_16357_)
  );
  AND2_X1 _51712_ (
    .A1(_16355_),
    .A2(_16357_),
    .ZN(_16358_)
  );
  INV_X1 _51713_ (
    .A(_16358_),
    .ZN(_01182_)
  );
  AND2_X1 _51714_ (
    .A1(_12769_),
    .A2(_12943_),
    .ZN(_16359_)
  );
  INV_X1 _51715_ (
    .A(_16359_),
    .ZN(_16360_)
  );
  AND2_X1 _51716_ (
    .A1(\cpuregs[21] [5]),
    .A2(_12770_),
    .ZN(_16361_)
  );
  INV_X1 _51717_ (
    .A(_16361_),
    .ZN(_16362_)
  );
  AND2_X1 _51718_ (
    .A1(_16360_),
    .A2(_16362_),
    .ZN(_16363_)
  );
  INV_X1 _51719_ (
    .A(_16363_),
    .ZN(_01183_)
  );
  AND2_X1 _51720_ (
    .A1(_12769_),
    .A2(_12958_),
    .ZN(_16364_)
  );
  INV_X1 _51721_ (
    .A(_16364_),
    .ZN(_16365_)
  );
  AND2_X1 _51722_ (
    .A1(\cpuregs[21] [6]),
    .A2(_12770_),
    .ZN(_16366_)
  );
  INV_X1 _51723_ (
    .A(_16366_),
    .ZN(_16367_)
  );
  AND2_X1 _51724_ (
    .A1(_16365_),
    .A2(_16367_),
    .ZN(_16368_)
  );
  INV_X1 _51725_ (
    .A(_16368_),
    .ZN(_01184_)
  );
  AND2_X1 _51726_ (
    .A1(_12769_),
    .A2(_12973_),
    .ZN(_16369_)
  );
  INV_X1 _51727_ (
    .A(_16369_),
    .ZN(_16370_)
  );
  AND2_X1 _51728_ (
    .A1(\cpuregs[21] [7]),
    .A2(_12770_),
    .ZN(_16371_)
  );
  INV_X1 _51729_ (
    .A(_16371_),
    .ZN(_16372_)
  );
  AND2_X1 _51730_ (
    .A1(_16370_),
    .A2(_16372_),
    .ZN(_16373_)
  );
  INV_X1 _51731_ (
    .A(_16373_),
    .ZN(_01185_)
  );
  AND2_X1 _51732_ (
    .A1(_12769_),
    .A2(_12988_),
    .ZN(_16374_)
  );
  INV_X1 _51733_ (
    .A(_16374_),
    .ZN(_16375_)
  );
  AND2_X1 _51734_ (
    .A1(\cpuregs[21] [8]),
    .A2(_12770_),
    .ZN(_16376_)
  );
  INV_X1 _51735_ (
    .A(_16376_),
    .ZN(_16377_)
  );
  AND2_X1 _51736_ (
    .A1(_16375_),
    .A2(_16377_),
    .ZN(_16378_)
  );
  INV_X1 _51737_ (
    .A(_16378_),
    .ZN(_01186_)
  );
  AND2_X1 _51738_ (
    .A1(_12769_),
    .A2(_13003_),
    .ZN(_16379_)
  );
  INV_X1 _51739_ (
    .A(_16379_),
    .ZN(_16380_)
  );
  AND2_X1 _51740_ (
    .A1(\cpuregs[21] [9]),
    .A2(_12770_),
    .ZN(_16381_)
  );
  INV_X1 _51741_ (
    .A(_16381_),
    .ZN(_16382_)
  );
  AND2_X1 _51742_ (
    .A1(_16380_),
    .A2(_16382_),
    .ZN(_16383_)
  );
  INV_X1 _51743_ (
    .A(_16383_),
    .ZN(_01187_)
  );
  AND2_X1 _51744_ (
    .A1(_12769_),
    .A2(_13018_),
    .ZN(_16384_)
  );
  INV_X1 _51745_ (
    .A(_16384_),
    .ZN(_16385_)
  );
  AND2_X1 _51746_ (
    .A1(\cpuregs[21] [10]),
    .A2(_12770_),
    .ZN(_16386_)
  );
  INV_X1 _51747_ (
    .A(_16386_),
    .ZN(_16387_)
  );
  AND2_X1 _51748_ (
    .A1(_16385_),
    .A2(_16387_),
    .ZN(_16388_)
  );
  INV_X1 _51749_ (
    .A(_16388_),
    .ZN(_01188_)
  );
  AND2_X1 _51750_ (
    .A1(_12769_),
    .A2(_13033_),
    .ZN(_16389_)
  );
  INV_X1 _51751_ (
    .A(_16389_),
    .ZN(_16390_)
  );
  AND2_X1 _51752_ (
    .A1(\cpuregs[21] [11]),
    .A2(_12770_),
    .ZN(_16391_)
  );
  INV_X1 _51753_ (
    .A(_16391_),
    .ZN(_16392_)
  );
  AND2_X1 _51754_ (
    .A1(_16390_),
    .A2(_16392_),
    .ZN(_16393_)
  );
  INV_X1 _51755_ (
    .A(_16393_),
    .ZN(_01189_)
  );
  AND2_X1 _51756_ (
    .A1(_12769_),
    .A2(_13048_),
    .ZN(_16394_)
  );
  INV_X1 _51757_ (
    .A(_16394_),
    .ZN(_16395_)
  );
  AND2_X1 _51758_ (
    .A1(\cpuregs[21] [12]),
    .A2(_12770_),
    .ZN(_16396_)
  );
  INV_X1 _51759_ (
    .A(_16396_),
    .ZN(_16397_)
  );
  AND2_X1 _51760_ (
    .A1(_16395_),
    .A2(_16397_),
    .ZN(_16398_)
  );
  INV_X1 _51761_ (
    .A(_16398_),
    .ZN(_01190_)
  );
  AND2_X1 _51762_ (
    .A1(_12769_),
    .A2(_13063_),
    .ZN(_16399_)
  );
  INV_X1 _51763_ (
    .A(_16399_),
    .ZN(_16400_)
  );
  AND2_X1 _51764_ (
    .A1(\cpuregs[21] [13]),
    .A2(_12770_),
    .ZN(_16401_)
  );
  INV_X1 _51765_ (
    .A(_16401_),
    .ZN(_16402_)
  );
  AND2_X1 _51766_ (
    .A1(_16400_),
    .A2(_16402_),
    .ZN(_16403_)
  );
  INV_X1 _51767_ (
    .A(_16403_),
    .ZN(_01191_)
  );
  AND2_X1 _51768_ (
    .A1(_12769_),
    .A2(_13078_),
    .ZN(_16404_)
  );
  INV_X1 _51769_ (
    .A(_16404_),
    .ZN(_16405_)
  );
  AND2_X1 _51770_ (
    .A1(\cpuregs[21] [14]),
    .A2(_12770_),
    .ZN(_16406_)
  );
  INV_X1 _51771_ (
    .A(_16406_),
    .ZN(_16407_)
  );
  AND2_X1 _51772_ (
    .A1(_16405_),
    .A2(_16407_),
    .ZN(_16408_)
  );
  INV_X1 _51773_ (
    .A(_16408_),
    .ZN(_01192_)
  );
  AND2_X1 _51774_ (
    .A1(_12769_),
    .A2(_13093_),
    .ZN(_16409_)
  );
  INV_X1 _51775_ (
    .A(_16409_),
    .ZN(_16410_)
  );
  AND2_X1 _51776_ (
    .A1(\cpuregs[21] [15]),
    .A2(_12770_),
    .ZN(_16411_)
  );
  INV_X1 _51777_ (
    .A(_16411_),
    .ZN(_16412_)
  );
  AND2_X1 _51778_ (
    .A1(_16410_),
    .A2(_16412_),
    .ZN(_16413_)
  );
  INV_X1 _51779_ (
    .A(_16413_),
    .ZN(_01193_)
  );
  AND2_X1 _51780_ (
    .A1(_12769_),
    .A2(_13108_),
    .ZN(_16414_)
  );
  INV_X1 _51781_ (
    .A(_16414_),
    .ZN(_16415_)
  );
  AND2_X1 _51782_ (
    .A1(\cpuregs[21] [16]),
    .A2(_12770_),
    .ZN(_16416_)
  );
  INV_X1 _51783_ (
    .A(_16416_),
    .ZN(_16417_)
  );
  AND2_X1 _51784_ (
    .A1(_16415_),
    .A2(_16417_),
    .ZN(_16418_)
  );
  INV_X1 _51785_ (
    .A(_16418_),
    .ZN(_01194_)
  );
  AND2_X1 _51786_ (
    .A1(_12769_),
    .A2(_13123_),
    .ZN(_16419_)
  );
  INV_X1 _51787_ (
    .A(_16419_),
    .ZN(_16420_)
  );
  AND2_X1 _51788_ (
    .A1(\cpuregs[21] [17]),
    .A2(_12770_),
    .ZN(_16421_)
  );
  INV_X1 _51789_ (
    .A(_16421_),
    .ZN(_16422_)
  );
  AND2_X1 _51790_ (
    .A1(_16420_),
    .A2(_16422_),
    .ZN(_16423_)
  );
  INV_X1 _51791_ (
    .A(_16423_),
    .ZN(_01195_)
  );
  AND2_X1 _51792_ (
    .A1(_12769_),
    .A2(_13139_),
    .ZN(_16424_)
  );
  INV_X1 _51793_ (
    .A(_16424_),
    .ZN(_16425_)
  );
  AND2_X1 _51794_ (
    .A1(\cpuregs[21] [18]),
    .A2(_12770_),
    .ZN(_16426_)
  );
  INV_X1 _51795_ (
    .A(_16426_),
    .ZN(_16427_)
  );
  AND2_X1 _51796_ (
    .A1(_16425_),
    .A2(_16427_),
    .ZN(_16428_)
  );
  INV_X1 _51797_ (
    .A(_16428_),
    .ZN(_01196_)
  );
  AND2_X1 _51798_ (
    .A1(_12769_),
    .A2(_13154_),
    .ZN(_16429_)
  );
  INV_X1 _51799_ (
    .A(_16429_),
    .ZN(_16430_)
  );
  AND2_X1 _51800_ (
    .A1(\cpuregs[21] [19]),
    .A2(_12770_),
    .ZN(_16431_)
  );
  INV_X1 _51801_ (
    .A(_16431_),
    .ZN(_16432_)
  );
  AND2_X1 _51802_ (
    .A1(_16430_),
    .A2(_16432_),
    .ZN(_16433_)
  );
  INV_X1 _51803_ (
    .A(_16433_),
    .ZN(_01197_)
  );
  AND2_X1 _51804_ (
    .A1(_12769_),
    .A2(_13169_),
    .ZN(_16434_)
  );
  INV_X1 _51805_ (
    .A(_16434_),
    .ZN(_16435_)
  );
  AND2_X1 _51806_ (
    .A1(\cpuregs[21] [20]),
    .A2(_12770_),
    .ZN(_16436_)
  );
  INV_X1 _51807_ (
    .A(_16436_),
    .ZN(_16437_)
  );
  AND2_X1 _51808_ (
    .A1(_16435_),
    .A2(_16437_),
    .ZN(_16438_)
  );
  INV_X1 _51809_ (
    .A(_16438_),
    .ZN(_01198_)
  );
  AND2_X1 _51810_ (
    .A1(_12769_),
    .A2(_13184_),
    .ZN(_16439_)
  );
  INV_X1 _51811_ (
    .A(_16439_),
    .ZN(_16440_)
  );
  AND2_X1 _51812_ (
    .A1(\cpuregs[21] [21]),
    .A2(_12770_),
    .ZN(_16441_)
  );
  INV_X1 _51813_ (
    .A(_16441_),
    .ZN(_16442_)
  );
  AND2_X1 _51814_ (
    .A1(_16440_),
    .A2(_16442_),
    .ZN(_16443_)
  );
  INV_X1 _51815_ (
    .A(_16443_),
    .ZN(_01199_)
  );
  AND2_X1 _51816_ (
    .A1(_12769_),
    .A2(_13199_),
    .ZN(_16444_)
  );
  INV_X1 _51817_ (
    .A(_16444_),
    .ZN(_16445_)
  );
  AND2_X1 _51818_ (
    .A1(\cpuregs[21] [22]),
    .A2(_12770_),
    .ZN(_16446_)
  );
  INV_X1 _51819_ (
    .A(_16446_),
    .ZN(_16447_)
  );
  AND2_X1 _51820_ (
    .A1(_16445_),
    .A2(_16447_),
    .ZN(_16448_)
  );
  INV_X1 _51821_ (
    .A(_16448_),
    .ZN(_01200_)
  );
  AND2_X1 _51822_ (
    .A1(_12769_),
    .A2(_13214_),
    .ZN(_16449_)
  );
  INV_X1 _51823_ (
    .A(_16449_),
    .ZN(_16450_)
  );
  AND2_X1 _51824_ (
    .A1(\cpuregs[21] [23]),
    .A2(_12770_),
    .ZN(_16451_)
  );
  INV_X1 _51825_ (
    .A(_16451_),
    .ZN(_16452_)
  );
  AND2_X1 _51826_ (
    .A1(_16450_),
    .A2(_16452_),
    .ZN(_16453_)
  );
  INV_X1 _51827_ (
    .A(_16453_),
    .ZN(_01201_)
  );
  AND2_X1 _51828_ (
    .A1(_12769_),
    .A2(_13229_),
    .ZN(_16454_)
  );
  INV_X1 _51829_ (
    .A(_16454_),
    .ZN(_16455_)
  );
  AND2_X1 _51830_ (
    .A1(\cpuregs[21] [24]),
    .A2(_12770_),
    .ZN(_16456_)
  );
  INV_X1 _51831_ (
    .A(_16456_),
    .ZN(_16457_)
  );
  AND2_X1 _51832_ (
    .A1(_16455_),
    .A2(_16457_),
    .ZN(_16458_)
  );
  INV_X1 _51833_ (
    .A(_16458_),
    .ZN(_01202_)
  );
  AND2_X1 _51834_ (
    .A1(_12769_),
    .A2(_13244_),
    .ZN(_16459_)
  );
  INV_X1 _51835_ (
    .A(_16459_),
    .ZN(_16460_)
  );
  AND2_X1 _51836_ (
    .A1(\cpuregs[21] [25]),
    .A2(_12770_),
    .ZN(_16461_)
  );
  INV_X1 _51837_ (
    .A(_16461_),
    .ZN(_16462_)
  );
  AND2_X1 _51838_ (
    .A1(_16460_),
    .A2(_16462_),
    .ZN(_16463_)
  );
  INV_X1 _51839_ (
    .A(_16463_),
    .ZN(_01203_)
  );
  AND2_X1 _51840_ (
    .A1(_12769_),
    .A2(_13259_),
    .ZN(_16464_)
  );
  INV_X1 _51841_ (
    .A(_16464_),
    .ZN(_16465_)
  );
  AND2_X1 _51842_ (
    .A1(\cpuregs[21] [26]),
    .A2(_12770_),
    .ZN(_16466_)
  );
  INV_X1 _51843_ (
    .A(_16466_),
    .ZN(_16467_)
  );
  AND2_X1 _51844_ (
    .A1(_16465_),
    .A2(_16467_),
    .ZN(_16468_)
  );
  INV_X1 _51845_ (
    .A(_16468_),
    .ZN(_01204_)
  );
  AND2_X1 _51846_ (
    .A1(_12769_),
    .A2(_13274_),
    .ZN(_16469_)
  );
  INV_X1 _51847_ (
    .A(_16469_),
    .ZN(_16470_)
  );
  AND2_X1 _51848_ (
    .A1(\cpuregs[21] [27]),
    .A2(_12770_),
    .ZN(_16471_)
  );
  INV_X1 _51849_ (
    .A(_16471_),
    .ZN(_16472_)
  );
  AND2_X1 _51850_ (
    .A1(_16470_),
    .A2(_16472_),
    .ZN(_16473_)
  );
  INV_X1 _51851_ (
    .A(_16473_),
    .ZN(_01205_)
  );
  AND2_X1 _51852_ (
    .A1(_12769_),
    .A2(_13289_),
    .ZN(_16474_)
  );
  INV_X1 _51853_ (
    .A(_16474_),
    .ZN(_16475_)
  );
  AND2_X1 _51854_ (
    .A1(\cpuregs[21] [28]),
    .A2(_12770_),
    .ZN(_16476_)
  );
  INV_X1 _51855_ (
    .A(_16476_),
    .ZN(_16477_)
  );
  AND2_X1 _51856_ (
    .A1(_16475_),
    .A2(_16477_),
    .ZN(_16478_)
  );
  INV_X1 _51857_ (
    .A(_16478_),
    .ZN(_01206_)
  );
  AND2_X1 _51858_ (
    .A1(_12769_),
    .A2(_13304_),
    .ZN(_16479_)
  );
  INV_X1 _51859_ (
    .A(_16479_),
    .ZN(_16480_)
  );
  AND2_X1 _51860_ (
    .A1(\cpuregs[21] [29]),
    .A2(_12770_),
    .ZN(_16481_)
  );
  INV_X1 _51861_ (
    .A(_16481_),
    .ZN(_16482_)
  );
  AND2_X1 _51862_ (
    .A1(_16480_),
    .A2(_16482_),
    .ZN(_16483_)
  );
  INV_X1 _51863_ (
    .A(_16483_),
    .ZN(_01207_)
  );
  AND2_X1 _51864_ (
    .A1(_12769_),
    .A2(_13319_),
    .ZN(_16484_)
  );
  INV_X1 _51865_ (
    .A(_16484_),
    .ZN(_16485_)
  );
  AND2_X1 _51866_ (
    .A1(\cpuregs[21] [30]),
    .A2(_12770_),
    .ZN(_16486_)
  );
  INV_X1 _51867_ (
    .A(_16486_),
    .ZN(_16487_)
  );
  AND2_X1 _51868_ (
    .A1(_16485_),
    .A2(_16487_),
    .ZN(_16488_)
  );
  INV_X1 _51869_ (
    .A(_16488_),
    .ZN(_01208_)
  );
  AND2_X1 _51870_ (
    .A1(_12650_),
    .A2(_12874_),
    .ZN(_16489_)
  );
  INV_X1 _51871_ (
    .A(_16489_),
    .ZN(_16490_)
  );
  AND2_X1 _51872_ (
    .A1(\cpuregs[7] [0]),
    .A2(_12651_),
    .ZN(_16491_)
  );
  INV_X1 _51873_ (
    .A(_16491_),
    .ZN(_16492_)
  );
  AND2_X1 _51874_ (
    .A1(_16490_),
    .A2(_16492_),
    .ZN(_16493_)
  );
  INV_X1 _51875_ (
    .A(_16493_),
    .ZN(_01209_)
  );
  AND2_X1 _51876_ (
    .A1(_12650_),
    .A2(_12886_),
    .ZN(_16494_)
  );
  INV_X1 _51877_ (
    .A(_16494_),
    .ZN(_16495_)
  );
  AND2_X1 _51878_ (
    .A1(\cpuregs[7] [1]),
    .A2(_12651_),
    .ZN(_16496_)
  );
  INV_X1 _51879_ (
    .A(_16496_),
    .ZN(_16497_)
  );
  AND2_X1 _51880_ (
    .A1(_16495_),
    .A2(_16497_),
    .ZN(_16498_)
  );
  INV_X1 _51881_ (
    .A(_16498_),
    .ZN(_01210_)
  );
  AND2_X1 _51882_ (
    .A1(_12650_),
    .A2(_12900_),
    .ZN(_16499_)
  );
  INV_X1 _51883_ (
    .A(_16499_),
    .ZN(_16500_)
  );
  AND2_X1 _51884_ (
    .A1(\cpuregs[7] [2]),
    .A2(_12651_),
    .ZN(_16501_)
  );
  INV_X1 _51885_ (
    .A(_16501_),
    .ZN(_16502_)
  );
  AND2_X1 _51886_ (
    .A1(_16500_),
    .A2(_16502_),
    .ZN(_16503_)
  );
  INV_X1 _51887_ (
    .A(_16503_),
    .ZN(_01211_)
  );
  AND2_X1 _51888_ (
    .A1(_12650_),
    .A2(_12913_),
    .ZN(_16504_)
  );
  INV_X1 _51889_ (
    .A(_16504_),
    .ZN(_16505_)
  );
  AND2_X1 _51890_ (
    .A1(\cpuregs[7] [3]),
    .A2(_12651_),
    .ZN(_16506_)
  );
  INV_X1 _51891_ (
    .A(_16506_),
    .ZN(_16507_)
  );
  AND2_X1 _51892_ (
    .A1(_16505_),
    .A2(_16507_),
    .ZN(_16508_)
  );
  INV_X1 _51893_ (
    .A(_16508_),
    .ZN(_01212_)
  );
  AND2_X1 _51894_ (
    .A1(\cpuregs[7] [4]),
    .A2(_12651_),
    .ZN(_16509_)
  );
  INV_X1 _51895_ (
    .A(_16509_),
    .ZN(_16510_)
  );
  AND2_X1 _51896_ (
    .A1(_12650_),
    .A2(_12928_),
    .ZN(_16511_)
  );
  INV_X1 _51897_ (
    .A(_16511_),
    .ZN(_16512_)
  );
  AND2_X1 _51898_ (
    .A1(_16510_),
    .A2(_16512_),
    .ZN(_16513_)
  );
  INV_X1 _51899_ (
    .A(_16513_),
    .ZN(_01213_)
  );
  AND2_X1 _51900_ (
    .A1(_12650_),
    .A2(_12943_),
    .ZN(_16514_)
  );
  INV_X1 _51901_ (
    .A(_16514_),
    .ZN(_16515_)
  );
  AND2_X1 _51902_ (
    .A1(\cpuregs[7] [5]),
    .A2(_12651_),
    .ZN(_16516_)
  );
  INV_X1 _51903_ (
    .A(_16516_),
    .ZN(_16517_)
  );
  AND2_X1 _51904_ (
    .A1(_16515_),
    .A2(_16517_),
    .ZN(_16518_)
  );
  INV_X1 _51905_ (
    .A(_16518_),
    .ZN(_01214_)
  );
  AND2_X1 _51906_ (
    .A1(_12650_),
    .A2(_12958_),
    .ZN(_16519_)
  );
  INV_X1 _51907_ (
    .A(_16519_),
    .ZN(_16520_)
  );
  AND2_X1 _51908_ (
    .A1(\cpuregs[7] [6]),
    .A2(_12651_),
    .ZN(_16521_)
  );
  INV_X1 _51909_ (
    .A(_16521_),
    .ZN(_16522_)
  );
  AND2_X1 _51910_ (
    .A1(_16520_),
    .A2(_16522_),
    .ZN(_16523_)
  );
  INV_X1 _51911_ (
    .A(_16523_),
    .ZN(_01215_)
  );
  AND2_X1 _51912_ (
    .A1(_12650_),
    .A2(_12973_),
    .ZN(_16524_)
  );
  INV_X1 _51913_ (
    .A(_16524_),
    .ZN(_16525_)
  );
  AND2_X1 _51914_ (
    .A1(\cpuregs[7] [7]),
    .A2(_12651_),
    .ZN(_16526_)
  );
  INV_X1 _51915_ (
    .A(_16526_),
    .ZN(_16527_)
  );
  AND2_X1 _51916_ (
    .A1(_16525_),
    .A2(_16527_),
    .ZN(_16528_)
  );
  INV_X1 _51917_ (
    .A(_16528_),
    .ZN(_01216_)
  );
  AND2_X1 _51918_ (
    .A1(_12650_),
    .A2(_12988_),
    .ZN(_16529_)
  );
  INV_X1 _51919_ (
    .A(_16529_),
    .ZN(_16530_)
  );
  AND2_X1 _51920_ (
    .A1(\cpuregs[7] [8]),
    .A2(_12651_),
    .ZN(_16531_)
  );
  INV_X1 _51921_ (
    .A(_16531_),
    .ZN(_16532_)
  );
  AND2_X1 _51922_ (
    .A1(_16530_),
    .A2(_16532_),
    .ZN(_16533_)
  );
  INV_X1 _51923_ (
    .A(_16533_),
    .ZN(_01217_)
  );
  AND2_X1 _51924_ (
    .A1(_12650_),
    .A2(_13003_),
    .ZN(_16534_)
  );
  INV_X1 _51925_ (
    .A(_16534_),
    .ZN(_16535_)
  );
  AND2_X1 _51926_ (
    .A1(\cpuregs[7] [9]),
    .A2(_12651_),
    .ZN(_16536_)
  );
  INV_X1 _51927_ (
    .A(_16536_),
    .ZN(_16537_)
  );
  AND2_X1 _51928_ (
    .A1(_16535_),
    .A2(_16537_),
    .ZN(_16538_)
  );
  INV_X1 _51929_ (
    .A(_16538_),
    .ZN(_01218_)
  );
  AND2_X1 _51930_ (
    .A1(_12650_),
    .A2(_13018_),
    .ZN(_16539_)
  );
  INV_X1 _51931_ (
    .A(_16539_),
    .ZN(_16540_)
  );
  AND2_X1 _51932_ (
    .A1(\cpuregs[7] [10]),
    .A2(_12651_),
    .ZN(_16541_)
  );
  INV_X1 _51933_ (
    .A(_16541_),
    .ZN(_16542_)
  );
  AND2_X1 _51934_ (
    .A1(_16540_),
    .A2(_16542_),
    .ZN(_16543_)
  );
  INV_X1 _51935_ (
    .A(_16543_),
    .ZN(_01219_)
  );
  AND2_X1 _51936_ (
    .A1(_12650_),
    .A2(_13033_),
    .ZN(_16544_)
  );
  INV_X1 _51937_ (
    .A(_16544_),
    .ZN(_16545_)
  );
  AND2_X1 _51938_ (
    .A1(\cpuregs[7] [11]),
    .A2(_12651_),
    .ZN(_16546_)
  );
  INV_X1 _51939_ (
    .A(_16546_),
    .ZN(_16547_)
  );
  AND2_X1 _51940_ (
    .A1(_16545_),
    .A2(_16547_),
    .ZN(_16548_)
  );
  INV_X1 _51941_ (
    .A(_16548_),
    .ZN(_01220_)
  );
  AND2_X1 _51942_ (
    .A1(_12650_),
    .A2(_13048_),
    .ZN(_16549_)
  );
  INV_X1 _51943_ (
    .A(_16549_),
    .ZN(_16550_)
  );
  AND2_X1 _51944_ (
    .A1(\cpuregs[7] [12]),
    .A2(_12651_),
    .ZN(_16551_)
  );
  INV_X1 _51945_ (
    .A(_16551_),
    .ZN(_16552_)
  );
  AND2_X1 _51946_ (
    .A1(_16550_),
    .A2(_16552_),
    .ZN(_16553_)
  );
  INV_X1 _51947_ (
    .A(_16553_),
    .ZN(_01221_)
  );
  AND2_X1 _51948_ (
    .A1(_12650_),
    .A2(_13063_),
    .ZN(_16554_)
  );
  INV_X1 _51949_ (
    .A(_16554_),
    .ZN(_16555_)
  );
  AND2_X1 _51950_ (
    .A1(\cpuregs[7] [13]),
    .A2(_12651_),
    .ZN(_16556_)
  );
  INV_X1 _51951_ (
    .A(_16556_),
    .ZN(_16557_)
  );
  AND2_X1 _51952_ (
    .A1(_16555_),
    .A2(_16557_),
    .ZN(_16558_)
  );
  INV_X1 _51953_ (
    .A(_16558_),
    .ZN(_01222_)
  );
  AND2_X1 _51954_ (
    .A1(_12650_),
    .A2(_13078_),
    .ZN(_16559_)
  );
  INV_X1 _51955_ (
    .A(_16559_),
    .ZN(_16560_)
  );
  AND2_X1 _51956_ (
    .A1(\cpuregs[7] [14]),
    .A2(_12651_),
    .ZN(_16561_)
  );
  INV_X1 _51957_ (
    .A(_16561_),
    .ZN(_16562_)
  );
  AND2_X1 _51958_ (
    .A1(_16560_),
    .A2(_16562_),
    .ZN(_16563_)
  );
  INV_X1 _51959_ (
    .A(_16563_),
    .ZN(_01223_)
  );
  AND2_X1 _51960_ (
    .A1(_12650_),
    .A2(_13093_),
    .ZN(_16564_)
  );
  INV_X1 _51961_ (
    .A(_16564_),
    .ZN(_16565_)
  );
  AND2_X1 _51962_ (
    .A1(\cpuregs[7] [15]),
    .A2(_12651_),
    .ZN(_16566_)
  );
  INV_X1 _51963_ (
    .A(_16566_),
    .ZN(_16567_)
  );
  AND2_X1 _51964_ (
    .A1(_16565_),
    .A2(_16567_),
    .ZN(_16568_)
  );
  INV_X1 _51965_ (
    .A(_16568_),
    .ZN(_01224_)
  );
  AND2_X1 _51966_ (
    .A1(_12650_),
    .A2(_13108_),
    .ZN(_16569_)
  );
  INV_X1 _51967_ (
    .A(_16569_),
    .ZN(_16570_)
  );
  AND2_X1 _51968_ (
    .A1(\cpuregs[7] [16]),
    .A2(_12651_),
    .ZN(_16571_)
  );
  INV_X1 _51969_ (
    .A(_16571_),
    .ZN(_16572_)
  );
  AND2_X1 _51970_ (
    .A1(_16570_),
    .A2(_16572_),
    .ZN(_16573_)
  );
  INV_X1 _51971_ (
    .A(_16573_),
    .ZN(_01225_)
  );
  AND2_X1 _51972_ (
    .A1(_12650_),
    .A2(_13123_),
    .ZN(_16574_)
  );
  INV_X1 _51973_ (
    .A(_16574_),
    .ZN(_16575_)
  );
  AND2_X1 _51974_ (
    .A1(\cpuregs[7] [17]),
    .A2(_12651_),
    .ZN(_16576_)
  );
  INV_X1 _51975_ (
    .A(_16576_),
    .ZN(_16577_)
  );
  AND2_X1 _51976_ (
    .A1(_16575_),
    .A2(_16577_),
    .ZN(_16578_)
  );
  INV_X1 _51977_ (
    .A(_16578_),
    .ZN(_01226_)
  );
  AND2_X1 _51978_ (
    .A1(_12650_),
    .A2(_13139_),
    .ZN(_16579_)
  );
  INV_X1 _51979_ (
    .A(_16579_),
    .ZN(_16580_)
  );
  AND2_X1 _51980_ (
    .A1(\cpuregs[7] [18]),
    .A2(_12651_),
    .ZN(_16581_)
  );
  INV_X1 _51981_ (
    .A(_16581_),
    .ZN(_16582_)
  );
  AND2_X1 _51982_ (
    .A1(_16580_),
    .A2(_16582_),
    .ZN(_16583_)
  );
  INV_X1 _51983_ (
    .A(_16583_),
    .ZN(_01227_)
  );
  AND2_X1 _51984_ (
    .A1(_12650_),
    .A2(_13154_),
    .ZN(_16584_)
  );
  INV_X1 _51985_ (
    .A(_16584_),
    .ZN(_16585_)
  );
  AND2_X1 _51986_ (
    .A1(\cpuregs[7] [19]),
    .A2(_12651_),
    .ZN(_16586_)
  );
  INV_X1 _51987_ (
    .A(_16586_),
    .ZN(_16587_)
  );
  AND2_X1 _51988_ (
    .A1(_16585_),
    .A2(_16587_),
    .ZN(_16588_)
  );
  INV_X1 _51989_ (
    .A(_16588_),
    .ZN(_01228_)
  );
  AND2_X1 _51990_ (
    .A1(_12650_),
    .A2(_13169_),
    .ZN(_16589_)
  );
  INV_X1 _51991_ (
    .A(_16589_),
    .ZN(_16590_)
  );
  AND2_X1 _51992_ (
    .A1(\cpuregs[7] [20]),
    .A2(_12651_),
    .ZN(_16591_)
  );
  INV_X1 _51993_ (
    .A(_16591_),
    .ZN(_16592_)
  );
  AND2_X1 _51994_ (
    .A1(_16590_),
    .A2(_16592_),
    .ZN(_16593_)
  );
  INV_X1 _51995_ (
    .A(_16593_),
    .ZN(_01229_)
  );
  AND2_X1 _51996_ (
    .A1(_12650_),
    .A2(_13184_),
    .ZN(_16594_)
  );
  INV_X1 _51997_ (
    .A(_16594_),
    .ZN(_16595_)
  );
  AND2_X1 _51998_ (
    .A1(\cpuregs[7] [21]),
    .A2(_12651_),
    .ZN(_16596_)
  );
  INV_X1 _51999_ (
    .A(_16596_),
    .ZN(_16597_)
  );
  AND2_X1 _52000_ (
    .A1(_16595_),
    .A2(_16597_),
    .ZN(_16598_)
  );
  INV_X1 _52001_ (
    .A(_16598_),
    .ZN(_01230_)
  );
  AND2_X1 _52002_ (
    .A1(_12650_),
    .A2(_13199_),
    .ZN(_16599_)
  );
  INV_X1 _52003_ (
    .A(_16599_),
    .ZN(_16600_)
  );
  AND2_X1 _52004_ (
    .A1(\cpuregs[7] [22]),
    .A2(_12651_),
    .ZN(_16601_)
  );
  INV_X1 _52005_ (
    .A(_16601_),
    .ZN(_16602_)
  );
  AND2_X1 _52006_ (
    .A1(_16600_),
    .A2(_16602_),
    .ZN(_16603_)
  );
  INV_X1 _52007_ (
    .A(_16603_),
    .ZN(_01231_)
  );
  AND2_X1 _52008_ (
    .A1(_12650_),
    .A2(_13214_),
    .ZN(_16604_)
  );
  INV_X1 _52009_ (
    .A(_16604_),
    .ZN(_16605_)
  );
  AND2_X1 _52010_ (
    .A1(\cpuregs[7] [23]),
    .A2(_12651_),
    .ZN(_16606_)
  );
  INV_X1 _52011_ (
    .A(_16606_),
    .ZN(_16607_)
  );
  AND2_X1 _52012_ (
    .A1(_16605_),
    .A2(_16607_),
    .ZN(_16608_)
  );
  INV_X1 _52013_ (
    .A(_16608_),
    .ZN(_01232_)
  );
  AND2_X1 _52014_ (
    .A1(_12650_),
    .A2(_13229_),
    .ZN(_16609_)
  );
  INV_X1 _52015_ (
    .A(_16609_),
    .ZN(_16610_)
  );
  AND2_X1 _52016_ (
    .A1(\cpuregs[7] [24]),
    .A2(_12651_),
    .ZN(_16611_)
  );
  INV_X1 _52017_ (
    .A(_16611_),
    .ZN(_16612_)
  );
  AND2_X1 _52018_ (
    .A1(_16610_),
    .A2(_16612_),
    .ZN(_16613_)
  );
  INV_X1 _52019_ (
    .A(_16613_),
    .ZN(_01233_)
  );
  AND2_X1 _52020_ (
    .A1(_12650_),
    .A2(_13244_),
    .ZN(_16614_)
  );
  INV_X1 _52021_ (
    .A(_16614_),
    .ZN(_16615_)
  );
  AND2_X1 _52022_ (
    .A1(\cpuregs[7] [25]),
    .A2(_12651_),
    .ZN(_16616_)
  );
  INV_X1 _52023_ (
    .A(_16616_),
    .ZN(_16617_)
  );
  AND2_X1 _52024_ (
    .A1(_16615_),
    .A2(_16617_),
    .ZN(_16618_)
  );
  INV_X1 _52025_ (
    .A(_16618_),
    .ZN(_01234_)
  );
  AND2_X1 _52026_ (
    .A1(_12650_),
    .A2(_13259_),
    .ZN(_16619_)
  );
  INV_X1 _52027_ (
    .A(_16619_),
    .ZN(_16620_)
  );
  AND2_X1 _52028_ (
    .A1(\cpuregs[7] [26]),
    .A2(_12651_),
    .ZN(_16621_)
  );
  INV_X1 _52029_ (
    .A(_16621_),
    .ZN(_16622_)
  );
  AND2_X1 _52030_ (
    .A1(_16620_),
    .A2(_16622_),
    .ZN(_16623_)
  );
  INV_X1 _52031_ (
    .A(_16623_),
    .ZN(_01235_)
  );
  AND2_X1 _52032_ (
    .A1(_12650_),
    .A2(_13274_),
    .ZN(_16624_)
  );
  INV_X1 _52033_ (
    .A(_16624_),
    .ZN(_16625_)
  );
  AND2_X1 _52034_ (
    .A1(\cpuregs[7] [27]),
    .A2(_12651_),
    .ZN(_16626_)
  );
  INV_X1 _52035_ (
    .A(_16626_),
    .ZN(_16627_)
  );
  AND2_X1 _52036_ (
    .A1(_16625_),
    .A2(_16627_),
    .ZN(_16628_)
  );
  INV_X1 _52037_ (
    .A(_16628_),
    .ZN(_01236_)
  );
  AND2_X1 _52038_ (
    .A1(_12650_),
    .A2(_13289_),
    .ZN(_16629_)
  );
  INV_X1 _52039_ (
    .A(_16629_),
    .ZN(_16630_)
  );
  AND2_X1 _52040_ (
    .A1(\cpuregs[7] [28]),
    .A2(_12651_),
    .ZN(_16631_)
  );
  INV_X1 _52041_ (
    .A(_16631_),
    .ZN(_16632_)
  );
  AND2_X1 _52042_ (
    .A1(_16630_),
    .A2(_16632_),
    .ZN(_16633_)
  );
  INV_X1 _52043_ (
    .A(_16633_),
    .ZN(_01237_)
  );
  AND2_X1 _52044_ (
    .A1(_12650_),
    .A2(_13304_),
    .ZN(_16634_)
  );
  INV_X1 _52045_ (
    .A(_16634_),
    .ZN(_16635_)
  );
  AND2_X1 _52046_ (
    .A1(\cpuregs[7] [29]),
    .A2(_12651_),
    .ZN(_16636_)
  );
  INV_X1 _52047_ (
    .A(_16636_),
    .ZN(_16637_)
  );
  AND2_X1 _52048_ (
    .A1(_16635_),
    .A2(_16637_),
    .ZN(_16638_)
  );
  INV_X1 _52049_ (
    .A(_16638_),
    .ZN(_01238_)
  );
  AND2_X1 _52050_ (
    .A1(_12650_),
    .A2(_13319_),
    .ZN(_16639_)
  );
  INV_X1 _52051_ (
    .A(_16639_),
    .ZN(_16640_)
  );
  AND2_X1 _52052_ (
    .A1(\cpuregs[7] [30]),
    .A2(_12651_),
    .ZN(_16641_)
  );
  INV_X1 _52053_ (
    .A(_16641_),
    .ZN(_16642_)
  );
  AND2_X1 _52054_ (
    .A1(_16640_),
    .A2(_16642_),
    .ZN(_16643_)
  );
  INV_X1 _52055_ (
    .A(_16643_),
    .ZN(_01239_)
  );
  AND2_X1 _52056_ (
    .A1(_12658_),
    .A2(_12874_),
    .ZN(_16644_)
  );
  INV_X1 _52057_ (
    .A(_16644_),
    .ZN(_16645_)
  );
  AND2_X1 _52058_ (
    .A1(\cpuregs[6] [0]),
    .A2(_12659_),
    .ZN(_16646_)
  );
  INV_X1 _52059_ (
    .A(_16646_),
    .ZN(_16647_)
  );
  AND2_X1 _52060_ (
    .A1(_16645_),
    .A2(_16647_),
    .ZN(_16648_)
  );
  INV_X1 _52061_ (
    .A(_16648_),
    .ZN(_01240_)
  );
  AND2_X1 _52062_ (
    .A1(_12658_),
    .A2(_12886_),
    .ZN(_16649_)
  );
  INV_X1 _52063_ (
    .A(_16649_),
    .ZN(_16650_)
  );
  AND2_X1 _52064_ (
    .A1(\cpuregs[6] [1]),
    .A2(_12659_),
    .ZN(_16651_)
  );
  INV_X1 _52065_ (
    .A(_16651_),
    .ZN(_16652_)
  );
  AND2_X1 _52066_ (
    .A1(_16650_),
    .A2(_16652_),
    .ZN(_16653_)
  );
  INV_X1 _52067_ (
    .A(_16653_),
    .ZN(_01241_)
  );
  AND2_X1 _52068_ (
    .A1(_12658_),
    .A2(_12900_),
    .ZN(_16654_)
  );
  INV_X1 _52069_ (
    .A(_16654_),
    .ZN(_16655_)
  );
  AND2_X1 _52070_ (
    .A1(\cpuregs[6] [2]),
    .A2(_12659_),
    .ZN(_16656_)
  );
  INV_X1 _52071_ (
    .A(_16656_),
    .ZN(_16657_)
  );
  AND2_X1 _52072_ (
    .A1(_16655_),
    .A2(_16657_),
    .ZN(_16658_)
  );
  INV_X1 _52073_ (
    .A(_16658_),
    .ZN(_01242_)
  );
  AND2_X1 _52074_ (
    .A1(_12658_),
    .A2(_12913_),
    .ZN(_16659_)
  );
  INV_X1 _52075_ (
    .A(_16659_),
    .ZN(_16660_)
  );
  AND2_X1 _52076_ (
    .A1(\cpuregs[6] [3]),
    .A2(_12659_),
    .ZN(_16661_)
  );
  INV_X1 _52077_ (
    .A(_16661_),
    .ZN(_16662_)
  );
  AND2_X1 _52078_ (
    .A1(_16660_),
    .A2(_16662_),
    .ZN(_16663_)
  );
  INV_X1 _52079_ (
    .A(_16663_),
    .ZN(_01243_)
  );
  AND2_X1 _52080_ (
    .A1(\cpuregs[6] [4]),
    .A2(_12659_),
    .ZN(_16664_)
  );
  INV_X1 _52081_ (
    .A(_16664_),
    .ZN(_16665_)
  );
  AND2_X1 _52082_ (
    .A1(_12658_),
    .A2(_12928_),
    .ZN(_16666_)
  );
  INV_X1 _52083_ (
    .A(_16666_),
    .ZN(_16667_)
  );
  AND2_X1 _52084_ (
    .A1(_16665_),
    .A2(_16667_),
    .ZN(_16668_)
  );
  INV_X1 _52085_ (
    .A(_16668_),
    .ZN(_01244_)
  );
  AND2_X1 _52086_ (
    .A1(_12658_),
    .A2(_12943_),
    .ZN(_16669_)
  );
  INV_X1 _52087_ (
    .A(_16669_),
    .ZN(_16670_)
  );
  AND2_X1 _52088_ (
    .A1(\cpuregs[6] [5]),
    .A2(_12659_),
    .ZN(_16671_)
  );
  INV_X1 _52089_ (
    .A(_16671_),
    .ZN(_16672_)
  );
  AND2_X1 _52090_ (
    .A1(_16670_),
    .A2(_16672_),
    .ZN(_16673_)
  );
  INV_X1 _52091_ (
    .A(_16673_),
    .ZN(_01245_)
  );
  AND2_X1 _52092_ (
    .A1(_12658_),
    .A2(_12958_),
    .ZN(_16674_)
  );
  INV_X1 _52093_ (
    .A(_16674_),
    .ZN(_16675_)
  );
  AND2_X1 _52094_ (
    .A1(\cpuregs[6] [6]),
    .A2(_12659_),
    .ZN(_16676_)
  );
  INV_X1 _52095_ (
    .A(_16676_),
    .ZN(_16677_)
  );
  AND2_X1 _52096_ (
    .A1(_16675_),
    .A2(_16677_),
    .ZN(_16678_)
  );
  INV_X1 _52097_ (
    .A(_16678_),
    .ZN(_01246_)
  );
  AND2_X1 _52098_ (
    .A1(_12658_),
    .A2(_12973_),
    .ZN(_16679_)
  );
  INV_X1 _52099_ (
    .A(_16679_),
    .ZN(_16680_)
  );
  AND2_X1 _52100_ (
    .A1(\cpuregs[6] [7]),
    .A2(_12659_),
    .ZN(_16681_)
  );
  INV_X1 _52101_ (
    .A(_16681_),
    .ZN(_16682_)
  );
  AND2_X1 _52102_ (
    .A1(_16680_),
    .A2(_16682_),
    .ZN(_16683_)
  );
  INV_X1 _52103_ (
    .A(_16683_),
    .ZN(_01247_)
  );
  AND2_X1 _52104_ (
    .A1(_12658_),
    .A2(_12988_),
    .ZN(_16684_)
  );
  INV_X1 _52105_ (
    .A(_16684_),
    .ZN(_16685_)
  );
  AND2_X1 _52106_ (
    .A1(\cpuregs[6] [8]),
    .A2(_12659_),
    .ZN(_16686_)
  );
  INV_X1 _52107_ (
    .A(_16686_),
    .ZN(_16687_)
  );
  AND2_X1 _52108_ (
    .A1(_16685_),
    .A2(_16687_),
    .ZN(_16688_)
  );
  INV_X1 _52109_ (
    .A(_16688_),
    .ZN(_01248_)
  );
  AND2_X1 _52110_ (
    .A1(_12658_),
    .A2(_13003_),
    .ZN(_16689_)
  );
  INV_X1 _52111_ (
    .A(_16689_),
    .ZN(_16690_)
  );
  AND2_X1 _52112_ (
    .A1(\cpuregs[6] [9]),
    .A2(_12659_),
    .ZN(_16691_)
  );
  INV_X1 _52113_ (
    .A(_16691_),
    .ZN(_16692_)
  );
  AND2_X1 _52114_ (
    .A1(_16690_),
    .A2(_16692_),
    .ZN(_16693_)
  );
  INV_X1 _52115_ (
    .A(_16693_),
    .ZN(_01249_)
  );
  AND2_X1 _52116_ (
    .A1(_12658_),
    .A2(_13018_),
    .ZN(_16694_)
  );
  INV_X1 _52117_ (
    .A(_16694_),
    .ZN(_16695_)
  );
  AND2_X1 _52118_ (
    .A1(\cpuregs[6] [10]),
    .A2(_12659_),
    .ZN(_16696_)
  );
  INV_X1 _52119_ (
    .A(_16696_),
    .ZN(_16697_)
  );
  AND2_X1 _52120_ (
    .A1(_16695_),
    .A2(_16697_),
    .ZN(_16698_)
  );
  INV_X1 _52121_ (
    .A(_16698_),
    .ZN(_01250_)
  );
  AND2_X1 _52122_ (
    .A1(_12658_),
    .A2(_13033_),
    .ZN(_16699_)
  );
  INV_X1 _52123_ (
    .A(_16699_),
    .ZN(_16700_)
  );
  AND2_X1 _52124_ (
    .A1(\cpuregs[6] [11]),
    .A2(_12659_),
    .ZN(_16701_)
  );
  INV_X1 _52125_ (
    .A(_16701_),
    .ZN(_16702_)
  );
  AND2_X1 _52126_ (
    .A1(_16700_),
    .A2(_16702_),
    .ZN(_16703_)
  );
  INV_X1 _52127_ (
    .A(_16703_),
    .ZN(_01251_)
  );
  AND2_X1 _52128_ (
    .A1(_12658_),
    .A2(_13048_),
    .ZN(_16704_)
  );
  INV_X1 _52129_ (
    .A(_16704_),
    .ZN(_16705_)
  );
  AND2_X1 _52130_ (
    .A1(\cpuregs[6] [12]),
    .A2(_12659_),
    .ZN(_16706_)
  );
  INV_X1 _52131_ (
    .A(_16706_),
    .ZN(_16707_)
  );
  AND2_X1 _52132_ (
    .A1(_16705_),
    .A2(_16707_),
    .ZN(_16708_)
  );
  INV_X1 _52133_ (
    .A(_16708_),
    .ZN(_01252_)
  );
  AND2_X1 _52134_ (
    .A1(_12658_),
    .A2(_13063_),
    .ZN(_16709_)
  );
  INV_X1 _52135_ (
    .A(_16709_),
    .ZN(_16710_)
  );
  AND2_X1 _52136_ (
    .A1(\cpuregs[6] [13]),
    .A2(_12659_),
    .ZN(_16711_)
  );
  INV_X1 _52137_ (
    .A(_16711_),
    .ZN(_16712_)
  );
  AND2_X1 _52138_ (
    .A1(_16710_),
    .A2(_16712_),
    .ZN(_16713_)
  );
  INV_X1 _52139_ (
    .A(_16713_),
    .ZN(_01253_)
  );
  AND2_X1 _52140_ (
    .A1(\cpuregs[6] [14]),
    .A2(_12659_),
    .ZN(_16714_)
  );
  INV_X1 _52141_ (
    .A(_16714_),
    .ZN(_16715_)
  );
  AND2_X1 _52142_ (
    .A1(_12658_),
    .A2(_13078_),
    .ZN(_16716_)
  );
  INV_X1 _52143_ (
    .A(_16716_),
    .ZN(_16717_)
  );
  AND2_X1 _52144_ (
    .A1(_16715_),
    .A2(_16717_),
    .ZN(_16718_)
  );
  INV_X1 _52145_ (
    .A(_16718_),
    .ZN(_01254_)
  );
  AND2_X1 _52146_ (
    .A1(_12658_),
    .A2(_13093_),
    .ZN(_16719_)
  );
  INV_X1 _52147_ (
    .A(_16719_),
    .ZN(_16720_)
  );
  AND2_X1 _52148_ (
    .A1(\cpuregs[6] [15]),
    .A2(_12659_),
    .ZN(_16721_)
  );
  INV_X1 _52149_ (
    .A(_16721_),
    .ZN(_16722_)
  );
  AND2_X1 _52150_ (
    .A1(_16720_),
    .A2(_16722_),
    .ZN(_16723_)
  );
  INV_X1 _52151_ (
    .A(_16723_),
    .ZN(_01255_)
  );
  AND2_X1 _52152_ (
    .A1(_12658_),
    .A2(_13108_),
    .ZN(_16724_)
  );
  INV_X1 _52153_ (
    .A(_16724_),
    .ZN(_16725_)
  );
  AND2_X1 _52154_ (
    .A1(\cpuregs[6] [16]),
    .A2(_12659_),
    .ZN(_16726_)
  );
  INV_X1 _52155_ (
    .A(_16726_),
    .ZN(_16727_)
  );
  AND2_X1 _52156_ (
    .A1(_16725_),
    .A2(_16727_),
    .ZN(_16728_)
  );
  INV_X1 _52157_ (
    .A(_16728_),
    .ZN(_01256_)
  );
  AND2_X1 _52158_ (
    .A1(_12658_),
    .A2(_13123_),
    .ZN(_16729_)
  );
  INV_X1 _52159_ (
    .A(_16729_),
    .ZN(_16730_)
  );
  AND2_X1 _52160_ (
    .A1(\cpuregs[6] [17]),
    .A2(_12659_),
    .ZN(_16731_)
  );
  INV_X1 _52161_ (
    .A(_16731_),
    .ZN(_16732_)
  );
  AND2_X1 _52162_ (
    .A1(_16730_),
    .A2(_16732_),
    .ZN(_16733_)
  );
  INV_X1 _52163_ (
    .A(_16733_),
    .ZN(_01257_)
  );
  AND2_X1 _52164_ (
    .A1(_12658_),
    .A2(_13139_),
    .ZN(_16734_)
  );
  INV_X1 _52165_ (
    .A(_16734_),
    .ZN(_16735_)
  );
  AND2_X1 _52166_ (
    .A1(\cpuregs[6] [18]),
    .A2(_12659_),
    .ZN(_16736_)
  );
  INV_X1 _52167_ (
    .A(_16736_),
    .ZN(_16737_)
  );
  AND2_X1 _52168_ (
    .A1(_16735_),
    .A2(_16737_),
    .ZN(_16738_)
  );
  INV_X1 _52169_ (
    .A(_16738_),
    .ZN(_01258_)
  );
  AND2_X1 _52170_ (
    .A1(_12658_),
    .A2(_13154_),
    .ZN(_16739_)
  );
  INV_X1 _52171_ (
    .A(_16739_),
    .ZN(_16740_)
  );
  AND2_X1 _52172_ (
    .A1(\cpuregs[6] [19]),
    .A2(_12659_),
    .ZN(_16741_)
  );
  INV_X1 _52173_ (
    .A(_16741_),
    .ZN(_16742_)
  );
  AND2_X1 _52174_ (
    .A1(_16740_),
    .A2(_16742_),
    .ZN(_16743_)
  );
  INV_X1 _52175_ (
    .A(_16743_),
    .ZN(_01259_)
  );
  AND2_X1 _52176_ (
    .A1(_12658_),
    .A2(_13169_),
    .ZN(_16744_)
  );
  INV_X1 _52177_ (
    .A(_16744_),
    .ZN(_16745_)
  );
  AND2_X1 _52178_ (
    .A1(\cpuregs[6] [20]),
    .A2(_12659_),
    .ZN(_16746_)
  );
  INV_X1 _52179_ (
    .A(_16746_),
    .ZN(_16747_)
  );
  AND2_X1 _52180_ (
    .A1(_16745_),
    .A2(_16747_),
    .ZN(_16748_)
  );
  INV_X1 _52181_ (
    .A(_16748_),
    .ZN(_01260_)
  );
  AND2_X1 _52182_ (
    .A1(_12658_),
    .A2(_13184_),
    .ZN(_16749_)
  );
  INV_X1 _52183_ (
    .A(_16749_),
    .ZN(_16750_)
  );
  AND2_X1 _52184_ (
    .A1(\cpuregs[6] [21]),
    .A2(_12659_),
    .ZN(_16751_)
  );
  INV_X1 _52185_ (
    .A(_16751_),
    .ZN(_16752_)
  );
  AND2_X1 _52186_ (
    .A1(_16750_),
    .A2(_16752_),
    .ZN(_16753_)
  );
  INV_X1 _52187_ (
    .A(_16753_),
    .ZN(_01261_)
  );
  AND2_X1 _52188_ (
    .A1(_12658_),
    .A2(_13199_),
    .ZN(_16754_)
  );
  INV_X1 _52189_ (
    .A(_16754_),
    .ZN(_16755_)
  );
  AND2_X1 _52190_ (
    .A1(\cpuregs[6] [22]),
    .A2(_12659_),
    .ZN(_16756_)
  );
  INV_X1 _52191_ (
    .A(_16756_),
    .ZN(_16757_)
  );
  AND2_X1 _52192_ (
    .A1(_16755_),
    .A2(_16757_),
    .ZN(_16758_)
  );
  INV_X1 _52193_ (
    .A(_16758_),
    .ZN(_01262_)
  );
  AND2_X1 _52194_ (
    .A1(_12658_),
    .A2(_13214_),
    .ZN(_16759_)
  );
  INV_X1 _52195_ (
    .A(_16759_),
    .ZN(_16760_)
  );
  AND2_X1 _52196_ (
    .A1(\cpuregs[6] [23]),
    .A2(_12659_),
    .ZN(_16761_)
  );
  INV_X1 _52197_ (
    .A(_16761_),
    .ZN(_16762_)
  );
  AND2_X1 _52198_ (
    .A1(_16760_),
    .A2(_16762_),
    .ZN(_16763_)
  );
  INV_X1 _52199_ (
    .A(_16763_),
    .ZN(_01263_)
  );
  AND2_X1 _52200_ (
    .A1(_12658_),
    .A2(_13229_),
    .ZN(_16764_)
  );
  INV_X1 _52201_ (
    .A(_16764_),
    .ZN(_16765_)
  );
  AND2_X1 _52202_ (
    .A1(\cpuregs[6] [24]),
    .A2(_12659_),
    .ZN(_16766_)
  );
  INV_X1 _52203_ (
    .A(_16766_),
    .ZN(_16767_)
  );
  AND2_X1 _52204_ (
    .A1(_16765_),
    .A2(_16767_),
    .ZN(_16768_)
  );
  INV_X1 _52205_ (
    .A(_16768_),
    .ZN(_01264_)
  );
  AND2_X1 _52206_ (
    .A1(_12658_),
    .A2(_13244_),
    .ZN(_16769_)
  );
  INV_X1 _52207_ (
    .A(_16769_),
    .ZN(_16770_)
  );
  AND2_X1 _52208_ (
    .A1(\cpuregs[6] [25]),
    .A2(_12659_),
    .ZN(_16771_)
  );
  INV_X1 _52209_ (
    .A(_16771_),
    .ZN(_16772_)
  );
  AND2_X1 _52210_ (
    .A1(_16770_),
    .A2(_16772_),
    .ZN(_16773_)
  );
  INV_X1 _52211_ (
    .A(_16773_),
    .ZN(_01265_)
  );
  AND2_X1 _52212_ (
    .A1(_12658_),
    .A2(_13259_),
    .ZN(_16774_)
  );
  INV_X1 _52213_ (
    .A(_16774_),
    .ZN(_16775_)
  );
  AND2_X1 _52214_ (
    .A1(\cpuregs[6] [26]),
    .A2(_12659_),
    .ZN(_16776_)
  );
  INV_X1 _52215_ (
    .A(_16776_),
    .ZN(_16777_)
  );
  AND2_X1 _52216_ (
    .A1(_16775_),
    .A2(_16777_),
    .ZN(_16778_)
  );
  INV_X1 _52217_ (
    .A(_16778_),
    .ZN(_01266_)
  );
  AND2_X1 _52218_ (
    .A1(_12658_),
    .A2(_13274_),
    .ZN(_16779_)
  );
  INV_X1 _52219_ (
    .A(_16779_),
    .ZN(_16780_)
  );
  AND2_X1 _52220_ (
    .A1(\cpuregs[6] [27]),
    .A2(_12659_),
    .ZN(_16781_)
  );
  INV_X1 _52221_ (
    .A(_16781_),
    .ZN(_16782_)
  );
  AND2_X1 _52222_ (
    .A1(_16780_),
    .A2(_16782_),
    .ZN(_16783_)
  );
  INV_X1 _52223_ (
    .A(_16783_),
    .ZN(_01267_)
  );
  AND2_X1 _52224_ (
    .A1(_12658_),
    .A2(_13289_),
    .ZN(_16784_)
  );
  INV_X1 _52225_ (
    .A(_16784_),
    .ZN(_16785_)
  );
  AND2_X1 _52226_ (
    .A1(\cpuregs[6] [28]),
    .A2(_12659_),
    .ZN(_16786_)
  );
  INV_X1 _52227_ (
    .A(_16786_),
    .ZN(_16787_)
  );
  AND2_X1 _52228_ (
    .A1(_16785_),
    .A2(_16787_),
    .ZN(_16788_)
  );
  INV_X1 _52229_ (
    .A(_16788_),
    .ZN(_01268_)
  );
  AND2_X1 _52230_ (
    .A1(_12658_),
    .A2(_13304_),
    .ZN(_16789_)
  );
  INV_X1 _52231_ (
    .A(_16789_),
    .ZN(_16790_)
  );
  AND2_X1 _52232_ (
    .A1(\cpuregs[6] [29]),
    .A2(_12659_),
    .ZN(_16791_)
  );
  INV_X1 _52233_ (
    .A(_16791_),
    .ZN(_16792_)
  );
  AND2_X1 _52234_ (
    .A1(_16790_),
    .A2(_16792_),
    .ZN(_16793_)
  );
  INV_X1 _52235_ (
    .A(_16793_),
    .ZN(_01269_)
  );
  AND2_X1 _52236_ (
    .A1(_12658_),
    .A2(_13319_),
    .ZN(_16794_)
  );
  INV_X1 _52237_ (
    .A(_16794_),
    .ZN(_16795_)
  );
  AND2_X1 _52238_ (
    .A1(\cpuregs[6] [30]),
    .A2(_12659_),
    .ZN(_16796_)
  );
  INV_X1 _52239_ (
    .A(_16796_),
    .ZN(_16797_)
  );
  AND2_X1 _52240_ (
    .A1(_16795_),
    .A2(_16797_),
    .ZN(_16798_)
  );
  INV_X1 _52241_ (
    .A(_16798_),
    .ZN(_01270_)
  );
  AND2_X1 _52242_ (
    .A1(_12739_),
    .A2(_12874_),
    .ZN(_16799_)
  );
  INV_X1 _52243_ (
    .A(_16799_),
    .ZN(_16800_)
  );
  AND2_X1 _52244_ (
    .A1(\cpuregs[25] [0]),
    .A2(_12740_),
    .ZN(_16801_)
  );
  INV_X1 _52245_ (
    .A(_16801_),
    .ZN(_16802_)
  );
  AND2_X1 _52246_ (
    .A1(_16800_),
    .A2(_16802_),
    .ZN(_16803_)
  );
  INV_X1 _52247_ (
    .A(_16803_),
    .ZN(_01271_)
  );
  AND2_X1 _52248_ (
    .A1(_12739_),
    .A2(_12886_),
    .ZN(_16804_)
  );
  INV_X1 _52249_ (
    .A(_16804_),
    .ZN(_16805_)
  );
  AND2_X1 _52250_ (
    .A1(\cpuregs[25] [1]),
    .A2(_12740_),
    .ZN(_16806_)
  );
  INV_X1 _52251_ (
    .A(_16806_),
    .ZN(_16807_)
  );
  AND2_X1 _52252_ (
    .A1(_16805_),
    .A2(_16807_),
    .ZN(_16808_)
  );
  INV_X1 _52253_ (
    .A(_16808_),
    .ZN(_01272_)
  );
  AND2_X1 _52254_ (
    .A1(\cpuregs[25] [2]),
    .A2(_12740_),
    .ZN(_16809_)
  );
  INV_X1 _52255_ (
    .A(_16809_),
    .ZN(_16810_)
  );
  AND2_X1 _52256_ (
    .A1(_12739_),
    .A2(_12900_),
    .ZN(_16811_)
  );
  INV_X1 _52257_ (
    .A(_16811_),
    .ZN(_16812_)
  );
  AND2_X1 _52258_ (
    .A1(_16810_),
    .A2(_16812_),
    .ZN(_16813_)
  );
  INV_X1 _52259_ (
    .A(_16813_),
    .ZN(_01273_)
  );
  AND2_X1 _52260_ (
    .A1(_12739_),
    .A2(_12913_),
    .ZN(_16814_)
  );
  INV_X1 _52261_ (
    .A(_16814_),
    .ZN(_16815_)
  );
  AND2_X1 _52262_ (
    .A1(\cpuregs[25] [3]),
    .A2(_12740_),
    .ZN(_16816_)
  );
  INV_X1 _52263_ (
    .A(_16816_),
    .ZN(_16817_)
  );
  AND2_X1 _52264_ (
    .A1(_16815_),
    .A2(_16817_),
    .ZN(_16818_)
  );
  INV_X1 _52265_ (
    .A(_16818_),
    .ZN(_01274_)
  );
  AND2_X1 _52266_ (
    .A1(\cpuregs[25] [4]),
    .A2(_12740_),
    .ZN(_16819_)
  );
  INV_X1 _52267_ (
    .A(_16819_),
    .ZN(_16820_)
  );
  AND2_X1 _52268_ (
    .A1(_12739_),
    .A2(_12928_),
    .ZN(_16821_)
  );
  INV_X1 _52269_ (
    .A(_16821_),
    .ZN(_16822_)
  );
  AND2_X1 _52270_ (
    .A1(_16820_),
    .A2(_16822_),
    .ZN(_16823_)
  );
  INV_X1 _52271_ (
    .A(_16823_),
    .ZN(_01275_)
  );
  AND2_X1 _52272_ (
    .A1(_12739_),
    .A2(_12943_),
    .ZN(_16824_)
  );
  INV_X1 _52273_ (
    .A(_16824_),
    .ZN(_16825_)
  );
  AND2_X1 _52274_ (
    .A1(\cpuregs[25] [5]),
    .A2(_12740_),
    .ZN(_16826_)
  );
  INV_X1 _52275_ (
    .A(_16826_),
    .ZN(_16827_)
  );
  AND2_X1 _52276_ (
    .A1(_16825_),
    .A2(_16827_),
    .ZN(_16828_)
  );
  INV_X1 _52277_ (
    .A(_16828_),
    .ZN(_01276_)
  );
  AND2_X1 _52278_ (
    .A1(_12739_),
    .A2(_12958_),
    .ZN(_16829_)
  );
  INV_X1 _52279_ (
    .A(_16829_),
    .ZN(_16830_)
  );
  AND2_X1 _52280_ (
    .A1(\cpuregs[25] [6]),
    .A2(_12740_),
    .ZN(_16831_)
  );
  INV_X1 _52281_ (
    .A(_16831_),
    .ZN(_16832_)
  );
  AND2_X1 _52282_ (
    .A1(_16830_),
    .A2(_16832_),
    .ZN(_16833_)
  );
  INV_X1 _52283_ (
    .A(_16833_),
    .ZN(_01277_)
  );
  AND2_X1 _52284_ (
    .A1(_12739_),
    .A2(_12973_),
    .ZN(_16834_)
  );
  INV_X1 _52285_ (
    .A(_16834_),
    .ZN(_16835_)
  );
  AND2_X1 _52286_ (
    .A1(\cpuregs[25] [7]),
    .A2(_12740_),
    .ZN(_16836_)
  );
  INV_X1 _52287_ (
    .A(_16836_),
    .ZN(_16837_)
  );
  AND2_X1 _52288_ (
    .A1(_16835_),
    .A2(_16837_),
    .ZN(_16838_)
  );
  INV_X1 _52289_ (
    .A(_16838_),
    .ZN(_01278_)
  );
  AND2_X1 _52290_ (
    .A1(_12739_),
    .A2(_12988_),
    .ZN(_16839_)
  );
  INV_X1 _52291_ (
    .A(_16839_),
    .ZN(_16840_)
  );
  AND2_X1 _52292_ (
    .A1(\cpuregs[25] [8]),
    .A2(_12740_),
    .ZN(_16841_)
  );
  INV_X1 _52293_ (
    .A(_16841_),
    .ZN(_16842_)
  );
  AND2_X1 _52294_ (
    .A1(_16840_),
    .A2(_16842_),
    .ZN(_16843_)
  );
  INV_X1 _52295_ (
    .A(_16843_),
    .ZN(_01279_)
  );
  AND2_X1 _52296_ (
    .A1(_12739_),
    .A2(_13003_),
    .ZN(_16844_)
  );
  INV_X1 _52297_ (
    .A(_16844_),
    .ZN(_16845_)
  );
  AND2_X1 _52298_ (
    .A1(\cpuregs[25] [9]),
    .A2(_12740_),
    .ZN(_16846_)
  );
  INV_X1 _52299_ (
    .A(_16846_),
    .ZN(_16847_)
  );
  AND2_X1 _52300_ (
    .A1(_16845_),
    .A2(_16847_),
    .ZN(_16848_)
  );
  INV_X1 _52301_ (
    .A(_16848_),
    .ZN(_01280_)
  );
  AND2_X1 _52302_ (
    .A1(_12739_),
    .A2(_13018_),
    .ZN(_16849_)
  );
  INV_X1 _52303_ (
    .A(_16849_),
    .ZN(_16850_)
  );
  AND2_X1 _52304_ (
    .A1(\cpuregs[25] [10]),
    .A2(_12740_),
    .ZN(_16851_)
  );
  INV_X1 _52305_ (
    .A(_16851_),
    .ZN(_16852_)
  );
  AND2_X1 _52306_ (
    .A1(_16850_),
    .A2(_16852_),
    .ZN(_16853_)
  );
  INV_X1 _52307_ (
    .A(_16853_),
    .ZN(_01281_)
  );
  AND2_X1 _52308_ (
    .A1(_12739_),
    .A2(_13033_),
    .ZN(_16854_)
  );
  INV_X1 _52309_ (
    .A(_16854_),
    .ZN(_16855_)
  );
  AND2_X1 _52310_ (
    .A1(\cpuregs[25] [11]),
    .A2(_12740_),
    .ZN(_16856_)
  );
  INV_X1 _52311_ (
    .A(_16856_),
    .ZN(_16857_)
  );
  AND2_X1 _52312_ (
    .A1(_16855_),
    .A2(_16857_),
    .ZN(_16858_)
  );
  INV_X1 _52313_ (
    .A(_16858_),
    .ZN(_01282_)
  );
  AND2_X1 _52314_ (
    .A1(_12739_),
    .A2(_13048_),
    .ZN(_16859_)
  );
  INV_X1 _52315_ (
    .A(_16859_),
    .ZN(_16860_)
  );
  AND2_X1 _52316_ (
    .A1(\cpuregs[25] [12]),
    .A2(_12740_),
    .ZN(_16861_)
  );
  INV_X1 _52317_ (
    .A(_16861_),
    .ZN(_16862_)
  );
  AND2_X1 _52318_ (
    .A1(_16860_),
    .A2(_16862_),
    .ZN(_16863_)
  );
  INV_X1 _52319_ (
    .A(_16863_),
    .ZN(_01283_)
  );
  AND2_X1 _52320_ (
    .A1(_12739_),
    .A2(_13063_),
    .ZN(_16864_)
  );
  INV_X1 _52321_ (
    .A(_16864_),
    .ZN(_16865_)
  );
  AND2_X1 _52322_ (
    .A1(\cpuregs[25] [13]),
    .A2(_12740_),
    .ZN(_16866_)
  );
  INV_X1 _52323_ (
    .A(_16866_),
    .ZN(_16867_)
  );
  AND2_X1 _52324_ (
    .A1(_16865_),
    .A2(_16867_),
    .ZN(_16868_)
  );
  INV_X1 _52325_ (
    .A(_16868_),
    .ZN(_01284_)
  );
  AND2_X1 _52326_ (
    .A1(_12739_),
    .A2(_13078_),
    .ZN(_16869_)
  );
  INV_X1 _52327_ (
    .A(_16869_),
    .ZN(_16870_)
  );
  AND2_X1 _52328_ (
    .A1(\cpuregs[25] [14]),
    .A2(_12740_),
    .ZN(_16871_)
  );
  INV_X1 _52329_ (
    .A(_16871_),
    .ZN(_16872_)
  );
  AND2_X1 _52330_ (
    .A1(_16870_),
    .A2(_16872_),
    .ZN(_16873_)
  );
  INV_X1 _52331_ (
    .A(_16873_),
    .ZN(_01285_)
  );
  AND2_X1 _52332_ (
    .A1(_12739_),
    .A2(_13093_),
    .ZN(_16874_)
  );
  INV_X1 _52333_ (
    .A(_16874_),
    .ZN(_16875_)
  );
  AND2_X1 _52334_ (
    .A1(\cpuregs[25] [15]),
    .A2(_12740_),
    .ZN(_16876_)
  );
  INV_X1 _52335_ (
    .A(_16876_),
    .ZN(_16877_)
  );
  AND2_X1 _52336_ (
    .A1(_16875_),
    .A2(_16877_),
    .ZN(_16878_)
  );
  INV_X1 _52337_ (
    .A(_16878_),
    .ZN(_01286_)
  );
  AND2_X1 _52338_ (
    .A1(_12739_),
    .A2(_13108_),
    .ZN(_16879_)
  );
  INV_X1 _52339_ (
    .A(_16879_),
    .ZN(_16880_)
  );
  AND2_X1 _52340_ (
    .A1(\cpuregs[25] [16]),
    .A2(_12740_),
    .ZN(_16881_)
  );
  INV_X1 _52341_ (
    .A(_16881_),
    .ZN(_16882_)
  );
  AND2_X1 _52342_ (
    .A1(_16880_),
    .A2(_16882_),
    .ZN(_16883_)
  );
  INV_X1 _52343_ (
    .A(_16883_),
    .ZN(_01287_)
  );
  AND2_X1 _52344_ (
    .A1(_12739_),
    .A2(_13123_),
    .ZN(_16884_)
  );
  INV_X1 _52345_ (
    .A(_16884_),
    .ZN(_16885_)
  );
  AND2_X1 _52346_ (
    .A1(\cpuregs[25] [17]),
    .A2(_12740_),
    .ZN(_16886_)
  );
  INV_X1 _52347_ (
    .A(_16886_),
    .ZN(_16887_)
  );
  AND2_X1 _52348_ (
    .A1(_16885_),
    .A2(_16887_),
    .ZN(_16888_)
  );
  INV_X1 _52349_ (
    .A(_16888_),
    .ZN(_01288_)
  );
  AND2_X1 _52350_ (
    .A1(_12739_),
    .A2(_13139_),
    .ZN(_16889_)
  );
  INV_X1 _52351_ (
    .A(_16889_),
    .ZN(_16890_)
  );
  AND2_X1 _52352_ (
    .A1(\cpuregs[25] [18]),
    .A2(_12740_),
    .ZN(_16891_)
  );
  INV_X1 _52353_ (
    .A(_16891_),
    .ZN(_16892_)
  );
  AND2_X1 _52354_ (
    .A1(_16890_),
    .A2(_16892_),
    .ZN(_16893_)
  );
  INV_X1 _52355_ (
    .A(_16893_),
    .ZN(_01289_)
  );
  AND2_X1 _52356_ (
    .A1(_12739_),
    .A2(_13154_),
    .ZN(_16894_)
  );
  INV_X1 _52357_ (
    .A(_16894_),
    .ZN(_16895_)
  );
  AND2_X1 _52358_ (
    .A1(\cpuregs[25] [19]),
    .A2(_12740_),
    .ZN(_16896_)
  );
  INV_X1 _52359_ (
    .A(_16896_),
    .ZN(_16897_)
  );
  AND2_X1 _52360_ (
    .A1(_16895_),
    .A2(_16897_),
    .ZN(_16898_)
  );
  INV_X1 _52361_ (
    .A(_16898_),
    .ZN(_01290_)
  );
  AND2_X1 _52362_ (
    .A1(_12739_),
    .A2(_13169_),
    .ZN(_16899_)
  );
  INV_X1 _52363_ (
    .A(_16899_),
    .ZN(_16900_)
  );
  AND2_X1 _52364_ (
    .A1(\cpuregs[25] [20]),
    .A2(_12740_),
    .ZN(_16901_)
  );
  INV_X1 _52365_ (
    .A(_16901_),
    .ZN(_16902_)
  );
  AND2_X1 _52366_ (
    .A1(_16900_),
    .A2(_16902_),
    .ZN(_16903_)
  );
  INV_X1 _52367_ (
    .A(_16903_),
    .ZN(_01291_)
  );
  AND2_X1 _52368_ (
    .A1(_12739_),
    .A2(_13184_),
    .ZN(_16904_)
  );
  INV_X1 _52369_ (
    .A(_16904_),
    .ZN(_16905_)
  );
  AND2_X1 _52370_ (
    .A1(\cpuregs[25] [21]),
    .A2(_12740_),
    .ZN(_16906_)
  );
  INV_X1 _52371_ (
    .A(_16906_),
    .ZN(_16907_)
  );
  AND2_X1 _52372_ (
    .A1(_16905_),
    .A2(_16907_),
    .ZN(_16908_)
  );
  INV_X1 _52373_ (
    .A(_16908_),
    .ZN(_01292_)
  );
  AND2_X1 _52374_ (
    .A1(_12739_),
    .A2(_13199_),
    .ZN(_16909_)
  );
  INV_X1 _52375_ (
    .A(_16909_),
    .ZN(_16910_)
  );
  AND2_X1 _52376_ (
    .A1(\cpuregs[25] [22]),
    .A2(_12740_),
    .ZN(_16911_)
  );
  INV_X1 _52377_ (
    .A(_16911_),
    .ZN(_16912_)
  );
  AND2_X1 _52378_ (
    .A1(_16910_),
    .A2(_16912_),
    .ZN(_16913_)
  );
  INV_X1 _52379_ (
    .A(_16913_),
    .ZN(_01293_)
  );
  AND2_X1 _52380_ (
    .A1(_12739_),
    .A2(_13214_),
    .ZN(_16914_)
  );
  INV_X1 _52381_ (
    .A(_16914_),
    .ZN(_16915_)
  );
  AND2_X1 _52382_ (
    .A1(\cpuregs[25] [23]),
    .A2(_12740_),
    .ZN(_16916_)
  );
  INV_X1 _52383_ (
    .A(_16916_),
    .ZN(_16917_)
  );
  AND2_X1 _52384_ (
    .A1(_16915_),
    .A2(_16917_),
    .ZN(_16918_)
  );
  INV_X1 _52385_ (
    .A(_16918_),
    .ZN(_01294_)
  );
  AND2_X1 _52386_ (
    .A1(_12739_),
    .A2(_13229_),
    .ZN(_16919_)
  );
  INV_X1 _52387_ (
    .A(_16919_),
    .ZN(_16920_)
  );
  AND2_X1 _52388_ (
    .A1(\cpuregs[25] [24]),
    .A2(_12740_),
    .ZN(_16921_)
  );
  INV_X1 _52389_ (
    .A(_16921_),
    .ZN(_16922_)
  );
  AND2_X1 _52390_ (
    .A1(_16920_),
    .A2(_16922_),
    .ZN(_16923_)
  );
  INV_X1 _52391_ (
    .A(_16923_),
    .ZN(_01295_)
  );
  AND2_X1 _52392_ (
    .A1(_12739_),
    .A2(_13244_),
    .ZN(_16924_)
  );
  INV_X1 _52393_ (
    .A(_16924_),
    .ZN(_16925_)
  );
  AND2_X1 _52394_ (
    .A1(\cpuregs[25] [25]),
    .A2(_12740_),
    .ZN(_16926_)
  );
  INV_X1 _52395_ (
    .A(_16926_),
    .ZN(_16927_)
  );
  AND2_X1 _52396_ (
    .A1(_16925_),
    .A2(_16927_),
    .ZN(_16928_)
  );
  INV_X1 _52397_ (
    .A(_16928_),
    .ZN(_01296_)
  );
  AND2_X1 _52398_ (
    .A1(_12739_),
    .A2(_13259_),
    .ZN(_16929_)
  );
  INV_X1 _52399_ (
    .A(_16929_),
    .ZN(_16930_)
  );
  AND2_X1 _52400_ (
    .A1(\cpuregs[25] [26]),
    .A2(_12740_),
    .ZN(_16931_)
  );
  INV_X1 _52401_ (
    .A(_16931_),
    .ZN(_16932_)
  );
  AND2_X1 _52402_ (
    .A1(_16930_),
    .A2(_16932_),
    .ZN(_16933_)
  );
  INV_X1 _52403_ (
    .A(_16933_),
    .ZN(_01297_)
  );
  AND2_X1 _52404_ (
    .A1(_12739_),
    .A2(_13274_),
    .ZN(_16934_)
  );
  INV_X1 _52405_ (
    .A(_16934_),
    .ZN(_16935_)
  );
  AND2_X1 _52406_ (
    .A1(\cpuregs[25] [27]),
    .A2(_12740_),
    .ZN(_16936_)
  );
  INV_X1 _52407_ (
    .A(_16936_),
    .ZN(_16937_)
  );
  AND2_X1 _52408_ (
    .A1(_16935_),
    .A2(_16937_),
    .ZN(_16938_)
  );
  INV_X1 _52409_ (
    .A(_16938_),
    .ZN(_01298_)
  );
  AND2_X1 _52410_ (
    .A1(_12739_),
    .A2(_13289_),
    .ZN(_16939_)
  );
  INV_X1 _52411_ (
    .A(_16939_),
    .ZN(_16940_)
  );
  AND2_X1 _52412_ (
    .A1(\cpuregs[25] [28]),
    .A2(_12740_),
    .ZN(_16941_)
  );
  INV_X1 _52413_ (
    .A(_16941_),
    .ZN(_16942_)
  );
  AND2_X1 _52414_ (
    .A1(_16940_),
    .A2(_16942_),
    .ZN(_16943_)
  );
  INV_X1 _52415_ (
    .A(_16943_),
    .ZN(_01299_)
  );
  AND2_X1 _52416_ (
    .A1(_12739_),
    .A2(_13304_),
    .ZN(_16944_)
  );
  INV_X1 _52417_ (
    .A(_16944_),
    .ZN(_16945_)
  );
  AND2_X1 _52418_ (
    .A1(\cpuregs[25] [29]),
    .A2(_12740_),
    .ZN(_16946_)
  );
  INV_X1 _52419_ (
    .A(_16946_),
    .ZN(_16947_)
  );
  AND2_X1 _52420_ (
    .A1(_16945_),
    .A2(_16947_),
    .ZN(_16948_)
  );
  INV_X1 _52421_ (
    .A(_16948_),
    .ZN(_01300_)
  );
  AND2_X1 _52422_ (
    .A1(_12739_),
    .A2(_13319_),
    .ZN(_16949_)
  );
  INV_X1 _52423_ (
    .A(_16949_),
    .ZN(_16950_)
  );
  AND2_X1 _52424_ (
    .A1(\cpuregs[25] [30]),
    .A2(_12740_),
    .ZN(_16951_)
  );
  INV_X1 _52425_ (
    .A(_16951_),
    .ZN(_16952_)
  );
  AND2_X1 _52426_ (
    .A1(_16950_),
    .A2(_16952_),
    .ZN(_16953_)
  );
  INV_X1 _52427_ (
    .A(_16953_),
    .ZN(_01301_)
  );
  AND2_X1 _52428_ (
    .A1(_12696_),
    .A2(_12874_),
    .ZN(_16954_)
  );
  INV_X1 _52429_ (
    .A(_16954_),
    .ZN(_16955_)
  );
  AND2_X1 _52430_ (
    .A1(\cpuregs[30] [0]),
    .A2(_12697_),
    .ZN(_16956_)
  );
  INV_X1 _52431_ (
    .A(_16956_),
    .ZN(_16957_)
  );
  AND2_X1 _52432_ (
    .A1(_16955_),
    .A2(_16957_),
    .ZN(_16958_)
  );
  INV_X1 _52433_ (
    .A(_16958_),
    .ZN(_01302_)
  );
  AND2_X1 _52434_ (
    .A1(_12696_),
    .A2(_12886_),
    .ZN(_16959_)
  );
  INV_X1 _52435_ (
    .A(_16959_),
    .ZN(_16960_)
  );
  AND2_X1 _52436_ (
    .A1(\cpuregs[30] [1]),
    .A2(_12697_),
    .ZN(_16961_)
  );
  INV_X1 _52437_ (
    .A(_16961_),
    .ZN(_16962_)
  );
  AND2_X1 _52438_ (
    .A1(_16960_),
    .A2(_16962_),
    .ZN(_16963_)
  );
  INV_X1 _52439_ (
    .A(_16963_),
    .ZN(_01303_)
  );
  AND2_X1 _52440_ (
    .A1(_12696_),
    .A2(_12900_),
    .ZN(_16964_)
  );
  INV_X1 _52441_ (
    .A(_16964_),
    .ZN(_16965_)
  );
  AND2_X1 _52442_ (
    .A1(\cpuregs[30] [2]),
    .A2(_12697_),
    .ZN(_16966_)
  );
  INV_X1 _52443_ (
    .A(_16966_),
    .ZN(_16967_)
  );
  AND2_X1 _52444_ (
    .A1(_16965_),
    .A2(_16967_),
    .ZN(_16968_)
  );
  INV_X1 _52445_ (
    .A(_16968_),
    .ZN(_01304_)
  );
  AND2_X1 _52446_ (
    .A1(_12696_),
    .A2(_12913_),
    .ZN(_16969_)
  );
  INV_X1 _52447_ (
    .A(_16969_),
    .ZN(_16970_)
  );
  AND2_X1 _52448_ (
    .A1(\cpuregs[30] [3]),
    .A2(_12697_),
    .ZN(_16971_)
  );
  INV_X1 _52449_ (
    .A(_16971_),
    .ZN(_16972_)
  );
  AND2_X1 _52450_ (
    .A1(_16970_),
    .A2(_16972_),
    .ZN(_16973_)
  );
  INV_X1 _52451_ (
    .A(_16973_),
    .ZN(_01305_)
  );
  AND2_X1 _52452_ (
    .A1(_12696_),
    .A2(_12928_),
    .ZN(_16974_)
  );
  INV_X1 _52453_ (
    .A(_16974_),
    .ZN(_16975_)
  );
  AND2_X1 _52454_ (
    .A1(\cpuregs[30] [4]),
    .A2(_12697_),
    .ZN(_16976_)
  );
  INV_X1 _52455_ (
    .A(_16976_),
    .ZN(_16977_)
  );
  AND2_X1 _52456_ (
    .A1(_16975_),
    .A2(_16977_),
    .ZN(_16978_)
  );
  INV_X1 _52457_ (
    .A(_16978_),
    .ZN(_01306_)
  );
  AND2_X1 _52458_ (
    .A1(_12696_),
    .A2(_12943_),
    .ZN(_16979_)
  );
  INV_X1 _52459_ (
    .A(_16979_),
    .ZN(_16980_)
  );
  AND2_X1 _52460_ (
    .A1(\cpuregs[30] [5]),
    .A2(_12697_),
    .ZN(_16981_)
  );
  INV_X1 _52461_ (
    .A(_16981_),
    .ZN(_16982_)
  );
  AND2_X1 _52462_ (
    .A1(_16980_),
    .A2(_16982_),
    .ZN(_16983_)
  );
  INV_X1 _52463_ (
    .A(_16983_),
    .ZN(_01307_)
  );
  AND2_X1 _52464_ (
    .A1(_12696_),
    .A2(_12958_),
    .ZN(_16984_)
  );
  INV_X1 _52465_ (
    .A(_16984_),
    .ZN(_16985_)
  );
  AND2_X1 _52466_ (
    .A1(\cpuregs[30] [6]),
    .A2(_12697_),
    .ZN(_16986_)
  );
  INV_X1 _52467_ (
    .A(_16986_),
    .ZN(_16987_)
  );
  AND2_X1 _52468_ (
    .A1(_16985_),
    .A2(_16987_),
    .ZN(_16988_)
  );
  INV_X1 _52469_ (
    .A(_16988_),
    .ZN(_01308_)
  );
  AND2_X1 _52470_ (
    .A1(_12696_),
    .A2(_12973_),
    .ZN(_16989_)
  );
  INV_X1 _52471_ (
    .A(_16989_),
    .ZN(_16990_)
  );
  AND2_X1 _52472_ (
    .A1(\cpuregs[30] [7]),
    .A2(_12697_),
    .ZN(_16991_)
  );
  INV_X1 _52473_ (
    .A(_16991_),
    .ZN(_16992_)
  );
  AND2_X1 _52474_ (
    .A1(_16990_),
    .A2(_16992_),
    .ZN(_16993_)
  );
  INV_X1 _52475_ (
    .A(_16993_),
    .ZN(_01309_)
  );
  AND2_X1 _52476_ (
    .A1(_12696_),
    .A2(_12988_),
    .ZN(_16994_)
  );
  INV_X1 _52477_ (
    .A(_16994_),
    .ZN(_16995_)
  );
  AND2_X1 _52478_ (
    .A1(\cpuregs[30] [8]),
    .A2(_12697_),
    .ZN(_16996_)
  );
  INV_X1 _52479_ (
    .A(_16996_),
    .ZN(_16997_)
  );
  AND2_X1 _52480_ (
    .A1(_16995_),
    .A2(_16997_),
    .ZN(_16998_)
  );
  INV_X1 _52481_ (
    .A(_16998_),
    .ZN(_01310_)
  );
  AND2_X1 _52482_ (
    .A1(_12696_),
    .A2(_13003_),
    .ZN(_16999_)
  );
  INV_X1 _52483_ (
    .A(_16999_),
    .ZN(_17000_)
  );
  AND2_X1 _52484_ (
    .A1(\cpuregs[30] [9]),
    .A2(_12697_),
    .ZN(_17001_)
  );
  INV_X1 _52485_ (
    .A(_17001_),
    .ZN(_17002_)
  );
  AND2_X1 _52486_ (
    .A1(_17000_),
    .A2(_17002_),
    .ZN(_17003_)
  );
  INV_X1 _52487_ (
    .A(_17003_),
    .ZN(_01311_)
  );
  AND2_X1 _52488_ (
    .A1(_12696_),
    .A2(_13018_),
    .ZN(_17004_)
  );
  INV_X1 _52489_ (
    .A(_17004_),
    .ZN(_17005_)
  );
  AND2_X1 _52490_ (
    .A1(\cpuregs[30] [10]),
    .A2(_12697_),
    .ZN(_17006_)
  );
  INV_X1 _52491_ (
    .A(_17006_),
    .ZN(_17007_)
  );
  AND2_X1 _52492_ (
    .A1(_17005_),
    .A2(_17007_),
    .ZN(_17008_)
  );
  INV_X1 _52493_ (
    .A(_17008_),
    .ZN(_01312_)
  );
  AND2_X1 _52494_ (
    .A1(_12696_),
    .A2(_13033_),
    .ZN(_17009_)
  );
  INV_X1 _52495_ (
    .A(_17009_),
    .ZN(_17010_)
  );
  AND2_X1 _52496_ (
    .A1(\cpuregs[30] [11]),
    .A2(_12697_),
    .ZN(_17011_)
  );
  INV_X1 _52497_ (
    .A(_17011_),
    .ZN(_17012_)
  );
  AND2_X1 _52498_ (
    .A1(_17010_),
    .A2(_17012_),
    .ZN(_17013_)
  );
  INV_X1 _52499_ (
    .A(_17013_),
    .ZN(_01313_)
  );
  AND2_X1 _52500_ (
    .A1(_12696_),
    .A2(_13048_),
    .ZN(_17014_)
  );
  INV_X1 _52501_ (
    .A(_17014_),
    .ZN(_17015_)
  );
  AND2_X1 _52502_ (
    .A1(\cpuregs[30] [12]),
    .A2(_12697_),
    .ZN(_17016_)
  );
  INV_X1 _52503_ (
    .A(_17016_),
    .ZN(_17017_)
  );
  AND2_X1 _52504_ (
    .A1(_17015_),
    .A2(_17017_),
    .ZN(_17018_)
  );
  INV_X1 _52505_ (
    .A(_17018_),
    .ZN(_01314_)
  );
  AND2_X1 _52506_ (
    .A1(_12696_),
    .A2(_13063_),
    .ZN(_17019_)
  );
  INV_X1 _52507_ (
    .A(_17019_),
    .ZN(_17020_)
  );
  AND2_X1 _52508_ (
    .A1(\cpuregs[30] [13]),
    .A2(_12697_),
    .ZN(_17021_)
  );
  INV_X1 _52509_ (
    .A(_17021_),
    .ZN(_17022_)
  );
  AND2_X1 _52510_ (
    .A1(_17020_),
    .A2(_17022_),
    .ZN(_17023_)
  );
  INV_X1 _52511_ (
    .A(_17023_),
    .ZN(_01315_)
  );
  AND2_X1 _52512_ (
    .A1(\cpuregs[30] [14]),
    .A2(_12697_),
    .ZN(_17024_)
  );
  INV_X1 _52513_ (
    .A(_17024_),
    .ZN(_17025_)
  );
  AND2_X1 _52514_ (
    .A1(_12696_),
    .A2(_13078_),
    .ZN(_17026_)
  );
  INV_X1 _52515_ (
    .A(_17026_),
    .ZN(_17027_)
  );
  AND2_X1 _52516_ (
    .A1(_17025_),
    .A2(_17027_),
    .ZN(_17028_)
  );
  INV_X1 _52517_ (
    .A(_17028_),
    .ZN(_01316_)
  );
  AND2_X1 _52518_ (
    .A1(_12696_),
    .A2(_13093_),
    .ZN(_17029_)
  );
  INV_X1 _52519_ (
    .A(_17029_),
    .ZN(_17030_)
  );
  AND2_X1 _52520_ (
    .A1(\cpuregs[30] [15]),
    .A2(_12697_),
    .ZN(_17031_)
  );
  INV_X1 _52521_ (
    .A(_17031_),
    .ZN(_17032_)
  );
  AND2_X1 _52522_ (
    .A1(_17030_),
    .A2(_17032_),
    .ZN(_17033_)
  );
  INV_X1 _52523_ (
    .A(_17033_),
    .ZN(_01317_)
  );
  AND2_X1 _52524_ (
    .A1(\cpuregs[30] [16]),
    .A2(_12697_),
    .ZN(_17034_)
  );
  INV_X1 _52525_ (
    .A(_17034_),
    .ZN(_17035_)
  );
  AND2_X1 _52526_ (
    .A1(_12696_),
    .A2(_13108_),
    .ZN(_17036_)
  );
  INV_X1 _52527_ (
    .A(_17036_),
    .ZN(_17037_)
  );
  AND2_X1 _52528_ (
    .A1(_17035_),
    .A2(_17037_),
    .ZN(_17038_)
  );
  INV_X1 _52529_ (
    .A(_17038_),
    .ZN(_01318_)
  );
  AND2_X1 _52530_ (
    .A1(_12696_),
    .A2(_13123_),
    .ZN(_17039_)
  );
  INV_X1 _52531_ (
    .A(_17039_),
    .ZN(_17040_)
  );
  AND2_X1 _52532_ (
    .A1(\cpuregs[30] [17]),
    .A2(_12697_),
    .ZN(_17041_)
  );
  INV_X1 _52533_ (
    .A(_17041_),
    .ZN(_17042_)
  );
  AND2_X1 _52534_ (
    .A1(_17040_),
    .A2(_17042_),
    .ZN(_17043_)
  );
  INV_X1 _52535_ (
    .A(_17043_),
    .ZN(_01319_)
  );
  AND2_X1 _52536_ (
    .A1(_12696_),
    .A2(_13139_),
    .ZN(_17044_)
  );
  INV_X1 _52537_ (
    .A(_17044_),
    .ZN(_17045_)
  );
  AND2_X1 _52538_ (
    .A1(\cpuregs[30] [18]),
    .A2(_12697_),
    .ZN(_17046_)
  );
  INV_X1 _52539_ (
    .A(_17046_),
    .ZN(_17047_)
  );
  AND2_X1 _52540_ (
    .A1(_17045_),
    .A2(_17047_),
    .ZN(_17048_)
  );
  INV_X1 _52541_ (
    .A(_17048_),
    .ZN(_01320_)
  );
  AND2_X1 _52542_ (
    .A1(_12696_),
    .A2(_13154_),
    .ZN(_17049_)
  );
  INV_X1 _52543_ (
    .A(_17049_),
    .ZN(_17050_)
  );
  AND2_X1 _52544_ (
    .A1(\cpuregs[30] [19]),
    .A2(_12697_),
    .ZN(_17051_)
  );
  INV_X1 _52545_ (
    .A(_17051_),
    .ZN(_17052_)
  );
  AND2_X1 _52546_ (
    .A1(_17050_),
    .A2(_17052_),
    .ZN(_17053_)
  );
  INV_X1 _52547_ (
    .A(_17053_),
    .ZN(_01321_)
  );
  AND2_X1 _52548_ (
    .A1(_12696_),
    .A2(_13169_),
    .ZN(_17054_)
  );
  INV_X1 _52549_ (
    .A(_17054_),
    .ZN(_17055_)
  );
  AND2_X1 _52550_ (
    .A1(\cpuregs[30] [20]),
    .A2(_12697_),
    .ZN(_17056_)
  );
  INV_X1 _52551_ (
    .A(_17056_),
    .ZN(_17057_)
  );
  AND2_X1 _52552_ (
    .A1(_17055_),
    .A2(_17057_),
    .ZN(_17058_)
  );
  INV_X1 _52553_ (
    .A(_17058_),
    .ZN(_01322_)
  );
  AND2_X1 _52554_ (
    .A1(_12696_),
    .A2(_13184_),
    .ZN(_17059_)
  );
  INV_X1 _52555_ (
    .A(_17059_),
    .ZN(_17060_)
  );
  AND2_X1 _52556_ (
    .A1(\cpuregs[30] [21]),
    .A2(_12697_),
    .ZN(_17061_)
  );
  INV_X1 _52557_ (
    .A(_17061_),
    .ZN(_17062_)
  );
  AND2_X1 _52558_ (
    .A1(_17060_),
    .A2(_17062_),
    .ZN(_17063_)
  );
  INV_X1 _52559_ (
    .A(_17063_),
    .ZN(_01323_)
  );
  AND2_X1 _52560_ (
    .A1(_12696_),
    .A2(_13199_),
    .ZN(_17064_)
  );
  INV_X1 _52561_ (
    .A(_17064_),
    .ZN(_17065_)
  );
  AND2_X1 _52562_ (
    .A1(\cpuregs[30] [22]),
    .A2(_12697_),
    .ZN(_17066_)
  );
  INV_X1 _52563_ (
    .A(_17066_),
    .ZN(_17067_)
  );
  AND2_X1 _52564_ (
    .A1(_17065_),
    .A2(_17067_),
    .ZN(_17068_)
  );
  INV_X1 _52565_ (
    .A(_17068_),
    .ZN(_01324_)
  );
  AND2_X1 _52566_ (
    .A1(_12696_),
    .A2(_13214_),
    .ZN(_17069_)
  );
  INV_X1 _52567_ (
    .A(_17069_),
    .ZN(_17070_)
  );
  AND2_X1 _52568_ (
    .A1(\cpuregs[30] [23]),
    .A2(_12697_),
    .ZN(_17071_)
  );
  INV_X1 _52569_ (
    .A(_17071_),
    .ZN(_17072_)
  );
  AND2_X1 _52570_ (
    .A1(_17070_),
    .A2(_17072_),
    .ZN(_17073_)
  );
  INV_X1 _52571_ (
    .A(_17073_),
    .ZN(_01325_)
  );
  AND2_X1 _52572_ (
    .A1(_12696_),
    .A2(_13229_),
    .ZN(_17074_)
  );
  INV_X1 _52573_ (
    .A(_17074_),
    .ZN(_17075_)
  );
  AND2_X1 _52574_ (
    .A1(\cpuregs[30] [24]),
    .A2(_12697_),
    .ZN(_17076_)
  );
  INV_X1 _52575_ (
    .A(_17076_),
    .ZN(_17077_)
  );
  AND2_X1 _52576_ (
    .A1(_17075_),
    .A2(_17077_),
    .ZN(_17078_)
  );
  INV_X1 _52577_ (
    .A(_17078_),
    .ZN(_01326_)
  );
  AND2_X1 _52578_ (
    .A1(_12696_),
    .A2(_13244_),
    .ZN(_17079_)
  );
  INV_X1 _52579_ (
    .A(_17079_),
    .ZN(_17080_)
  );
  AND2_X1 _52580_ (
    .A1(\cpuregs[30] [25]),
    .A2(_12697_),
    .ZN(_17081_)
  );
  INV_X1 _52581_ (
    .A(_17081_),
    .ZN(_17082_)
  );
  AND2_X1 _52582_ (
    .A1(_17080_),
    .A2(_17082_),
    .ZN(_17083_)
  );
  INV_X1 _52583_ (
    .A(_17083_),
    .ZN(_01327_)
  );
  AND2_X1 _52584_ (
    .A1(_12696_),
    .A2(_13259_),
    .ZN(_17084_)
  );
  INV_X1 _52585_ (
    .A(_17084_),
    .ZN(_17085_)
  );
  AND2_X1 _52586_ (
    .A1(\cpuregs[30] [26]),
    .A2(_12697_),
    .ZN(_17086_)
  );
  INV_X1 _52587_ (
    .A(_17086_),
    .ZN(_17087_)
  );
  AND2_X1 _52588_ (
    .A1(_17085_),
    .A2(_17087_),
    .ZN(_17088_)
  );
  INV_X1 _52589_ (
    .A(_17088_),
    .ZN(_01328_)
  );
  AND2_X1 _52590_ (
    .A1(_12696_),
    .A2(_13274_),
    .ZN(_17089_)
  );
  INV_X1 _52591_ (
    .A(_17089_),
    .ZN(_17090_)
  );
  AND2_X1 _52592_ (
    .A1(\cpuregs[30] [27]),
    .A2(_12697_),
    .ZN(_17091_)
  );
  INV_X1 _52593_ (
    .A(_17091_),
    .ZN(_17092_)
  );
  AND2_X1 _52594_ (
    .A1(_17090_),
    .A2(_17092_),
    .ZN(_17093_)
  );
  INV_X1 _52595_ (
    .A(_17093_),
    .ZN(_01329_)
  );
  AND2_X1 _52596_ (
    .A1(_12696_),
    .A2(_13289_),
    .ZN(_17094_)
  );
  INV_X1 _52597_ (
    .A(_17094_),
    .ZN(_17095_)
  );
  AND2_X1 _52598_ (
    .A1(\cpuregs[30] [28]),
    .A2(_12697_),
    .ZN(_17096_)
  );
  INV_X1 _52599_ (
    .A(_17096_),
    .ZN(_17097_)
  );
  AND2_X1 _52600_ (
    .A1(_17095_),
    .A2(_17097_),
    .ZN(_17098_)
  );
  INV_X1 _52601_ (
    .A(_17098_),
    .ZN(_01330_)
  );
  AND2_X1 _52602_ (
    .A1(_12696_),
    .A2(_13304_),
    .ZN(_17099_)
  );
  INV_X1 _52603_ (
    .A(_17099_),
    .ZN(_17100_)
  );
  AND2_X1 _52604_ (
    .A1(\cpuregs[30] [29]),
    .A2(_12697_),
    .ZN(_17101_)
  );
  INV_X1 _52605_ (
    .A(_17101_),
    .ZN(_17102_)
  );
  AND2_X1 _52606_ (
    .A1(_17100_),
    .A2(_17102_),
    .ZN(_17103_)
  );
  INV_X1 _52607_ (
    .A(_17103_),
    .ZN(_01331_)
  );
  AND2_X1 _52608_ (
    .A1(_12696_),
    .A2(_13319_),
    .ZN(_17104_)
  );
  INV_X1 _52609_ (
    .A(_17104_),
    .ZN(_17105_)
  );
  AND2_X1 _52610_ (
    .A1(\cpuregs[30] [30]),
    .A2(_12697_),
    .ZN(_17106_)
  );
  INV_X1 _52611_ (
    .A(_17106_),
    .ZN(_17107_)
  );
  AND2_X1 _52612_ (
    .A1(_17105_),
    .A2(_17107_),
    .ZN(_17108_)
  );
  INV_X1 _52613_ (
    .A(_17108_),
    .ZN(_01332_)
  );
  AND2_X1 _52614_ (
    .A1(_12732_),
    .A2(_12872_),
    .ZN(_17109_)
  );
  INV_X1 _52615_ (
    .A(_17109_),
    .ZN(_17110_)
  );
  AND2_X1 _52616_ (
    .A1(_21865_),
    .A2(_12733_),
    .ZN(_17111_)
  );
  INV_X1 _52617_ (
    .A(_17111_),
    .ZN(_17112_)
  );
  AND2_X1 _52618_ (
    .A1(_17110_),
    .A2(_17112_),
    .ZN(_01333_)
  );
  AND2_X1 _52619_ (
    .A1(_12732_),
    .A2(_12884_),
    .ZN(_17113_)
  );
  INV_X1 _52620_ (
    .A(_17113_),
    .ZN(_17114_)
  );
  AND2_X1 _52621_ (
    .A1(_21866_),
    .A2(_12733_),
    .ZN(_17115_)
  );
  INV_X1 _52622_ (
    .A(_17115_),
    .ZN(_17116_)
  );
  AND2_X1 _52623_ (
    .A1(_17114_),
    .A2(_17116_),
    .ZN(_01334_)
  );
  AND2_X1 _52624_ (
    .A1(_12732_),
    .A2(_12898_),
    .ZN(_17117_)
  );
  INV_X1 _52625_ (
    .A(_17117_),
    .ZN(_17118_)
  );
  AND2_X1 _52626_ (
    .A1(_21867_),
    .A2(_12733_),
    .ZN(_17119_)
  );
  INV_X1 _52627_ (
    .A(_17119_),
    .ZN(_17120_)
  );
  AND2_X1 _52628_ (
    .A1(_17118_),
    .A2(_17120_),
    .ZN(_01335_)
  );
  AND2_X1 _52629_ (
    .A1(_12732_),
    .A2(_12913_),
    .ZN(_17121_)
  );
  INV_X1 _52630_ (
    .A(_17121_),
    .ZN(_17122_)
  );
  AND2_X1 _52631_ (
    .A1(\cpuregs[26] [3]),
    .A2(_12733_),
    .ZN(_17123_)
  );
  INV_X1 _52632_ (
    .A(_17123_),
    .ZN(_17124_)
  );
  AND2_X1 _52633_ (
    .A1(_17122_),
    .A2(_17124_),
    .ZN(_17125_)
  );
  INV_X1 _52634_ (
    .A(_17125_),
    .ZN(_01336_)
  );
  AND2_X1 _52635_ (
    .A1(_12732_),
    .A2(_12928_),
    .ZN(_17126_)
  );
  INV_X1 _52636_ (
    .A(_17126_),
    .ZN(_17127_)
  );
  AND2_X1 _52637_ (
    .A1(\cpuregs[26] [4]),
    .A2(_12733_),
    .ZN(_17128_)
  );
  INV_X1 _52638_ (
    .A(_17128_),
    .ZN(_17129_)
  );
  AND2_X1 _52639_ (
    .A1(_17127_),
    .A2(_17129_),
    .ZN(_17130_)
  );
  INV_X1 _52640_ (
    .A(_17130_),
    .ZN(_01337_)
  );
  AND2_X1 _52641_ (
    .A1(_12732_),
    .A2(_12941_),
    .ZN(_17131_)
  );
  INV_X1 _52642_ (
    .A(_17131_),
    .ZN(_17132_)
  );
  AND2_X1 _52643_ (
    .A1(_21868_),
    .A2(_12733_),
    .ZN(_17133_)
  );
  INV_X1 _52644_ (
    .A(_17133_),
    .ZN(_17134_)
  );
  AND2_X1 _52645_ (
    .A1(_17132_),
    .A2(_17134_),
    .ZN(_01338_)
  );
  AND2_X1 _52646_ (
    .A1(_12732_),
    .A2(_12956_),
    .ZN(_17135_)
  );
  INV_X1 _52647_ (
    .A(_17135_),
    .ZN(_17136_)
  );
  AND2_X1 _52648_ (
    .A1(_21869_),
    .A2(_12733_),
    .ZN(_17137_)
  );
  INV_X1 _52649_ (
    .A(_17137_),
    .ZN(_17138_)
  );
  AND2_X1 _52650_ (
    .A1(_17136_),
    .A2(_17138_),
    .ZN(_01339_)
  );
  AND2_X1 _52651_ (
    .A1(_12732_),
    .A2(_12971_),
    .ZN(_17139_)
  );
  INV_X1 _52652_ (
    .A(_17139_),
    .ZN(_17140_)
  );
  AND2_X1 _52653_ (
    .A1(_21870_),
    .A2(_12733_),
    .ZN(_17141_)
  );
  INV_X1 _52654_ (
    .A(_17141_),
    .ZN(_17142_)
  );
  AND2_X1 _52655_ (
    .A1(_17140_),
    .A2(_17142_),
    .ZN(_01340_)
  );
  AND2_X1 _52656_ (
    .A1(_12732_),
    .A2(_12986_),
    .ZN(_17143_)
  );
  INV_X1 _52657_ (
    .A(_17143_),
    .ZN(_17144_)
  );
  AND2_X1 _52658_ (
    .A1(_21871_),
    .A2(_12733_),
    .ZN(_17145_)
  );
  INV_X1 _52659_ (
    .A(_17145_),
    .ZN(_17146_)
  );
  AND2_X1 _52660_ (
    .A1(_17144_),
    .A2(_17146_),
    .ZN(_01341_)
  );
  AND2_X1 _52661_ (
    .A1(_12732_),
    .A2(_13001_),
    .ZN(_17147_)
  );
  INV_X1 _52662_ (
    .A(_17147_),
    .ZN(_17148_)
  );
  AND2_X1 _52663_ (
    .A1(_21872_),
    .A2(_12733_),
    .ZN(_17149_)
  );
  INV_X1 _52664_ (
    .A(_17149_),
    .ZN(_17150_)
  );
  AND2_X1 _52665_ (
    .A1(_17148_),
    .A2(_17150_),
    .ZN(_01342_)
  );
  AND2_X1 _52666_ (
    .A1(_12732_),
    .A2(_13016_),
    .ZN(_17151_)
  );
  INV_X1 _52667_ (
    .A(_17151_),
    .ZN(_17152_)
  );
  AND2_X1 _52668_ (
    .A1(_21873_),
    .A2(_12733_),
    .ZN(_17153_)
  );
  INV_X1 _52669_ (
    .A(_17153_),
    .ZN(_17154_)
  );
  AND2_X1 _52670_ (
    .A1(_17152_),
    .A2(_17154_),
    .ZN(_01343_)
  );
  AND2_X1 _52671_ (
    .A1(_12732_),
    .A2(_13031_),
    .ZN(_17155_)
  );
  INV_X1 _52672_ (
    .A(_17155_),
    .ZN(_17156_)
  );
  AND2_X1 _52673_ (
    .A1(_21874_),
    .A2(_12733_),
    .ZN(_17157_)
  );
  INV_X1 _52674_ (
    .A(_17157_),
    .ZN(_17158_)
  );
  AND2_X1 _52675_ (
    .A1(_17156_),
    .A2(_17158_),
    .ZN(_01344_)
  );
  AND2_X1 _52676_ (
    .A1(_12732_),
    .A2(_13046_),
    .ZN(_17159_)
  );
  INV_X1 _52677_ (
    .A(_17159_),
    .ZN(_17160_)
  );
  AND2_X1 _52678_ (
    .A1(_21875_),
    .A2(_12733_),
    .ZN(_17161_)
  );
  INV_X1 _52679_ (
    .A(_17161_),
    .ZN(_17162_)
  );
  AND2_X1 _52680_ (
    .A1(_17160_),
    .A2(_17162_),
    .ZN(_01345_)
  );
  AND2_X1 _52681_ (
    .A1(_12732_),
    .A2(_13061_),
    .ZN(_17163_)
  );
  INV_X1 _52682_ (
    .A(_17163_),
    .ZN(_17164_)
  );
  AND2_X1 _52683_ (
    .A1(_21876_),
    .A2(_12733_),
    .ZN(_17165_)
  );
  INV_X1 _52684_ (
    .A(_17165_),
    .ZN(_17166_)
  );
  AND2_X1 _52685_ (
    .A1(_17164_),
    .A2(_17166_),
    .ZN(_01346_)
  );
  AND2_X1 _52686_ (
    .A1(_12732_),
    .A2(_13078_),
    .ZN(_17167_)
  );
  INV_X1 _52687_ (
    .A(_17167_),
    .ZN(_17168_)
  );
  AND2_X1 _52688_ (
    .A1(\cpuregs[26] [14]),
    .A2(_12733_),
    .ZN(_17169_)
  );
  INV_X1 _52689_ (
    .A(_17169_),
    .ZN(_17170_)
  );
  AND2_X1 _52690_ (
    .A1(_17168_),
    .A2(_17170_),
    .ZN(_17171_)
  );
  INV_X1 _52691_ (
    .A(_17171_),
    .ZN(_01347_)
  );
  AND2_X1 _52692_ (
    .A1(_12732_),
    .A2(_13091_),
    .ZN(_17172_)
  );
  INV_X1 _52693_ (
    .A(_17172_),
    .ZN(_17173_)
  );
  AND2_X1 _52694_ (
    .A1(_21877_),
    .A2(_12733_),
    .ZN(_17174_)
  );
  INV_X1 _52695_ (
    .A(_17174_),
    .ZN(_17175_)
  );
  AND2_X1 _52696_ (
    .A1(_17173_),
    .A2(_17175_),
    .ZN(_01348_)
  );
  AND2_X1 _52697_ (
    .A1(\cpuregs[26] [16]),
    .A2(_12733_),
    .ZN(_17176_)
  );
  INV_X1 _52698_ (
    .A(_17176_),
    .ZN(_17177_)
  );
  AND2_X1 _52699_ (
    .A1(_12732_),
    .A2(_13108_),
    .ZN(_17178_)
  );
  INV_X1 _52700_ (
    .A(_17178_),
    .ZN(_17179_)
  );
  AND2_X1 _52701_ (
    .A1(_17177_),
    .A2(_17179_),
    .ZN(_17180_)
  );
  INV_X1 _52702_ (
    .A(_17180_),
    .ZN(_01349_)
  );
  AND2_X1 _52703_ (
    .A1(_12732_),
    .A2(_13121_),
    .ZN(_17181_)
  );
  INV_X1 _52704_ (
    .A(_17181_),
    .ZN(_17182_)
  );
  AND2_X1 _52705_ (
    .A1(_21879_),
    .A2(_12733_),
    .ZN(_17183_)
  );
  INV_X1 _52706_ (
    .A(_17183_),
    .ZN(_17184_)
  );
  AND2_X1 _52707_ (
    .A1(_17182_),
    .A2(_17184_),
    .ZN(_01350_)
  );
  AND2_X1 _52708_ (
    .A1(_12732_),
    .A2(_13139_),
    .ZN(_17185_)
  );
  INV_X1 _52709_ (
    .A(_17185_),
    .ZN(_17186_)
  );
  AND2_X1 _52710_ (
    .A1(\cpuregs[26] [18]),
    .A2(_12733_),
    .ZN(_17187_)
  );
  INV_X1 _52711_ (
    .A(_17187_),
    .ZN(_17188_)
  );
  AND2_X1 _52712_ (
    .A1(_17186_),
    .A2(_17188_),
    .ZN(_17189_)
  );
  INV_X1 _52713_ (
    .A(_17189_),
    .ZN(_01351_)
  );
  AND2_X1 _52714_ (
    .A1(_12732_),
    .A2(_13152_),
    .ZN(_17190_)
  );
  INV_X1 _52715_ (
    .A(_17190_),
    .ZN(_17191_)
  );
  AND2_X1 _52716_ (
    .A1(_21880_),
    .A2(_12733_),
    .ZN(_17192_)
  );
  INV_X1 _52717_ (
    .A(_17192_),
    .ZN(_17193_)
  );
  AND2_X1 _52718_ (
    .A1(_17191_),
    .A2(_17193_),
    .ZN(_01352_)
  );
  AND2_X1 _52719_ (
    .A1(_12732_),
    .A2(_13169_),
    .ZN(_17194_)
  );
  INV_X1 _52720_ (
    .A(_17194_),
    .ZN(_17195_)
  );
  AND2_X1 _52721_ (
    .A1(\cpuregs[26] [20]),
    .A2(_12733_),
    .ZN(_17196_)
  );
  INV_X1 _52722_ (
    .A(_17196_),
    .ZN(_17197_)
  );
  AND2_X1 _52723_ (
    .A1(_17195_),
    .A2(_17197_),
    .ZN(_17198_)
  );
  INV_X1 _52724_ (
    .A(_17198_),
    .ZN(_01353_)
  );
  AND2_X1 _52725_ (
    .A1(_12732_),
    .A2(_13182_),
    .ZN(_17199_)
  );
  INV_X1 _52726_ (
    .A(_17199_),
    .ZN(_17200_)
  );
  AND2_X1 _52727_ (
    .A1(_21881_),
    .A2(_12733_),
    .ZN(_17201_)
  );
  INV_X1 _52728_ (
    .A(_17201_),
    .ZN(_17202_)
  );
  AND2_X1 _52729_ (
    .A1(_17200_),
    .A2(_17202_),
    .ZN(_01354_)
  );
  AND2_X1 _52730_ (
    .A1(_12732_),
    .A2(_13199_),
    .ZN(_17203_)
  );
  INV_X1 _52731_ (
    .A(_17203_),
    .ZN(_17204_)
  );
  AND2_X1 _52732_ (
    .A1(\cpuregs[26] [22]),
    .A2(_12733_),
    .ZN(_17205_)
  );
  INV_X1 _52733_ (
    .A(_17205_),
    .ZN(_17206_)
  );
  AND2_X1 _52734_ (
    .A1(_17204_),
    .A2(_17206_),
    .ZN(_17207_)
  );
  INV_X1 _52735_ (
    .A(_17207_),
    .ZN(_01355_)
  );
  AND2_X1 _52736_ (
    .A1(_12732_),
    .A2(_13212_),
    .ZN(_17208_)
  );
  INV_X1 _52737_ (
    .A(_17208_),
    .ZN(_17209_)
  );
  AND2_X1 _52738_ (
    .A1(_21882_),
    .A2(_12733_),
    .ZN(_17210_)
  );
  INV_X1 _52739_ (
    .A(_17210_),
    .ZN(_17211_)
  );
  AND2_X1 _52740_ (
    .A1(_17209_),
    .A2(_17211_),
    .ZN(_01356_)
  );
  AND2_X1 _52741_ (
    .A1(_12732_),
    .A2(_13229_),
    .ZN(_17212_)
  );
  INV_X1 _52742_ (
    .A(_17212_),
    .ZN(_17213_)
  );
  AND2_X1 _52743_ (
    .A1(\cpuregs[26] [24]),
    .A2(_12733_),
    .ZN(_17214_)
  );
  INV_X1 _52744_ (
    .A(_17214_),
    .ZN(_17215_)
  );
  AND2_X1 _52745_ (
    .A1(_17213_),
    .A2(_17215_),
    .ZN(_17216_)
  );
  INV_X1 _52746_ (
    .A(_17216_),
    .ZN(_01357_)
  );
  AND2_X1 _52747_ (
    .A1(_12732_),
    .A2(_13242_),
    .ZN(_17217_)
  );
  INV_X1 _52748_ (
    .A(_17217_),
    .ZN(_17218_)
  );
  AND2_X1 _52749_ (
    .A1(_21883_),
    .A2(_12733_),
    .ZN(_17219_)
  );
  INV_X1 _52750_ (
    .A(_17219_),
    .ZN(_17220_)
  );
  AND2_X1 _52751_ (
    .A1(_17218_),
    .A2(_17220_),
    .ZN(_01358_)
  );
  AND2_X1 _52752_ (
    .A1(_12732_),
    .A2(_13257_),
    .ZN(_17221_)
  );
  INV_X1 _52753_ (
    .A(_17221_),
    .ZN(_17222_)
  );
  AND2_X1 _52754_ (
    .A1(_21884_),
    .A2(_12733_),
    .ZN(_17223_)
  );
  INV_X1 _52755_ (
    .A(_17223_),
    .ZN(_17224_)
  );
  AND2_X1 _52756_ (
    .A1(_17222_),
    .A2(_17224_),
    .ZN(_01359_)
  );
  AND2_X1 _52757_ (
    .A1(_12732_),
    .A2(_13272_),
    .ZN(_17225_)
  );
  INV_X1 _52758_ (
    .A(_17225_),
    .ZN(_17226_)
  );
  AND2_X1 _52759_ (
    .A1(_21885_),
    .A2(_12733_),
    .ZN(_17227_)
  );
  INV_X1 _52760_ (
    .A(_17227_),
    .ZN(_17228_)
  );
  AND2_X1 _52761_ (
    .A1(_17226_),
    .A2(_17228_),
    .ZN(_01360_)
  );
  AND2_X1 _52762_ (
    .A1(_12732_),
    .A2(_13289_),
    .ZN(_17229_)
  );
  INV_X1 _52763_ (
    .A(_17229_),
    .ZN(_17230_)
  );
  AND2_X1 _52764_ (
    .A1(\cpuregs[26] [28]),
    .A2(_12733_),
    .ZN(_17231_)
  );
  INV_X1 _52765_ (
    .A(_17231_),
    .ZN(_17232_)
  );
  AND2_X1 _52766_ (
    .A1(_17230_),
    .A2(_17232_),
    .ZN(_17233_)
  );
  INV_X1 _52767_ (
    .A(_17233_),
    .ZN(_01361_)
  );
  AND2_X1 _52768_ (
    .A1(_12732_),
    .A2(_13302_),
    .ZN(_17234_)
  );
  INV_X1 _52769_ (
    .A(_17234_),
    .ZN(_17235_)
  );
  AND2_X1 _52770_ (
    .A1(_21887_),
    .A2(_12733_),
    .ZN(_17236_)
  );
  INV_X1 _52771_ (
    .A(_17236_),
    .ZN(_17237_)
  );
  AND2_X1 _52772_ (
    .A1(_17235_),
    .A2(_17237_),
    .ZN(_01362_)
  );
  AND2_X1 _52773_ (
    .A1(_12732_),
    .A2(_13317_),
    .ZN(_17238_)
  );
  INV_X1 _52774_ (
    .A(_17238_),
    .ZN(_17239_)
  );
  AND2_X1 _52775_ (
    .A1(_21888_),
    .A2(_12733_),
    .ZN(_17240_)
  );
  INV_X1 _52776_ (
    .A(_17240_),
    .ZN(_17241_)
  );
  AND2_X1 _52777_ (
    .A1(_17239_),
    .A2(_17241_),
    .ZN(_01363_)
  );
  AND2_X1 _52778_ (
    .A1(_12710_),
    .A2(_12874_),
    .ZN(_17242_)
  );
  INV_X1 _52779_ (
    .A(_17242_),
    .ZN(_17243_)
  );
  AND2_X1 _52780_ (
    .A1(\cpuregs[29] [0]),
    .A2(_12711_),
    .ZN(_17244_)
  );
  INV_X1 _52781_ (
    .A(_17244_),
    .ZN(_17245_)
  );
  AND2_X1 _52782_ (
    .A1(_17243_),
    .A2(_17245_),
    .ZN(_17246_)
  );
  INV_X1 _52783_ (
    .A(_17246_),
    .ZN(_01364_)
  );
  AND2_X1 _52784_ (
    .A1(_12710_),
    .A2(_12886_),
    .ZN(_17247_)
  );
  INV_X1 _52785_ (
    .A(_17247_),
    .ZN(_17248_)
  );
  AND2_X1 _52786_ (
    .A1(\cpuregs[29] [1]),
    .A2(_12711_),
    .ZN(_17249_)
  );
  INV_X1 _52787_ (
    .A(_17249_),
    .ZN(_17250_)
  );
  AND2_X1 _52788_ (
    .A1(_17248_),
    .A2(_17250_),
    .ZN(_17251_)
  );
  INV_X1 _52789_ (
    .A(_17251_),
    .ZN(_01365_)
  );
  AND2_X1 _52790_ (
    .A1(\cpuregs[29] [2]),
    .A2(_12711_),
    .ZN(_17252_)
  );
  INV_X1 _52791_ (
    .A(_17252_),
    .ZN(_17253_)
  );
  AND2_X1 _52792_ (
    .A1(_12710_),
    .A2(_12900_),
    .ZN(_17254_)
  );
  INV_X1 _52793_ (
    .A(_17254_),
    .ZN(_17255_)
  );
  AND2_X1 _52794_ (
    .A1(_17253_),
    .A2(_17255_),
    .ZN(_17256_)
  );
  INV_X1 _52795_ (
    .A(_17256_),
    .ZN(_01366_)
  );
  AND2_X1 _52796_ (
    .A1(_12710_),
    .A2(_12913_),
    .ZN(_17257_)
  );
  INV_X1 _52797_ (
    .A(_17257_),
    .ZN(_17258_)
  );
  AND2_X1 _52798_ (
    .A1(\cpuregs[29] [3]),
    .A2(_12711_),
    .ZN(_17259_)
  );
  INV_X1 _52799_ (
    .A(_17259_),
    .ZN(_17260_)
  );
  AND2_X1 _52800_ (
    .A1(_17258_),
    .A2(_17260_),
    .ZN(_17261_)
  );
  INV_X1 _52801_ (
    .A(_17261_),
    .ZN(_01367_)
  );
  AND2_X1 _52802_ (
    .A1(_12710_),
    .A2(_12928_),
    .ZN(_17262_)
  );
  INV_X1 _52803_ (
    .A(_17262_),
    .ZN(_17263_)
  );
  AND2_X1 _52804_ (
    .A1(\cpuregs[29] [4]),
    .A2(_12711_),
    .ZN(_17264_)
  );
  INV_X1 _52805_ (
    .A(_17264_),
    .ZN(_17265_)
  );
  AND2_X1 _52806_ (
    .A1(_17263_),
    .A2(_17265_),
    .ZN(_17266_)
  );
  INV_X1 _52807_ (
    .A(_17266_),
    .ZN(_01368_)
  );
  AND2_X1 _52808_ (
    .A1(_12710_),
    .A2(_12943_),
    .ZN(_17267_)
  );
  INV_X1 _52809_ (
    .A(_17267_),
    .ZN(_17268_)
  );
  AND2_X1 _52810_ (
    .A1(\cpuregs[29] [5]),
    .A2(_12711_),
    .ZN(_17269_)
  );
  INV_X1 _52811_ (
    .A(_17269_),
    .ZN(_17270_)
  );
  AND2_X1 _52812_ (
    .A1(_17268_),
    .A2(_17270_),
    .ZN(_17271_)
  );
  INV_X1 _52813_ (
    .A(_17271_),
    .ZN(_01369_)
  );
  AND2_X1 _52814_ (
    .A1(_12710_),
    .A2(_12958_),
    .ZN(_17272_)
  );
  INV_X1 _52815_ (
    .A(_17272_),
    .ZN(_17273_)
  );
  AND2_X1 _52816_ (
    .A1(\cpuregs[29] [6]),
    .A2(_12711_),
    .ZN(_17274_)
  );
  INV_X1 _52817_ (
    .A(_17274_),
    .ZN(_17275_)
  );
  AND2_X1 _52818_ (
    .A1(_17273_),
    .A2(_17275_),
    .ZN(_17276_)
  );
  INV_X1 _52819_ (
    .A(_17276_),
    .ZN(_01370_)
  );
  AND2_X1 _52820_ (
    .A1(_12710_),
    .A2(_12973_),
    .ZN(_17277_)
  );
  INV_X1 _52821_ (
    .A(_17277_),
    .ZN(_17278_)
  );
  AND2_X1 _52822_ (
    .A1(\cpuregs[29] [7]),
    .A2(_12711_),
    .ZN(_17279_)
  );
  INV_X1 _52823_ (
    .A(_17279_),
    .ZN(_17280_)
  );
  AND2_X1 _52824_ (
    .A1(_17278_),
    .A2(_17280_),
    .ZN(_17281_)
  );
  INV_X1 _52825_ (
    .A(_17281_),
    .ZN(_01371_)
  );
  AND2_X1 _52826_ (
    .A1(_12710_),
    .A2(_12988_),
    .ZN(_17282_)
  );
  INV_X1 _52827_ (
    .A(_17282_),
    .ZN(_17283_)
  );
  AND2_X1 _52828_ (
    .A1(\cpuregs[29] [8]),
    .A2(_12711_),
    .ZN(_17284_)
  );
  INV_X1 _52829_ (
    .A(_17284_),
    .ZN(_17285_)
  );
  AND2_X1 _52830_ (
    .A1(_17283_),
    .A2(_17285_),
    .ZN(_17286_)
  );
  INV_X1 _52831_ (
    .A(_17286_),
    .ZN(_01372_)
  );
  AND2_X1 _52832_ (
    .A1(_12710_),
    .A2(_13003_),
    .ZN(_17287_)
  );
  INV_X1 _52833_ (
    .A(_17287_),
    .ZN(_17288_)
  );
  AND2_X1 _52834_ (
    .A1(\cpuregs[29] [9]),
    .A2(_12711_),
    .ZN(_17289_)
  );
  INV_X1 _52835_ (
    .A(_17289_),
    .ZN(_17290_)
  );
  AND2_X1 _52836_ (
    .A1(_17288_),
    .A2(_17290_),
    .ZN(_17291_)
  );
  INV_X1 _52837_ (
    .A(_17291_),
    .ZN(_01373_)
  );
  AND2_X1 _52838_ (
    .A1(_12710_),
    .A2(_13018_),
    .ZN(_17292_)
  );
  INV_X1 _52839_ (
    .A(_17292_),
    .ZN(_17293_)
  );
  AND2_X1 _52840_ (
    .A1(\cpuregs[29] [10]),
    .A2(_12711_),
    .ZN(_17294_)
  );
  INV_X1 _52841_ (
    .A(_17294_),
    .ZN(_17295_)
  );
  AND2_X1 _52842_ (
    .A1(_17293_),
    .A2(_17295_),
    .ZN(_17296_)
  );
  INV_X1 _52843_ (
    .A(_17296_),
    .ZN(_01374_)
  );
  AND2_X1 _52844_ (
    .A1(_12710_),
    .A2(_13033_),
    .ZN(_17297_)
  );
  INV_X1 _52845_ (
    .A(_17297_),
    .ZN(_17298_)
  );
  AND2_X1 _52846_ (
    .A1(\cpuregs[29] [11]),
    .A2(_12711_),
    .ZN(_17299_)
  );
  INV_X1 _52847_ (
    .A(_17299_),
    .ZN(_17300_)
  );
  AND2_X1 _52848_ (
    .A1(_17298_),
    .A2(_17300_),
    .ZN(_17301_)
  );
  INV_X1 _52849_ (
    .A(_17301_),
    .ZN(_01375_)
  );
  AND2_X1 _52850_ (
    .A1(_12710_),
    .A2(_13048_),
    .ZN(_17302_)
  );
  INV_X1 _52851_ (
    .A(_17302_),
    .ZN(_17303_)
  );
  AND2_X1 _52852_ (
    .A1(\cpuregs[29] [12]),
    .A2(_12711_),
    .ZN(_17304_)
  );
  INV_X1 _52853_ (
    .A(_17304_),
    .ZN(_17305_)
  );
  AND2_X1 _52854_ (
    .A1(_17303_),
    .A2(_17305_),
    .ZN(_17306_)
  );
  INV_X1 _52855_ (
    .A(_17306_),
    .ZN(_01376_)
  );
  AND2_X1 _52856_ (
    .A1(_12710_),
    .A2(_13063_),
    .ZN(_17307_)
  );
  INV_X1 _52857_ (
    .A(_17307_),
    .ZN(_17308_)
  );
  AND2_X1 _52858_ (
    .A1(\cpuregs[29] [13]),
    .A2(_12711_),
    .ZN(_17309_)
  );
  INV_X1 _52859_ (
    .A(_17309_),
    .ZN(_17310_)
  );
  AND2_X1 _52860_ (
    .A1(_17308_),
    .A2(_17310_),
    .ZN(_17311_)
  );
  INV_X1 _52861_ (
    .A(_17311_),
    .ZN(_01377_)
  );
  AND2_X1 _52862_ (
    .A1(_12710_),
    .A2(_13078_),
    .ZN(_17312_)
  );
  INV_X1 _52863_ (
    .A(_17312_),
    .ZN(_17313_)
  );
  AND2_X1 _52864_ (
    .A1(\cpuregs[29] [14]),
    .A2(_12711_),
    .ZN(_17314_)
  );
  INV_X1 _52865_ (
    .A(_17314_),
    .ZN(_17315_)
  );
  AND2_X1 _52866_ (
    .A1(_17313_),
    .A2(_17315_),
    .ZN(_17316_)
  );
  INV_X1 _52867_ (
    .A(_17316_),
    .ZN(_01378_)
  );
  AND2_X1 _52868_ (
    .A1(_12710_),
    .A2(_13093_),
    .ZN(_17317_)
  );
  INV_X1 _52869_ (
    .A(_17317_),
    .ZN(_17318_)
  );
  AND2_X1 _52870_ (
    .A1(\cpuregs[29] [15]),
    .A2(_12711_),
    .ZN(_17319_)
  );
  INV_X1 _52871_ (
    .A(_17319_),
    .ZN(_17320_)
  );
  AND2_X1 _52872_ (
    .A1(_17318_),
    .A2(_17320_),
    .ZN(_17321_)
  );
  INV_X1 _52873_ (
    .A(_17321_),
    .ZN(_01379_)
  );
  AND2_X1 _52874_ (
    .A1(_12710_),
    .A2(_13108_),
    .ZN(_17322_)
  );
  INV_X1 _52875_ (
    .A(_17322_),
    .ZN(_17323_)
  );
  AND2_X1 _52876_ (
    .A1(\cpuregs[29] [16]),
    .A2(_12711_),
    .ZN(_17324_)
  );
  INV_X1 _52877_ (
    .A(_17324_),
    .ZN(_17325_)
  );
  AND2_X1 _52878_ (
    .A1(_17323_),
    .A2(_17325_),
    .ZN(_17326_)
  );
  INV_X1 _52879_ (
    .A(_17326_),
    .ZN(_01380_)
  );
  AND2_X1 _52880_ (
    .A1(_12710_),
    .A2(_13123_),
    .ZN(_17327_)
  );
  INV_X1 _52881_ (
    .A(_17327_),
    .ZN(_17328_)
  );
  AND2_X1 _52882_ (
    .A1(\cpuregs[29] [17]),
    .A2(_12711_),
    .ZN(_17329_)
  );
  INV_X1 _52883_ (
    .A(_17329_),
    .ZN(_17330_)
  );
  AND2_X1 _52884_ (
    .A1(_17328_),
    .A2(_17330_),
    .ZN(_17331_)
  );
  INV_X1 _52885_ (
    .A(_17331_),
    .ZN(_01381_)
  );
  AND2_X1 _52886_ (
    .A1(_12710_),
    .A2(_13139_),
    .ZN(_17332_)
  );
  INV_X1 _52887_ (
    .A(_17332_),
    .ZN(_17333_)
  );
  AND2_X1 _52888_ (
    .A1(\cpuregs[29] [18]),
    .A2(_12711_),
    .ZN(_17334_)
  );
  INV_X1 _52889_ (
    .A(_17334_),
    .ZN(_17335_)
  );
  AND2_X1 _52890_ (
    .A1(_17333_),
    .A2(_17335_),
    .ZN(_17336_)
  );
  INV_X1 _52891_ (
    .A(_17336_),
    .ZN(_01382_)
  );
  AND2_X1 _52892_ (
    .A1(_12710_),
    .A2(_13154_),
    .ZN(_17337_)
  );
  INV_X1 _52893_ (
    .A(_17337_),
    .ZN(_17338_)
  );
  AND2_X1 _52894_ (
    .A1(\cpuregs[29] [19]),
    .A2(_12711_),
    .ZN(_17339_)
  );
  INV_X1 _52895_ (
    .A(_17339_),
    .ZN(_17340_)
  );
  AND2_X1 _52896_ (
    .A1(_17338_),
    .A2(_17340_),
    .ZN(_17341_)
  );
  INV_X1 _52897_ (
    .A(_17341_),
    .ZN(_01383_)
  );
  AND2_X1 _52898_ (
    .A1(_12710_),
    .A2(_13169_),
    .ZN(_17342_)
  );
  INV_X1 _52899_ (
    .A(_17342_),
    .ZN(_17343_)
  );
  AND2_X1 _52900_ (
    .A1(\cpuregs[29] [20]),
    .A2(_12711_),
    .ZN(_17344_)
  );
  INV_X1 _52901_ (
    .A(_17344_),
    .ZN(_17345_)
  );
  AND2_X1 _52902_ (
    .A1(_17343_),
    .A2(_17345_),
    .ZN(_17346_)
  );
  INV_X1 _52903_ (
    .A(_17346_),
    .ZN(_01384_)
  );
  AND2_X1 _52904_ (
    .A1(_12710_),
    .A2(_13184_),
    .ZN(_17347_)
  );
  INV_X1 _52905_ (
    .A(_17347_),
    .ZN(_17348_)
  );
  AND2_X1 _52906_ (
    .A1(\cpuregs[29] [21]),
    .A2(_12711_),
    .ZN(_17349_)
  );
  INV_X1 _52907_ (
    .A(_17349_),
    .ZN(_17350_)
  );
  AND2_X1 _52908_ (
    .A1(_17348_),
    .A2(_17350_),
    .ZN(_17351_)
  );
  INV_X1 _52909_ (
    .A(_17351_),
    .ZN(_01385_)
  );
  AND2_X1 _52910_ (
    .A1(_12710_),
    .A2(_13199_),
    .ZN(_17352_)
  );
  INV_X1 _52911_ (
    .A(_17352_),
    .ZN(_17353_)
  );
  AND2_X1 _52912_ (
    .A1(\cpuregs[29] [22]),
    .A2(_12711_),
    .ZN(_17354_)
  );
  INV_X1 _52913_ (
    .A(_17354_),
    .ZN(_17355_)
  );
  AND2_X1 _52914_ (
    .A1(_17353_),
    .A2(_17355_),
    .ZN(_17356_)
  );
  INV_X1 _52915_ (
    .A(_17356_),
    .ZN(_01386_)
  );
  AND2_X1 _52916_ (
    .A1(_12710_),
    .A2(_13214_),
    .ZN(_17357_)
  );
  INV_X1 _52917_ (
    .A(_17357_),
    .ZN(_17358_)
  );
  AND2_X1 _52918_ (
    .A1(\cpuregs[29] [23]),
    .A2(_12711_),
    .ZN(_17359_)
  );
  INV_X1 _52919_ (
    .A(_17359_),
    .ZN(_17360_)
  );
  AND2_X1 _52920_ (
    .A1(_17358_),
    .A2(_17360_),
    .ZN(_17361_)
  );
  INV_X1 _52921_ (
    .A(_17361_),
    .ZN(_01387_)
  );
  AND2_X1 _52922_ (
    .A1(_12710_),
    .A2(_13229_),
    .ZN(_17362_)
  );
  INV_X1 _52923_ (
    .A(_17362_),
    .ZN(_17363_)
  );
  AND2_X1 _52924_ (
    .A1(\cpuregs[29] [24]),
    .A2(_12711_),
    .ZN(_17364_)
  );
  INV_X1 _52925_ (
    .A(_17364_),
    .ZN(_17365_)
  );
  AND2_X1 _52926_ (
    .A1(_17363_),
    .A2(_17365_),
    .ZN(_17366_)
  );
  INV_X1 _52927_ (
    .A(_17366_),
    .ZN(_01388_)
  );
  AND2_X1 _52928_ (
    .A1(_12710_),
    .A2(_13244_),
    .ZN(_17367_)
  );
  INV_X1 _52929_ (
    .A(_17367_),
    .ZN(_17368_)
  );
  AND2_X1 _52930_ (
    .A1(\cpuregs[29] [25]),
    .A2(_12711_),
    .ZN(_17369_)
  );
  INV_X1 _52931_ (
    .A(_17369_),
    .ZN(_17370_)
  );
  AND2_X1 _52932_ (
    .A1(_17368_),
    .A2(_17370_),
    .ZN(_17371_)
  );
  INV_X1 _52933_ (
    .A(_17371_),
    .ZN(_01389_)
  );
  AND2_X1 _52934_ (
    .A1(_12710_),
    .A2(_13259_),
    .ZN(_17372_)
  );
  INV_X1 _52935_ (
    .A(_17372_),
    .ZN(_17373_)
  );
  AND2_X1 _52936_ (
    .A1(\cpuregs[29] [26]),
    .A2(_12711_),
    .ZN(_17374_)
  );
  INV_X1 _52937_ (
    .A(_17374_),
    .ZN(_17375_)
  );
  AND2_X1 _52938_ (
    .A1(_17373_),
    .A2(_17375_),
    .ZN(_17376_)
  );
  INV_X1 _52939_ (
    .A(_17376_),
    .ZN(_01390_)
  );
  AND2_X1 _52940_ (
    .A1(_12710_),
    .A2(_13274_),
    .ZN(_17377_)
  );
  INV_X1 _52941_ (
    .A(_17377_),
    .ZN(_17378_)
  );
  AND2_X1 _52942_ (
    .A1(\cpuregs[29] [27]),
    .A2(_12711_),
    .ZN(_17379_)
  );
  INV_X1 _52943_ (
    .A(_17379_),
    .ZN(_17380_)
  );
  AND2_X1 _52944_ (
    .A1(_17378_),
    .A2(_17380_),
    .ZN(_17381_)
  );
  INV_X1 _52945_ (
    .A(_17381_),
    .ZN(_01391_)
  );
  AND2_X1 _52946_ (
    .A1(_12710_),
    .A2(_13289_),
    .ZN(_17382_)
  );
  INV_X1 _52947_ (
    .A(_17382_),
    .ZN(_17383_)
  );
  AND2_X1 _52948_ (
    .A1(\cpuregs[29] [28]),
    .A2(_12711_),
    .ZN(_17384_)
  );
  INV_X1 _52949_ (
    .A(_17384_),
    .ZN(_17385_)
  );
  AND2_X1 _52950_ (
    .A1(_17383_),
    .A2(_17385_),
    .ZN(_17386_)
  );
  INV_X1 _52951_ (
    .A(_17386_),
    .ZN(_01392_)
  );
  AND2_X1 _52952_ (
    .A1(_12710_),
    .A2(_13304_),
    .ZN(_17387_)
  );
  INV_X1 _52953_ (
    .A(_17387_),
    .ZN(_17388_)
  );
  AND2_X1 _52954_ (
    .A1(\cpuregs[29] [29]),
    .A2(_12711_),
    .ZN(_17389_)
  );
  INV_X1 _52955_ (
    .A(_17389_),
    .ZN(_17390_)
  );
  AND2_X1 _52956_ (
    .A1(_17388_),
    .A2(_17390_),
    .ZN(_17391_)
  );
  INV_X1 _52957_ (
    .A(_17391_),
    .ZN(_01393_)
  );
  AND2_X1 _52958_ (
    .A1(_12710_),
    .A2(_13319_),
    .ZN(_17392_)
  );
  INV_X1 _52959_ (
    .A(_17392_),
    .ZN(_17393_)
  );
  AND2_X1 _52960_ (
    .A1(\cpuregs[29] [30]),
    .A2(_12711_),
    .ZN(_17394_)
  );
  INV_X1 _52961_ (
    .A(_17394_),
    .ZN(_17395_)
  );
  AND2_X1 _52962_ (
    .A1(_17393_),
    .A2(_17395_),
    .ZN(_17396_)
  );
  INV_X1 _52963_ (
    .A(_17396_),
    .ZN(_01394_)
  );
  AND2_X1 _52964_ (
    .A1(_12717_),
    .A2(_12874_),
    .ZN(_17397_)
  );
  INV_X1 _52965_ (
    .A(_17397_),
    .ZN(_17398_)
  );
  AND2_X1 _52966_ (
    .A1(\cpuregs[28] [0]),
    .A2(_12718_),
    .ZN(_17399_)
  );
  INV_X1 _52967_ (
    .A(_17399_),
    .ZN(_17400_)
  );
  AND2_X1 _52968_ (
    .A1(_17398_),
    .A2(_17400_),
    .ZN(_17401_)
  );
  INV_X1 _52969_ (
    .A(_17401_),
    .ZN(_01395_)
  );
  AND2_X1 _52970_ (
    .A1(_12717_),
    .A2(_12886_),
    .ZN(_17402_)
  );
  INV_X1 _52971_ (
    .A(_17402_),
    .ZN(_17403_)
  );
  AND2_X1 _52972_ (
    .A1(\cpuregs[28] [1]),
    .A2(_12718_),
    .ZN(_17404_)
  );
  INV_X1 _52973_ (
    .A(_17404_),
    .ZN(_17405_)
  );
  AND2_X1 _52974_ (
    .A1(_17403_),
    .A2(_17405_),
    .ZN(_17406_)
  );
  INV_X1 _52975_ (
    .A(_17406_),
    .ZN(_01396_)
  );
  AND2_X1 _52976_ (
    .A1(\cpuregs[28] [2]),
    .A2(_12718_),
    .ZN(_17407_)
  );
  INV_X1 _52977_ (
    .A(_17407_),
    .ZN(_17408_)
  );
  AND2_X1 _52978_ (
    .A1(_12717_),
    .A2(_12900_),
    .ZN(_17409_)
  );
  INV_X1 _52979_ (
    .A(_17409_),
    .ZN(_17410_)
  );
  AND2_X1 _52980_ (
    .A1(_17408_),
    .A2(_17410_),
    .ZN(_17411_)
  );
  INV_X1 _52981_ (
    .A(_17411_),
    .ZN(_01397_)
  );
  AND2_X1 _52982_ (
    .A1(_12717_),
    .A2(_12913_),
    .ZN(_17412_)
  );
  INV_X1 _52983_ (
    .A(_17412_),
    .ZN(_17413_)
  );
  AND2_X1 _52984_ (
    .A1(\cpuregs[28] [3]),
    .A2(_12718_),
    .ZN(_17414_)
  );
  INV_X1 _52985_ (
    .A(_17414_),
    .ZN(_17415_)
  );
  AND2_X1 _52986_ (
    .A1(_17413_),
    .A2(_17415_),
    .ZN(_17416_)
  );
  INV_X1 _52987_ (
    .A(_17416_),
    .ZN(_01398_)
  );
  AND2_X1 _52988_ (
    .A1(_12717_),
    .A2(_12928_),
    .ZN(_17417_)
  );
  INV_X1 _52989_ (
    .A(_17417_),
    .ZN(_17418_)
  );
  AND2_X1 _52990_ (
    .A1(\cpuregs[28] [4]),
    .A2(_12718_),
    .ZN(_17419_)
  );
  INV_X1 _52991_ (
    .A(_17419_),
    .ZN(_17420_)
  );
  AND2_X1 _52992_ (
    .A1(_17418_),
    .A2(_17420_),
    .ZN(_17421_)
  );
  INV_X1 _52993_ (
    .A(_17421_),
    .ZN(_01399_)
  );
  AND2_X1 _52994_ (
    .A1(_12717_),
    .A2(_12943_),
    .ZN(_17422_)
  );
  INV_X1 _52995_ (
    .A(_17422_),
    .ZN(_17423_)
  );
  AND2_X1 _52996_ (
    .A1(\cpuregs[28] [5]),
    .A2(_12718_),
    .ZN(_17424_)
  );
  INV_X1 _52997_ (
    .A(_17424_),
    .ZN(_17425_)
  );
  AND2_X1 _52998_ (
    .A1(_17423_),
    .A2(_17425_),
    .ZN(_17426_)
  );
  INV_X1 _52999_ (
    .A(_17426_),
    .ZN(_01400_)
  );
  AND2_X1 _53000_ (
    .A1(_12717_),
    .A2(_12958_),
    .ZN(_17427_)
  );
  INV_X1 _53001_ (
    .A(_17427_),
    .ZN(_17428_)
  );
  AND2_X1 _53002_ (
    .A1(\cpuregs[28] [6]),
    .A2(_12718_),
    .ZN(_17429_)
  );
  INV_X1 _53003_ (
    .A(_17429_),
    .ZN(_17430_)
  );
  AND2_X1 _53004_ (
    .A1(_17428_),
    .A2(_17430_),
    .ZN(_17431_)
  );
  INV_X1 _53005_ (
    .A(_17431_),
    .ZN(_01401_)
  );
  AND2_X1 _53006_ (
    .A1(_12717_),
    .A2(_12973_),
    .ZN(_17432_)
  );
  INV_X1 _53007_ (
    .A(_17432_),
    .ZN(_17433_)
  );
  AND2_X1 _53008_ (
    .A1(\cpuregs[28] [7]),
    .A2(_12718_),
    .ZN(_17434_)
  );
  INV_X1 _53009_ (
    .A(_17434_),
    .ZN(_17435_)
  );
  AND2_X1 _53010_ (
    .A1(_17433_),
    .A2(_17435_),
    .ZN(_17436_)
  );
  INV_X1 _53011_ (
    .A(_17436_),
    .ZN(_01402_)
  );
  AND2_X1 _53012_ (
    .A1(_12717_),
    .A2(_12988_),
    .ZN(_17437_)
  );
  INV_X1 _53013_ (
    .A(_17437_),
    .ZN(_17438_)
  );
  AND2_X1 _53014_ (
    .A1(\cpuregs[28] [8]),
    .A2(_12718_),
    .ZN(_17439_)
  );
  INV_X1 _53015_ (
    .A(_17439_),
    .ZN(_17440_)
  );
  AND2_X1 _53016_ (
    .A1(_17438_),
    .A2(_17440_),
    .ZN(_17441_)
  );
  INV_X1 _53017_ (
    .A(_17441_),
    .ZN(_01403_)
  );
  AND2_X1 _53018_ (
    .A1(_12717_),
    .A2(_13003_),
    .ZN(_17442_)
  );
  INV_X1 _53019_ (
    .A(_17442_),
    .ZN(_17443_)
  );
  AND2_X1 _53020_ (
    .A1(\cpuregs[28] [9]),
    .A2(_12718_),
    .ZN(_17444_)
  );
  INV_X1 _53021_ (
    .A(_17444_),
    .ZN(_17445_)
  );
  AND2_X1 _53022_ (
    .A1(_17443_),
    .A2(_17445_),
    .ZN(_17446_)
  );
  INV_X1 _53023_ (
    .A(_17446_),
    .ZN(_01404_)
  );
  AND2_X1 _53024_ (
    .A1(_12717_),
    .A2(_13018_),
    .ZN(_17447_)
  );
  INV_X1 _53025_ (
    .A(_17447_),
    .ZN(_17448_)
  );
  AND2_X1 _53026_ (
    .A1(\cpuregs[28] [10]),
    .A2(_12718_),
    .ZN(_17449_)
  );
  INV_X1 _53027_ (
    .A(_17449_),
    .ZN(_17450_)
  );
  AND2_X1 _53028_ (
    .A1(_17448_),
    .A2(_17450_),
    .ZN(_17451_)
  );
  INV_X1 _53029_ (
    .A(_17451_),
    .ZN(_01405_)
  );
  AND2_X1 _53030_ (
    .A1(_12717_),
    .A2(_13033_),
    .ZN(_17452_)
  );
  INV_X1 _53031_ (
    .A(_17452_),
    .ZN(_17453_)
  );
  AND2_X1 _53032_ (
    .A1(\cpuregs[28] [11]),
    .A2(_12718_),
    .ZN(_17454_)
  );
  INV_X1 _53033_ (
    .A(_17454_),
    .ZN(_17455_)
  );
  AND2_X1 _53034_ (
    .A1(_17453_),
    .A2(_17455_),
    .ZN(_17456_)
  );
  INV_X1 _53035_ (
    .A(_17456_),
    .ZN(_01406_)
  );
  AND2_X1 _53036_ (
    .A1(_12717_),
    .A2(_13048_),
    .ZN(_17457_)
  );
  INV_X1 _53037_ (
    .A(_17457_),
    .ZN(_17458_)
  );
  AND2_X1 _53038_ (
    .A1(\cpuregs[28] [12]),
    .A2(_12718_),
    .ZN(_17459_)
  );
  INV_X1 _53039_ (
    .A(_17459_),
    .ZN(_17460_)
  );
  AND2_X1 _53040_ (
    .A1(_17458_),
    .A2(_17460_),
    .ZN(_17461_)
  );
  INV_X1 _53041_ (
    .A(_17461_),
    .ZN(_01407_)
  );
  AND2_X1 _53042_ (
    .A1(_12717_),
    .A2(_13063_),
    .ZN(_17462_)
  );
  INV_X1 _53043_ (
    .A(_17462_),
    .ZN(_17463_)
  );
  AND2_X1 _53044_ (
    .A1(\cpuregs[28] [13]),
    .A2(_12718_),
    .ZN(_17464_)
  );
  INV_X1 _53045_ (
    .A(_17464_),
    .ZN(_17465_)
  );
  AND2_X1 _53046_ (
    .A1(_17463_),
    .A2(_17465_),
    .ZN(_17466_)
  );
  INV_X1 _53047_ (
    .A(_17466_),
    .ZN(_01408_)
  );
  AND2_X1 _53048_ (
    .A1(_12717_),
    .A2(_13078_),
    .ZN(_17467_)
  );
  INV_X1 _53049_ (
    .A(_17467_),
    .ZN(_17468_)
  );
  AND2_X1 _53050_ (
    .A1(\cpuregs[28] [14]),
    .A2(_12718_),
    .ZN(_17469_)
  );
  INV_X1 _53051_ (
    .A(_17469_),
    .ZN(_17470_)
  );
  AND2_X1 _53052_ (
    .A1(_17468_),
    .A2(_17470_),
    .ZN(_17471_)
  );
  INV_X1 _53053_ (
    .A(_17471_),
    .ZN(_01409_)
  );
  AND2_X1 _53054_ (
    .A1(_12717_),
    .A2(_13093_),
    .ZN(_17472_)
  );
  INV_X1 _53055_ (
    .A(_17472_),
    .ZN(_17473_)
  );
  AND2_X1 _53056_ (
    .A1(\cpuregs[28] [15]),
    .A2(_12718_),
    .ZN(_17474_)
  );
  INV_X1 _53057_ (
    .A(_17474_),
    .ZN(_17475_)
  );
  AND2_X1 _53058_ (
    .A1(_17473_),
    .A2(_17475_),
    .ZN(_17476_)
  );
  INV_X1 _53059_ (
    .A(_17476_),
    .ZN(_01410_)
  );
  AND2_X1 _53060_ (
    .A1(\cpuregs[28] [16]),
    .A2(_12718_),
    .ZN(_17477_)
  );
  INV_X1 _53061_ (
    .A(_17477_),
    .ZN(_17478_)
  );
  AND2_X1 _53062_ (
    .A1(_12717_),
    .A2(_13108_),
    .ZN(_17479_)
  );
  INV_X1 _53063_ (
    .A(_17479_),
    .ZN(_17480_)
  );
  AND2_X1 _53064_ (
    .A1(_17478_),
    .A2(_17480_),
    .ZN(_17481_)
  );
  INV_X1 _53065_ (
    .A(_17481_),
    .ZN(_01411_)
  );
  AND2_X1 _53066_ (
    .A1(_12717_),
    .A2(_13123_),
    .ZN(_17482_)
  );
  INV_X1 _53067_ (
    .A(_17482_),
    .ZN(_17483_)
  );
  AND2_X1 _53068_ (
    .A1(\cpuregs[28] [17]),
    .A2(_12718_),
    .ZN(_17484_)
  );
  INV_X1 _53069_ (
    .A(_17484_),
    .ZN(_17485_)
  );
  AND2_X1 _53070_ (
    .A1(_17483_),
    .A2(_17485_),
    .ZN(_17486_)
  );
  INV_X1 _53071_ (
    .A(_17486_),
    .ZN(_01412_)
  );
  AND2_X1 _53072_ (
    .A1(_12717_),
    .A2(_13139_),
    .ZN(_17487_)
  );
  INV_X1 _53073_ (
    .A(_17487_),
    .ZN(_17488_)
  );
  AND2_X1 _53074_ (
    .A1(\cpuregs[28] [18]),
    .A2(_12718_),
    .ZN(_17489_)
  );
  INV_X1 _53075_ (
    .A(_17489_),
    .ZN(_17490_)
  );
  AND2_X1 _53076_ (
    .A1(_17488_),
    .A2(_17490_),
    .ZN(_17491_)
  );
  INV_X1 _53077_ (
    .A(_17491_),
    .ZN(_01413_)
  );
  AND2_X1 _53078_ (
    .A1(_12717_),
    .A2(_13154_),
    .ZN(_17492_)
  );
  INV_X1 _53079_ (
    .A(_17492_),
    .ZN(_17493_)
  );
  AND2_X1 _53080_ (
    .A1(\cpuregs[28] [19]),
    .A2(_12718_),
    .ZN(_17494_)
  );
  INV_X1 _53081_ (
    .A(_17494_),
    .ZN(_17495_)
  );
  AND2_X1 _53082_ (
    .A1(_17493_),
    .A2(_17495_),
    .ZN(_17496_)
  );
  INV_X1 _53083_ (
    .A(_17496_),
    .ZN(_01414_)
  );
  AND2_X1 _53084_ (
    .A1(_12717_),
    .A2(_13169_),
    .ZN(_17497_)
  );
  INV_X1 _53085_ (
    .A(_17497_),
    .ZN(_17498_)
  );
  AND2_X1 _53086_ (
    .A1(\cpuregs[28] [20]),
    .A2(_12718_),
    .ZN(_17499_)
  );
  INV_X1 _53087_ (
    .A(_17499_),
    .ZN(_17500_)
  );
  AND2_X1 _53088_ (
    .A1(_17498_),
    .A2(_17500_),
    .ZN(_17501_)
  );
  INV_X1 _53089_ (
    .A(_17501_),
    .ZN(_01415_)
  );
  AND2_X1 _53090_ (
    .A1(_12717_),
    .A2(_13184_),
    .ZN(_17502_)
  );
  INV_X1 _53091_ (
    .A(_17502_),
    .ZN(_17503_)
  );
  AND2_X1 _53092_ (
    .A1(\cpuregs[28] [21]),
    .A2(_12718_),
    .ZN(_17504_)
  );
  INV_X1 _53093_ (
    .A(_17504_),
    .ZN(_17505_)
  );
  AND2_X1 _53094_ (
    .A1(_17503_),
    .A2(_17505_),
    .ZN(_17506_)
  );
  INV_X1 _53095_ (
    .A(_17506_),
    .ZN(_01416_)
  );
  AND2_X1 _53096_ (
    .A1(_12717_),
    .A2(_13199_),
    .ZN(_17507_)
  );
  INV_X1 _53097_ (
    .A(_17507_),
    .ZN(_17508_)
  );
  AND2_X1 _53098_ (
    .A1(\cpuregs[28] [22]),
    .A2(_12718_),
    .ZN(_17509_)
  );
  INV_X1 _53099_ (
    .A(_17509_),
    .ZN(_17510_)
  );
  AND2_X1 _53100_ (
    .A1(_17508_),
    .A2(_17510_),
    .ZN(_17511_)
  );
  INV_X1 _53101_ (
    .A(_17511_),
    .ZN(_01417_)
  );
  AND2_X1 _53102_ (
    .A1(_12717_),
    .A2(_13214_),
    .ZN(_17512_)
  );
  INV_X1 _53103_ (
    .A(_17512_),
    .ZN(_17513_)
  );
  AND2_X1 _53104_ (
    .A1(\cpuregs[28] [23]),
    .A2(_12718_),
    .ZN(_17514_)
  );
  INV_X1 _53105_ (
    .A(_17514_),
    .ZN(_17515_)
  );
  AND2_X1 _53106_ (
    .A1(_17513_),
    .A2(_17515_),
    .ZN(_17516_)
  );
  INV_X1 _53107_ (
    .A(_17516_),
    .ZN(_01418_)
  );
  AND2_X1 _53108_ (
    .A1(_12717_),
    .A2(_13229_),
    .ZN(_17517_)
  );
  INV_X1 _53109_ (
    .A(_17517_),
    .ZN(_17518_)
  );
  AND2_X1 _53110_ (
    .A1(\cpuregs[28] [24]),
    .A2(_12718_),
    .ZN(_17519_)
  );
  INV_X1 _53111_ (
    .A(_17519_),
    .ZN(_17520_)
  );
  AND2_X1 _53112_ (
    .A1(_17518_),
    .A2(_17520_),
    .ZN(_17521_)
  );
  INV_X1 _53113_ (
    .A(_17521_),
    .ZN(_01419_)
  );
  AND2_X1 _53114_ (
    .A1(_12717_),
    .A2(_13244_),
    .ZN(_17522_)
  );
  INV_X1 _53115_ (
    .A(_17522_),
    .ZN(_17523_)
  );
  AND2_X1 _53116_ (
    .A1(\cpuregs[28] [25]),
    .A2(_12718_),
    .ZN(_17524_)
  );
  INV_X1 _53117_ (
    .A(_17524_),
    .ZN(_17525_)
  );
  AND2_X1 _53118_ (
    .A1(_17523_),
    .A2(_17525_),
    .ZN(_17526_)
  );
  INV_X1 _53119_ (
    .A(_17526_),
    .ZN(_01420_)
  );
  AND2_X1 _53120_ (
    .A1(_12717_),
    .A2(_13259_),
    .ZN(_17527_)
  );
  INV_X1 _53121_ (
    .A(_17527_),
    .ZN(_17528_)
  );
  AND2_X1 _53122_ (
    .A1(\cpuregs[28] [26]),
    .A2(_12718_),
    .ZN(_17529_)
  );
  INV_X1 _53123_ (
    .A(_17529_),
    .ZN(_17530_)
  );
  AND2_X1 _53124_ (
    .A1(_17528_),
    .A2(_17530_),
    .ZN(_17531_)
  );
  INV_X1 _53125_ (
    .A(_17531_),
    .ZN(_01421_)
  );
  AND2_X1 _53126_ (
    .A1(_12717_),
    .A2(_13274_),
    .ZN(_17532_)
  );
  INV_X1 _53127_ (
    .A(_17532_),
    .ZN(_17533_)
  );
  AND2_X1 _53128_ (
    .A1(\cpuregs[28] [27]),
    .A2(_12718_),
    .ZN(_17534_)
  );
  INV_X1 _53129_ (
    .A(_17534_),
    .ZN(_17535_)
  );
  AND2_X1 _53130_ (
    .A1(_17533_),
    .A2(_17535_),
    .ZN(_17536_)
  );
  INV_X1 _53131_ (
    .A(_17536_),
    .ZN(_01422_)
  );
  AND2_X1 _53132_ (
    .A1(_12717_),
    .A2(_13289_),
    .ZN(_17537_)
  );
  INV_X1 _53133_ (
    .A(_17537_),
    .ZN(_17538_)
  );
  AND2_X1 _53134_ (
    .A1(\cpuregs[28] [28]),
    .A2(_12718_),
    .ZN(_17539_)
  );
  INV_X1 _53135_ (
    .A(_17539_),
    .ZN(_17540_)
  );
  AND2_X1 _53136_ (
    .A1(_17538_),
    .A2(_17540_),
    .ZN(_17541_)
  );
  INV_X1 _53137_ (
    .A(_17541_),
    .ZN(_01423_)
  );
  AND2_X1 _53138_ (
    .A1(_12717_),
    .A2(_13304_),
    .ZN(_17542_)
  );
  INV_X1 _53139_ (
    .A(_17542_),
    .ZN(_17543_)
  );
  AND2_X1 _53140_ (
    .A1(\cpuregs[28] [29]),
    .A2(_12718_),
    .ZN(_17544_)
  );
  INV_X1 _53141_ (
    .A(_17544_),
    .ZN(_17545_)
  );
  AND2_X1 _53142_ (
    .A1(_17543_),
    .A2(_17545_),
    .ZN(_17546_)
  );
  INV_X1 _53143_ (
    .A(_17546_),
    .ZN(_01424_)
  );
  AND2_X1 _53144_ (
    .A1(_12717_),
    .A2(_13319_),
    .ZN(_17547_)
  );
  INV_X1 _53145_ (
    .A(_17547_),
    .ZN(_17548_)
  );
  AND2_X1 _53146_ (
    .A1(\cpuregs[28] [30]),
    .A2(_12718_),
    .ZN(_17549_)
  );
  INV_X1 _53147_ (
    .A(_17549_),
    .ZN(_17550_)
  );
  AND2_X1 _53148_ (
    .A1(_17548_),
    .A2(_17550_),
    .ZN(_17551_)
  );
  INV_X1 _53149_ (
    .A(_17551_),
    .ZN(_01425_)
  );
  AND2_X1 _53150_ (
    .A1(_12725_),
    .A2(_12874_),
    .ZN(_17552_)
  );
  INV_X1 _53151_ (
    .A(_17552_),
    .ZN(_17553_)
  );
  AND2_X1 _53152_ (
    .A1(\cpuregs[27] [0]),
    .A2(_12726_),
    .ZN(_17554_)
  );
  INV_X1 _53153_ (
    .A(_17554_),
    .ZN(_17555_)
  );
  AND2_X1 _53154_ (
    .A1(_17553_),
    .A2(_17555_),
    .ZN(_17556_)
  );
  INV_X1 _53155_ (
    .A(_17556_),
    .ZN(_01426_)
  );
  AND2_X1 _53156_ (
    .A1(_12725_),
    .A2(_12886_),
    .ZN(_17557_)
  );
  INV_X1 _53157_ (
    .A(_17557_),
    .ZN(_17558_)
  );
  AND2_X1 _53158_ (
    .A1(\cpuregs[27] [1]),
    .A2(_12726_),
    .ZN(_17559_)
  );
  INV_X1 _53159_ (
    .A(_17559_),
    .ZN(_17560_)
  );
  AND2_X1 _53160_ (
    .A1(_17558_),
    .A2(_17560_),
    .ZN(_17561_)
  );
  INV_X1 _53161_ (
    .A(_17561_),
    .ZN(_01427_)
  );
  AND2_X1 _53162_ (
    .A1(_12725_),
    .A2(_12900_),
    .ZN(_17562_)
  );
  INV_X1 _53163_ (
    .A(_17562_),
    .ZN(_17563_)
  );
  AND2_X1 _53164_ (
    .A1(\cpuregs[27] [2]),
    .A2(_12726_),
    .ZN(_17564_)
  );
  INV_X1 _53165_ (
    .A(_17564_),
    .ZN(_17565_)
  );
  AND2_X1 _53166_ (
    .A1(_17563_),
    .A2(_17565_),
    .ZN(_17566_)
  );
  INV_X1 _53167_ (
    .A(_17566_),
    .ZN(_01428_)
  );
  AND2_X1 _53168_ (
    .A1(_12725_),
    .A2(_12913_),
    .ZN(_17567_)
  );
  INV_X1 _53169_ (
    .A(_17567_),
    .ZN(_17568_)
  );
  AND2_X1 _53170_ (
    .A1(\cpuregs[27] [3]),
    .A2(_12726_),
    .ZN(_17569_)
  );
  INV_X1 _53171_ (
    .A(_17569_),
    .ZN(_17570_)
  );
  AND2_X1 _53172_ (
    .A1(_17568_),
    .A2(_17570_),
    .ZN(_17571_)
  );
  INV_X1 _53173_ (
    .A(_17571_),
    .ZN(_01429_)
  );
  AND2_X1 _53174_ (
    .A1(_12725_),
    .A2(_12928_),
    .ZN(_17572_)
  );
  INV_X1 _53175_ (
    .A(_17572_),
    .ZN(_17573_)
  );
  AND2_X1 _53176_ (
    .A1(\cpuregs[27] [4]),
    .A2(_12726_),
    .ZN(_17574_)
  );
  INV_X1 _53177_ (
    .A(_17574_),
    .ZN(_17575_)
  );
  AND2_X1 _53178_ (
    .A1(_17573_),
    .A2(_17575_),
    .ZN(_17576_)
  );
  INV_X1 _53179_ (
    .A(_17576_),
    .ZN(_01430_)
  );
  AND2_X1 _53180_ (
    .A1(_12725_),
    .A2(_12943_),
    .ZN(_17577_)
  );
  INV_X1 _53181_ (
    .A(_17577_),
    .ZN(_17578_)
  );
  AND2_X1 _53182_ (
    .A1(\cpuregs[27] [5]),
    .A2(_12726_),
    .ZN(_17579_)
  );
  INV_X1 _53183_ (
    .A(_17579_),
    .ZN(_17580_)
  );
  AND2_X1 _53184_ (
    .A1(_17578_),
    .A2(_17580_),
    .ZN(_17581_)
  );
  INV_X1 _53185_ (
    .A(_17581_),
    .ZN(_01431_)
  );
  AND2_X1 _53186_ (
    .A1(_12725_),
    .A2(_12958_),
    .ZN(_17582_)
  );
  INV_X1 _53187_ (
    .A(_17582_),
    .ZN(_17583_)
  );
  AND2_X1 _53188_ (
    .A1(\cpuregs[27] [6]),
    .A2(_12726_),
    .ZN(_17584_)
  );
  INV_X1 _53189_ (
    .A(_17584_),
    .ZN(_17585_)
  );
  AND2_X1 _53190_ (
    .A1(_17583_),
    .A2(_17585_),
    .ZN(_17586_)
  );
  INV_X1 _53191_ (
    .A(_17586_),
    .ZN(_01432_)
  );
  AND2_X1 _53192_ (
    .A1(_12725_),
    .A2(_12973_),
    .ZN(_17587_)
  );
  INV_X1 _53193_ (
    .A(_17587_),
    .ZN(_17588_)
  );
  AND2_X1 _53194_ (
    .A1(\cpuregs[27] [7]),
    .A2(_12726_),
    .ZN(_17589_)
  );
  INV_X1 _53195_ (
    .A(_17589_),
    .ZN(_17590_)
  );
  AND2_X1 _53196_ (
    .A1(_17588_),
    .A2(_17590_),
    .ZN(_17591_)
  );
  INV_X1 _53197_ (
    .A(_17591_),
    .ZN(_01433_)
  );
  AND2_X1 _53198_ (
    .A1(_12725_),
    .A2(_12988_),
    .ZN(_17592_)
  );
  INV_X1 _53199_ (
    .A(_17592_),
    .ZN(_17593_)
  );
  AND2_X1 _53200_ (
    .A1(\cpuregs[27] [8]),
    .A2(_12726_),
    .ZN(_17594_)
  );
  INV_X1 _53201_ (
    .A(_17594_),
    .ZN(_17595_)
  );
  AND2_X1 _53202_ (
    .A1(_17593_),
    .A2(_17595_),
    .ZN(_17596_)
  );
  INV_X1 _53203_ (
    .A(_17596_),
    .ZN(_01434_)
  );
  AND2_X1 _53204_ (
    .A1(_12725_),
    .A2(_13003_),
    .ZN(_17597_)
  );
  INV_X1 _53205_ (
    .A(_17597_),
    .ZN(_17598_)
  );
  AND2_X1 _53206_ (
    .A1(\cpuregs[27] [9]),
    .A2(_12726_),
    .ZN(_17599_)
  );
  INV_X1 _53207_ (
    .A(_17599_),
    .ZN(_17600_)
  );
  AND2_X1 _53208_ (
    .A1(_17598_),
    .A2(_17600_),
    .ZN(_17601_)
  );
  INV_X1 _53209_ (
    .A(_17601_),
    .ZN(_01435_)
  );
  AND2_X1 _53210_ (
    .A1(_12725_),
    .A2(_13018_),
    .ZN(_17602_)
  );
  INV_X1 _53211_ (
    .A(_17602_),
    .ZN(_17603_)
  );
  AND2_X1 _53212_ (
    .A1(\cpuregs[27] [10]),
    .A2(_12726_),
    .ZN(_17604_)
  );
  INV_X1 _53213_ (
    .A(_17604_),
    .ZN(_17605_)
  );
  AND2_X1 _53214_ (
    .A1(_17603_),
    .A2(_17605_),
    .ZN(_17606_)
  );
  INV_X1 _53215_ (
    .A(_17606_),
    .ZN(_01436_)
  );
  AND2_X1 _53216_ (
    .A1(_12725_),
    .A2(_13033_),
    .ZN(_17607_)
  );
  INV_X1 _53217_ (
    .A(_17607_),
    .ZN(_17608_)
  );
  AND2_X1 _53218_ (
    .A1(\cpuregs[27] [11]),
    .A2(_12726_),
    .ZN(_17609_)
  );
  INV_X1 _53219_ (
    .A(_17609_),
    .ZN(_17610_)
  );
  AND2_X1 _53220_ (
    .A1(_17608_),
    .A2(_17610_),
    .ZN(_17611_)
  );
  INV_X1 _53221_ (
    .A(_17611_),
    .ZN(_01437_)
  );
  AND2_X1 _53222_ (
    .A1(_12725_),
    .A2(_13048_),
    .ZN(_17612_)
  );
  INV_X1 _53223_ (
    .A(_17612_),
    .ZN(_17613_)
  );
  AND2_X1 _53224_ (
    .A1(\cpuregs[27] [12]),
    .A2(_12726_),
    .ZN(_17614_)
  );
  INV_X1 _53225_ (
    .A(_17614_),
    .ZN(_17615_)
  );
  AND2_X1 _53226_ (
    .A1(_17613_),
    .A2(_17615_),
    .ZN(_17616_)
  );
  INV_X1 _53227_ (
    .A(_17616_),
    .ZN(_01438_)
  );
  AND2_X1 _53228_ (
    .A1(_12725_),
    .A2(_13063_),
    .ZN(_17617_)
  );
  INV_X1 _53229_ (
    .A(_17617_),
    .ZN(_17618_)
  );
  AND2_X1 _53230_ (
    .A1(\cpuregs[27] [13]),
    .A2(_12726_),
    .ZN(_17619_)
  );
  INV_X1 _53231_ (
    .A(_17619_),
    .ZN(_17620_)
  );
  AND2_X1 _53232_ (
    .A1(_17618_),
    .A2(_17620_),
    .ZN(_17621_)
  );
  INV_X1 _53233_ (
    .A(_17621_),
    .ZN(_01439_)
  );
  AND2_X1 _53234_ (
    .A1(_12725_),
    .A2(_13078_),
    .ZN(_17622_)
  );
  INV_X1 _53235_ (
    .A(_17622_),
    .ZN(_17623_)
  );
  AND2_X1 _53236_ (
    .A1(\cpuregs[27] [14]),
    .A2(_12726_),
    .ZN(_17624_)
  );
  INV_X1 _53237_ (
    .A(_17624_),
    .ZN(_17625_)
  );
  AND2_X1 _53238_ (
    .A1(_17623_),
    .A2(_17625_),
    .ZN(_17626_)
  );
  INV_X1 _53239_ (
    .A(_17626_),
    .ZN(_01440_)
  );
  AND2_X1 _53240_ (
    .A1(_12725_),
    .A2(_13093_),
    .ZN(_17627_)
  );
  INV_X1 _53241_ (
    .A(_17627_),
    .ZN(_17628_)
  );
  AND2_X1 _53242_ (
    .A1(\cpuregs[27] [15]),
    .A2(_12726_),
    .ZN(_17629_)
  );
  INV_X1 _53243_ (
    .A(_17629_),
    .ZN(_17630_)
  );
  AND2_X1 _53244_ (
    .A1(_17628_),
    .A2(_17630_),
    .ZN(_17631_)
  );
  INV_X1 _53245_ (
    .A(_17631_),
    .ZN(_01441_)
  );
  AND2_X1 _53246_ (
    .A1(_12725_),
    .A2(_13108_),
    .ZN(_17632_)
  );
  INV_X1 _53247_ (
    .A(_17632_),
    .ZN(_17633_)
  );
  AND2_X1 _53248_ (
    .A1(\cpuregs[27] [16]),
    .A2(_12726_),
    .ZN(_17634_)
  );
  INV_X1 _53249_ (
    .A(_17634_),
    .ZN(_17635_)
  );
  AND2_X1 _53250_ (
    .A1(_17633_),
    .A2(_17635_),
    .ZN(_17636_)
  );
  INV_X1 _53251_ (
    .A(_17636_),
    .ZN(_01442_)
  );
  AND2_X1 _53252_ (
    .A1(_12725_),
    .A2(_13123_),
    .ZN(_17637_)
  );
  INV_X1 _53253_ (
    .A(_17637_),
    .ZN(_17638_)
  );
  AND2_X1 _53254_ (
    .A1(\cpuregs[27] [17]),
    .A2(_12726_),
    .ZN(_17639_)
  );
  INV_X1 _53255_ (
    .A(_17639_),
    .ZN(_17640_)
  );
  AND2_X1 _53256_ (
    .A1(_17638_),
    .A2(_17640_),
    .ZN(_17641_)
  );
  INV_X1 _53257_ (
    .A(_17641_),
    .ZN(_01443_)
  );
  AND2_X1 _53258_ (
    .A1(_12725_),
    .A2(_13139_),
    .ZN(_17642_)
  );
  INV_X1 _53259_ (
    .A(_17642_),
    .ZN(_17643_)
  );
  AND2_X1 _53260_ (
    .A1(\cpuregs[27] [18]),
    .A2(_12726_),
    .ZN(_17644_)
  );
  INV_X1 _53261_ (
    .A(_17644_),
    .ZN(_17645_)
  );
  AND2_X1 _53262_ (
    .A1(_17643_),
    .A2(_17645_),
    .ZN(_17646_)
  );
  INV_X1 _53263_ (
    .A(_17646_),
    .ZN(_01444_)
  );
  AND2_X1 _53264_ (
    .A1(_12725_),
    .A2(_13154_),
    .ZN(_17647_)
  );
  INV_X1 _53265_ (
    .A(_17647_),
    .ZN(_17648_)
  );
  AND2_X1 _53266_ (
    .A1(\cpuregs[27] [19]),
    .A2(_12726_),
    .ZN(_17649_)
  );
  INV_X1 _53267_ (
    .A(_17649_),
    .ZN(_17650_)
  );
  AND2_X1 _53268_ (
    .A1(_17648_),
    .A2(_17650_),
    .ZN(_17651_)
  );
  INV_X1 _53269_ (
    .A(_17651_),
    .ZN(_01445_)
  );
  AND2_X1 _53270_ (
    .A1(_12725_),
    .A2(_13169_),
    .ZN(_17652_)
  );
  INV_X1 _53271_ (
    .A(_17652_),
    .ZN(_17653_)
  );
  AND2_X1 _53272_ (
    .A1(\cpuregs[27] [20]),
    .A2(_12726_),
    .ZN(_17654_)
  );
  INV_X1 _53273_ (
    .A(_17654_),
    .ZN(_17655_)
  );
  AND2_X1 _53274_ (
    .A1(_17653_),
    .A2(_17655_),
    .ZN(_17656_)
  );
  INV_X1 _53275_ (
    .A(_17656_),
    .ZN(_01446_)
  );
  AND2_X1 _53276_ (
    .A1(_12725_),
    .A2(_13184_),
    .ZN(_17657_)
  );
  INV_X1 _53277_ (
    .A(_17657_),
    .ZN(_17658_)
  );
  AND2_X1 _53278_ (
    .A1(\cpuregs[27] [21]),
    .A2(_12726_),
    .ZN(_17659_)
  );
  INV_X1 _53279_ (
    .A(_17659_),
    .ZN(_17660_)
  );
  AND2_X1 _53280_ (
    .A1(_17658_),
    .A2(_17660_),
    .ZN(_17661_)
  );
  INV_X1 _53281_ (
    .A(_17661_),
    .ZN(_01447_)
  );
  AND2_X1 _53282_ (
    .A1(_12725_),
    .A2(_13199_),
    .ZN(_17662_)
  );
  INV_X1 _53283_ (
    .A(_17662_),
    .ZN(_17663_)
  );
  AND2_X1 _53284_ (
    .A1(\cpuregs[27] [22]),
    .A2(_12726_),
    .ZN(_17664_)
  );
  INV_X1 _53285_ (
    .A(_17664_),
    .ZN(_17665_)
  );
  AND2_X1 _53286_ (
    .A1(_17663_),
    .A2(_17665_),
    .ZN(_17666_)
  );
  INV_X1 _53287_ (
    .A(_17666_),
    .ZN(_01448_)
  );
  AND2_X1 _53288_ (
    .A1(_12725_),
    .A2(_13214_),
    .ZN(_17667_)
  );
  INV_X1 _53289_ (
    .A(_17667_),
    .ZN(_17668_)
  );
  AND2_X1 _53290_ (
    .A1(\cpuregs[27] [23]),
    .A2(_12726_),
    .ZN(_17669_)
  );
  INV_X1 _53291_ (
    .A(_17669_),
    .ZN(_17670_)
  );
  AND2_X1 _53292_ (
    .A1(_17668_),
    .A2(_17670_),
    .ZN(_17671_)
  );
  INV_X1 _53293_ (
    .A(_17671_),
    .ZN(_01449_)
  );
  AND2_X1 _53294_ (
    .A1(_12725_),
    .A2(_13229_),
    .ZN(_17672_)
  );
  INV_X1 _53295_ (
    .A(_17672_),
    .ZN(_17673_)
  );
  AND2_X1 _53296_ (
    .A1(\cpuregs[27] [24]),
    .A2(_12726_),
    .ZN(_17674_)
  );
  INV_X1 _53297_ (
    .A(_17674_),
    .ZN(_17675_)
  );
  AND2_X1 _53298_ (
    .A1(_17673_),
    .A2(_17675_),
    .ZN(_17676_)
  );
  INV_X1 _53299_ (
    .A(_17676_),
    .ZN(_01450_)
  );
  AND2_X1 _53300_ (
    .A1(_12725_),
    .A2(_13244_),
    .ZN(_17677_)
  );
  INV_X1 _53301_ (
    .A(_17677_),
    .ZN(_17678_)
  );
  AND2_X1 _53302_ (
    .A1(\cpuregs[27] [25]),
    .A2(_12726_),
    .ZN(_17679_)
  );
  INV_X1 _53303_ (
    .A(_17679_),
    .ZN(_17680_)
  );
  AND2_X1 _53304_ (
    .A1(_17678_),
    .A2(_17680_),
    .ZN(_17681_)
  );
  INV_X1 _53305_ (
    .A(_17681_),
    .ZN(_01451_)
  );
  AND2_X1 _53306_ (
    .A1(_12725_),
    .A2(_13259_),
    .ZN(_17682_)
  );
  INV_X1 _53307_ (
    .A(_17682_),
    .ZN(_17683_)
  );
  AND2_X1 _53308_ (
    .A1(\cpuregs[27] [26]),
    .A2(_12726_),
    .ZN(_17684_)
  );
  INV_X1 _53309_ (
    .A(_17684_),
    .ZN(_17685_)
  );
  AND2_X1 _53310_ (
    .A1(_17683_),
    .A2(_17685_),
    .ZN(_17686_)
  );
  INV_X1 _53311_ (
    .A(_17686_),
    .ZN(_01452_)
  );
  AND2_X1 _53312_ (
    .A1(_12725_),
    .A2(_13274_),
    .ZN(_17687_)
  );
  INV_X1 _53313_ (
    .A(_17687_),
    .ZN(_17688_)
  );
  AND2_X1 _53314_ (
    .A1(\cpuregs[27] [27]),
    .A2(_12726_),
    .ZN(_17689_)
  );
  INV_X1 _53315_ (
    .A(_17689_),
    .ZN(_17690_)
  );
  AND2_X1 _53316_ (
    .A1(_17688_),
    .A2(_17690_),
    .ZN(_17691_)
  );
  INV_X1 _53317_ (
    .A(_17691_),
    .ZN(_01453_)
  );
  AND2_X1 _53318_ (
    .A1(_12725_),
    .A2(_13289_),
    .ZN(_17692_)
  );
  INV_X1 _53319_ (
    .A(_17692_),
    .ZN(_17693_)
  );
  AND2_X1 _53320_ (
    .A1(\cpuregs[27] [28]),
    .A2(_12726_),
    .ZN(_17694_)
  );
  INV_X1 _53321_ (
    .A(_17694_),
    .ZN(_17695_)
  );
  AND2_X1 _53322_ (
    .A1(_17693_),
    .A2(_17695_),
    .ZN(_17696_)
  );
  INV_X1 _53323_ (
    .A(_17696_),
    .ZN(_01454_)
  );
  AND2_X1 _53324_ (
    .A1(_12725_),
    .A2(_13304_),
    .ZN(_17697_)
  );
  INV_X1 _53325_ (
    .A(_17697_),
    .ZN(_17698_)
  );
  AND2_X1 _53326_ (
    .A1(\cpuregs[27] [29]),
    .A2(_12726_),
    .ZN(_17699_)
  );
  INV_X1 _53327_ (
    .A(_17699_),
    .ZN(_17700_)
  );
  AND2_X1 _53328_ (
    .A1(_17698_),
    .A2(_17700_),
    .ZN(_17701_)
  );
  INV_X1 _53329_ (
    .A(_17701_),
    .ZN(_01455_)
  );
  AND2_X1 _53330_ (
    .A1(_12725_),
    .A2(_13319_),
    .ZN(_17702_)
  );
  INV_X1 _53331_ (
    .A(_17702_),
    .ZN(_17703_)
  );
  AND2_X1 _53332_ (
    .A1(\cpuregs[27] [30]),
    .A2(_12726_),
    .ZN(_17704_)
  );
  INV_X1 _53333_ (
    .A(_17704_),
    .ZN(_17705_)
  );
  AND2_X1 _53334_ (
    .A1(_17703_),
    .A2(_17705_),
    .ZN(_17706_)
  );
  INV_X1 _53335_ (
    .A(_17706_),
    .ZN(_01456_)
  );
  AND2_X1 _53336_ (
    .A1(_12689_),
    .A2(_12874_),
    .ZN(_17707_)
  );
  INV_X1 _53337_ (
    .A(_17707_),
    .ZN(_17708_)
  );
  AND2_X1 _53338_ (
    .A1(\cpuregs[31] [0]),
    .A2(_12690_),
    .ZN(_17709_)
  );
  INV_X1 _53339_ (
    .A(_17709_),
    .ZN(_17710_)
  );
  AND2_X1 _53340_ (
    .A1(_17708_),
    .A2(_17710_),
    .ZN(_17711_)
  );
  INV_X1 _53341_ (
    .A(_17711_),
    .ZN(_01457_)
  );
  AND2_X1 _53342_ (
    .A1(_12689_),
    .A2(_12886_),
    .ZN(_17712_)
  );
  INV_X1 _53343_ (
    .A(_17712_),
    .ZN(_17713_)
  );
  AND2_X1 _53344_ (
    .A1(\cpuregs[31] [1]),
    .A2(_12690_),
    .ZN(_17714_)
  );
  INV_X1 _53345_ (
    .A(_17714_),
    .ZN(_17715_)
  );
  AND2_X1 _53346_ (
    .A1(_17713_),
    .A2(_17715_),
    .ZN(_17716_)
  );
  INV_X1 _53347_ (
    .A(_17716_),
    .ZN(_01458_)
  );
  AND2_X1 _53348_ (
    .A1(_12689_),
    .A2(_12900_),
    .ZN(_17717_)
  );
  INV_X1 _53349_ (
    .A(_17717_),
    .ZN(_17718_)
  );
  AND2_X1 _53350_ (
    .A1(\cpuregs[31] [2]),
    .A2(_12690_),
    .ZN(_17719_)
  );
  INV_X1 _53351_ (
    .A(_17719_),
    .ZN(_17720_)
  );
  AND2_X1 _53352_ (
    .A1(_17718_),
    .A2(_17720_),
    .ZN(_17721_)
  );
  INV_X1 _53353_ (
    .A(_17721_),
    .ZN(_01459_)
  );
  AND2_X1 _53354_ (
    .A1(_12689_),
    .A2(_12913_),
    .ZN(_17722_)
  );
  INV_X1 _53355_ (
    .A(_17722_),
    .ZN(_17723_)
  );
  AND2_X1 _53356_ (
    .A1(\cpuregs[31] [3]),
    .A2(_12690_),
    .ZN(_17724_)
  );
  INV_X1 _53357_ (
    .A(_17724_),
    .ZN(_17725_)
  );
  AND2_X1 _53358_ (
    .A1(_17723_),
    .A2(_17725_),
    .ZN(_17726_)
  );
  INV_X1 _53359_ (
    .A(_17726_),
    .ZN(_01460_)
  );
  AND2_X1 _53360_ (
    .A1(_12689_),
    .A2(_12928_),
    .ZN(_17727_)
  );
  INV_X1 _53361_ (
    .A(_17727_),
    .ZN(_17728_)
  );
  AND2_X1 _53362_ (
    .A1(\cpuregs[31] [4]),
    .A2(_12690_),
    .ZN(_17729_)
  );
  INV_X1 _53363_ (
    .A(_17729_),
    .ZN(_17730_)
  );
  AND2_X1 _53364_ (
    .A1(_17728_),
    .A2(_17730_),
    .ZN(_17731_)
  );
  INV_X1 _53365_ (
    .A(_17731_),
    .ZN(_01461_)
  );
  AND2_X1 _53366_ (
    .A1(_12689_),
    .A2(_12943_),
    .ZN(_17732_)
  );
  INV_X1 _53367_ (
    .A(_17732_),
    .ZN(_17733_)
  );
  AND2_X1 _53368_ (
    .A1(\cpuregs[31] [5]),
    .A2(_12690_),
    .ZN(_17734_)
  );
  INV_X1 _53369_ (
    .A(_17734_),
    .ZN(_17735_)
  );
  AND2_X1 _53370_ (
    .A1(_17733_),
    .A2(_17735_),
    .ZN(_17736_)
  );
  INV_X1 _53371_ (
    .A(_17736_),
    .ZN(_01462_)
  );
  AND2_X1 _53372_ (
    .A1(_12689_),
    .A2(_12958_),
    .ZN(_17737_)
  );
  INV_X1 _53373_ (
    .A(_17737_),
    .ZN(_17738_)
  );
  AND2_X1 _53374_ (
    .A1(\cpuregs[31] [6]),
    .A2(_12690_),
    .ZN(_17739_)
  );
  INV_X1 _53375_ (
    .A(_17739_),
    .ZN(_17740_)
  );
  AND2_X1 _53376_ (
    .A1(_17738_),
    .A2(_17740_),
    .ZN(_17741_)
  );
  INV_X1 _53377_ (
    .A(_17741_),
    .ZN(_01463_)
  );
  AND2_X1 _53378_ (
    .A1(_12689_),
    .A2(_12973_),
    .ZN(_17742_)
  );
  INV_X1 _53379_ (
    .A(_17742_),
    .ZN(_17743_)
  );
  AND2_X1 _53380_ (
    .A1(\cpuregs[31] [7]),
    .A2(_12690_),
    .ZN(_17744_)
  );
  INV_X1 _53381_ (
    .A(_17744_),
    .ZN(_17745_)
  );
  AND2_X1 _53382_ (
    .A1(_17743_),
    .A2(_17745_),
    .ZN(_17746_)
  );
  INV_X1 _53383_ (
    .A(_17746_),
    .ZN(_01464_)
  );
  AND2_X1 _53384_ (
    .A1(_12689_),
    .A2(_12988_),
    .ZN(_17747_)
  );
  INV_X1 _53385_ (
    .A(_17747_),
    .ZN(_17748_)
  );
  AND2_X1 _53386_ (
    .A1(\cpuregs[31] [8]),
    .A2(_12690_),
    .ZN(_17749_)
  );
  INV_X1 _53387_ (
    .A(_17749_),
    .ZN(_17750_)
  );
  AND2_X1 _53388_ (
    .A1(_17748_),
    .A2(_17750_),
    .ZN(_17751_)
  );
  INV_X1 _53389_ (
    .A(_17751_),
    .ZN(_01465_)
  );
  AND2_X1 _53390_ (
    .A1(_12689_),
    .A2(_13003_),
    .ZN(_17752_)
  );
  INV_X1 _53391_ (
    .A(_17752_),
    .ZN(_17753_)
  );
  AND2_X1 _53392_ (
    .A1(\cpuregs[31] [9]),
    .A2(_12690_),
    .ZN(_17754_)
  );
  INV_X1 _53393_ (
    .A(_17754_),
    .ZN(_17755_)
  );
  AND2_X1 _53394_ (
    .A1(_17753_),
    .A2(_17755_),
    .ZN(_17756_)
  );
  INV_X1 _53395_ (
    .A(_17756_),
    .ZN(_01466_)
  );
  AND2_X1 _53396_ (
    .A1(_12689_),
    .A2(_13018_),
    .ZN(_17757_)
  );
  INV_X1 _53397_ (
    .A(_17757_),
    .ZN(_17758_)
  );
  AND2_X1 _53398_ (
    .A1(\cpuregs[31] [10]),
    .A2(_12690_),
    .ZN(_17759_)
  );
  INV_X1 _53399_ (
    .A(_17759_),
    .ZN(_17760_)
  );
  AND2_X1 _53400_ (
    .A1(_17758_),
    .A2(_17760_),
    .ZN(_17761_)
  );
  INV_X1 _53401_ (
    .A(_17761_),
    .ZN(_01467_)
  );
  AND2_X1 _53402_ (
    .A1(_12689_),
    .A2(_13033_),
    .ZN(_17762_)
  );
  INV_X1 _53403_ (
    .A(_17762_),
    .ZN(_17763_)
  );
  AND2_X1 _53404_ (
    .A1(\cpuregs[31] [11]),
    .A2(_12690_),
    .ZN(_17764_)
  );
  INV_X1 _53405_ (
    .A(_17764_),
    .ZN(_17765_)
  );
  AND2_X1 _53406_ (
    .A1(_17763_),
    .A2(_17765_),
    .ZN(_17766_)
  );
  INV_X1 _53407_ (
    .A(_17766_),
    .ZN(_01468_)
  );
  AND2_X1 _53408_ (
    .A1(_12689_),
    .A2(_13048_),
    .ZN(_17767_)
  );
  INV_X1 _53409_ (
    .A(_17767_),
    .ZN(_17768_)
  );
  AND2_X1 _53410_ (
    .A1(\cpuregs[31] [12]),
    .A2(_12690_),
    .ZN(_17769_)
  );
  INV_X1 _53411_ (
    .A(_17769_),
    .ZN(_17770_)
  );
  AND2_X1 _53412_ (
    .A1(_17768_),
    .A2(_17770_),
    .ZN(_17771_)
  );
  INV_X1 _53413_ (
    .A(_17771_),
    .ZN(_01469_)
  );
  AND2_X1 _53414_ (
    .A1(_12689_),
    .A2(_13063_),
    .ZN(_17772_)
  );
  INV_X1 _53415_ (
    .A(_17772_),
    .ZN(_17773_)
  );
  AND2_X1 _53416_ (
    .A1(\cpuregs[31] [13]),
    .A2(_12690_),
    .ZN(_17774_)
  );
  INV_X1 _53417_ (
    .A(_17774_),
    .ZN(_17775_)
  );
  AND2_X1 _53418_ (
    .A1(_17773_),
    .A2(_17775_),
    .ZN(_17776_)
  );
  INV_X1 _53419_ (
    .A(_17776_),
    .ZN(_01470_)
  );
  AND2_X1 _53420_ (
    .A1(_12689_),
    .A2(_13078_),
    .ZN(_17777_)
  );
  INV_X1 _53421_ (
    .A(_17777_),
    .ZN(_17778_)
  );
  AND2_X1 _53422_ (
    .A1(\cpuregs[31] [14]),
    .A2(_12690_),
    .ZN(_17779_)
  );
  INV_X1 _53423_ (
    .A(_17779_),
    .ZN(_17780_)
  );
  AND2_X1 _53424_ (
    .A1(_17778_),
    .A2(_17780_),
    .ZN(_17781_)
  );
  INV_X1 _53425_ (
    .A(_17781_),
    .ZN(_01471_)
  );
  AND2_X1 _53426_ (
    .A1(_12689_),
    .A2(_13093_),
    .ZN(_17782_)
  );
  INV_X1 _53427_ (
    .A(_17782_),
    .ZN(_17783_)
  );
  AND2_X1 _53428_ (
    .A1(\cpuregs[31] [15]),
    .A2(_12690_),
    .ZN(_17784_)
  );
  INV_X1 _53429_ (
    .A(_17784_),
    .ZN(_17785_)
  );
  AND2_X1 _53430_ (
    .A1(_17783_),
    .A2(_17785_),
    .ZN(_17786_)
  );
  INV_X1 _53431_ (
    .A(_17786_),
    .ZN(_01472_)
  );
  AND2_X1 _53432_ (
    .A1(_12689_),
    .A2(_13108_),
    .ZN(_17787_)
  );
  INV_X1 _53433_ (
    .A(_17787_),
    .ZN(_17788_)
  );
  AND2_X1 _53434_ (
    .A1(\cpuregs[31] [16]),
    .A2(_12690_),
    .ZN(_17789_)
  );
  INV_X1 _53435_ (
    .A(_17789_),
    .ZN(_17790_)
  );
  AND2_X1 _53436_ (
    .A1(_17788_),
    .A2(_17790_),
    .ZN(_17791_)
  );
  INV_X1 _53437_ (
    .A(_17791_),
    .ZN(_01473_)
  );
  AND2_X1 _53438_ (
    .A1(_12689_),
    .A2(_13123_),
    .ZN(_17792_)
  );
  INV_X1 _53439_ (
    .A(_17792_),
    .ZN(_17793_)
  );
  AND2_X1 _53440_ (
    .A1(\cpuregs[31] [17]),
    .A2(_12690_),
    .ZN(_17794_)
  );
  INV_X1 _53441_ (
    .A(_17794_),
    .ZN(_17795_)
  );
  AND2_X1 _53442_ (
    .A1(_17793_),
    .A2(_17795_),
    .ZN(_17796_)
  );
  INV_X1 _53443_ (
    .A(_17796_),
    .ZN(_01474_)
  );
  AND2_X1 _53444_ (
    .A1(_12689_),
    .A2(_13139_),
    .ZN(_17797_)
  );
  INV_X1 _53445_ (
    .A(_17797_),
    .ZN(_17798_)
  );
  AND2_X1 _53446_ (
    .A1(\cpuregs[31] [18]),
    .A2(_12690_),
    .ZN(_17799_)
  );
  INV_X1 _53447_ (
    .A(_17799_),
    .ZN(_17800_)
  );
  AND2_X1 _53448_ (
    .A1(_17798_),
    .A2(_17800_),
    .ZN(_17801_)
  );
  INV_X1 _53449_ (
    .A(_17801_),
    .ZN(_01475_)
  );
  AND2_X1 _53450_ (
    .A1(_12689_),
    .A2(_13154_),
    .ZN(_17802_)
  );
  INV_X1 _53451_ (
    .A(_17802_),
    .ZN(_17803_)
  );
  AND2_X1 _53452_ (
    .A1(\cpuregs[31] [19]),
    .A2(_12690_),
    .ZN(_17804_)
  );
  INV_X1 _53453_ (
    .A(_17804_),
    .ZN(_17805_)
  );
  AND2_X1 _53454_ (
    .A1(_17803_),
    .A2(_17805_),
    .ZN(_17806_)
  );
  INV_X1 _53455_ (
    .A(_17806_),
    .ZN(_01476_)
  );
  AND2_X1 _53456_ (
    .A1(_12689_),
    .A2(_13169_),
    .ZN(_17807_)
  );
  INV_X1 _53457_ (
    .A(_17807_),
    .ZN(_17808_)
  );
  AND2_X1 _53458_ (
    .A1(\cpuregs[31] [20]),
    .A2(_12690_),
    .ZN(_17809_)
  );
  INV_X1 _53459_ (
    .A(_17809_),
    .ZN(_17810_)
  );
  AND2_X1 _53460_ (
    .A1(_17808_),
    .A2(_17810_),
    .ZN(_17811_)
  );
  INV_X1 _53461_ (
    .A(_17811_),
    .ZN(_01477_)
  );
  AND2_X1 _53462_ (
    .A1(_12689_),
    .A2(_13184_),
    .ZN(_17812_)
  );
  INV_X1 _53463_ (
    .A(_17812_),
    .ZN(_17813_)
  );
  AND2_X1 _53464_ (
    .A1(\cpuregs[31] [21]),
    .A2(_12690_),
    .ZN(_17814_)
  );
  INV_X1 _53465_ (
    .A(_17814_),
    .ZN(_17815_)
  );
  AND2_X1 _53466_ (
    .A1(_17813_),
    .A2(_17815_),
    .ZN(_17816_)
  );
  INV_X1 _53467_ (
    .A(_17816_),
    .ZN(_01478_)
  );
  AND2_X1 _53468_ (
    .A1(_12689_),
    .A2(_13199_),
    .ZN(_17817_)
  );
  INV_X1 _53469_ (
    .A(_17817_),
    .ZN(_17818_)
  );
  AND2_X1 _53470_ (
    .A1(\cpuregs[31] [22]),
    .A2(_12690_),
    .ZN(_17819_)
  );
  INV_X1 _53471_ (
    .A(_17819_),
    .ZN(_17820_)
  );
  AND2_X1 _53472_ (
    .A1(_17818_),
    .A2(_17820_),
    .ZN(_17821_)
  );
  INV_X1 _53473_ (
    .A(_17821_),
    .ZN(_01479_)
  );
  AND2_X1 _53474_ (
    .A1(_12689_),
    .A2(_13214_),
    .ZN(_17822_)
  );
  INV_X1 _53475_ (
    .A(_17822_),
    .ZN(_17823_)
  );
  AND2_X1 _53476_ (
    .A1(\cpuregs[31] [23]),
    .A2(_12690_),
    .ZN(_17824_)
  );
  INV_X1 _53477_ (
    .A(_17824_),
    .ZN(_17825_)
  );
  AND2_X1 _53478_ (
    .A1(_17823_),
    .A2(_17825_),
    .ZN(_17826_)
  );
  INV_X1 _53479_ (
    .A(_17826_),
    .ZN(_01480_)
  );
  AND2_X1 _53480_ (
    .A1(_12689_),
    .A2(_13229_),
    .ZN(_17827_)
  );
  INV_X1 _53481_ (
    .A(_17827_),
    .ZN(_17828_)
  );
  AND2_X1 _53482_ (
    .A1(\cpuregs[31] [24]),
    .A2(_12690_),
    .ZN(_17829_)
  );
  INV_X1 _53483_ (
    .A(_17829_),
    .ZN(_17830_)
  );
  AND2_X1 _53484_ (
    .A1(_17828_),
    .A2(_17830_),
    .ZN(_17831_)
  );
  INV_X1 _53485_ (
    .A(_17831_),
    .ZN(_01481_)
  );
  AND2_X1 _53486_ (
    .A1(_12689_),
    .A2(_13244_),
    .ZN(_17832_)
  );
  INV_X1 _53487_ (
    .A(_17832_),
    .ZN(_17833_)
  );
  AND2_X1 _53488_ (
    .A1(\cpuregs[31] [25]),
    .A2(_12690_),
    .ZN(_17834_)
  );
  INV_X1 _53489_ (
    .A(_17834_),
    .ZN(_17835_)
  );
  AND2_X1 _53490_ (
    .A1(_17833_),
    .A2(_17835_),
    .ZN(_17836_)
  );
  INV_X1 _53491_ (
    .A(_17836_),
    .ZN(_01482_)
  );
  AND2_X1 _53492_ (
    .A1(_12689_),
    .A2(_13259_),
    .ZN(_17837_)
  );
  INV_X1 _53493_ (
    .A(_17837_),
    .ZN(_17838_)
  );
  AND2_X1 _53494_ (
    .A1(\cpuregs[31] [26]),
    .A2(_12690_),
    .ZN(_17839_)
  );
  INV_X1 _53495_ (
    .A(_17839_),
    .ZN(_17840_)
  );
  AND2_X1 _53496_ (
    .A1(_17838_),
    .A2(_17840_),
    .ZN(_17841_)
  );
  INV_X1 _53497_ (
    .A(_17841_),
    .ZN(_01483_)
  );
  AND2_X1 _53498_ (
    .A1(_12689_),
    .A2(_13274_),
    .ZN(_17842_)
  );
  INV_X1 _53499_ (
    .A(_17842_),
    .ZN(_17843_)
  );
  AND2_X1 _53500_ (
    .A1(\cpuregs[31] [27]),
    .A2(_12690_),
    .ZN(_17844_)
  );
  INV_X1 _53501_ (
    .A(_17844_),
    .ZN(_17845_)
  );
  AND2_X1 _53502_ (
    .A1(_17843_),
    .A2(_17845_),
    .ZN(_17846_)
  );
  INV_X1 _53503_ (
    .A(_17846_),
    .ZN(_01484_)
  );
  AND2_X1 _53504_ (
    .A1(_12689_),
    .A2(_13289_),
    .ZN(_17847_)
  );
  INV_X1 _53505_ (
    .A(_17847_),
    .ZN(_17848_)
  );
  AND2_X1 _53506_ (
    .A1(\cpuregs[31] [28]),
    .A2(_12690_),
    .ZN(_17849_)
  );
  INV_X1 _53507_ (
    .A(_17849_),
    .ZN(_17850_)
  );
  AND2_X1 _53508_ (
    .A1(_17848_),
    .A2(_17850_),
    .ZN(_17851_)
  );
  INV_X1 _53509_ (
    .A(_17851_),
    .ZN(_01485_)
  );
  AND2_X1 _53510_ (
    .A1(_12689_),
    .A2(_13304_),
    .ZN(_17852_)
  );
  INV_X1 _53511_ (
    .A(_17852_),
    .ZN(_17853_)
  );
  AND2_X1 _53512_ (
    .A1(\cpuregs[31] [29]),
    .A2(_12690_),
    .ZN(_17854_)
  );
  INV_X1 _53513_ (
    .A(_17854_),
    .ZN(_17855_)
  );
  AND2_X1 _53514_ (
    .A1(_17853_),
    .A2(_17855_),
    .ZN(_17856_)
  );
  INV_X1 _53515_ (
    .A(_17856_),
    .ZN(_01486_)
  );
  AND2_X1 _53516_ (
    .A1(_12689_),
    .A2(_13319_),
    .ZN(_17857_)
  );
  INV_X1 _53517_ (
    .A(_17857_),
    .ZN(_17858_)
  );
  AND2_X1 _53518_ (
    .A1(\cpuregs[31] [30]),
    .A2(_12690_),
    .ZN(_17859_)
  );
  INV_X1 _53519_ (
    .A(_17859_),
    .ZN(_17860_)
  );
  AND2_X1 _53520_ (
    .A1(_17858_),
    .A2(_17860_),
    .ZN(_17861_)
  );
  INV_X1 _53521_ (
    .A(_17861_),
    .ZN(_01487_)
  );
  AND2_X1 _53522_ (
    .A1(_21978_),
    .A2(_02901_),
    .ZN(_17862_)
  );
  INV_X1 _53523_ (
    .A(_17862_),
    .ZN(_17863_)
  );
  AND2_X1 _53524_ (
    .A1(mem_rdata_q[31]),
    .A2(_22523_),
    .ZN(_17864_)
  );
  INV_X1 _53525_ (
    .A(_17864_),
    .ZN(_17865_)
  );
  AND2_X1 _53526_ (
    .A1(mem_rdata_q[31]),
    .A2(_11684_),
    .ZN(_17866_)
  );
  INV_X1 _53527_ (
    .A(_17866_),
    .ZN(_17867_)
  );
  AND2_X1 _53528_ (
    .A1(_02900_),
    .A2(_17867_),
    .ZN(_17868_)
  );
  AND2_X1 _53529_ (
    .A1(instr_jal),
    .A2(decoded_imm_j[30]),
    .ZN(_17869_)
  );
  INV_X1 _53530_ (
    .A(_17869_),
    .ZN(_17870_)
  );
  AND2_X1 _53531_ (
    .A1(_21039_),
    .A2(_21290_),
    .ZN(_17871_)
  );
  INV_X1 _53532_ (
    .A(_17871_),
    .ZN(_17872_)
  );
  AND2_X1 _53533_ (
    .A1(mem_rdata_q[31]),
    .A2(_17872_),
    .ZN(_17873_)
  );
  INV_X1 _53534_ (
    .A(_17873_),
    .ZN(_17874_)
  );
  AND2_X1 _53535_ (
    .A1(_17870_),
    .A2(_17874_),
    .ZN(_17875_)
  );
  AND2_X1 _53536_ (
    .A1(_17868_),
    .A2(_17875_),
    .ZN(_17876_)
  );
  AND2_X1 _53537_ (
    .A1(_17865_),
    .A2(_17876_),
    .ZN(_17877_)
  );
  INV_X1 _53538_ (
    .A(_17877_),
    .ZN(_17878_)
  );
  AND2_X1 _53539_ (
    .A1(_17863_),
    .A2(_17878_),
    .ZN(_01519_)
  );
  AND2_X1 _53540_ (
    .A1(_21979_),
    .A2(_02901_),
    .ZN(_17879_)
  );
  INV_X1 _53541_ (
    .A(_17879_),
    .ZN(_17880_)
  );
  AND2_X1 _53542_ (
    .A1(mem_rdata_q[30]),
    .A2(_22523_),
    .ZN(_17881_)
  );
  INV_X1 _53543_ (
    .A(_17881_),
    .ZN(_17882_)
  );
  AND2_X1 _53544_ (
    .A1(_17876_),
    .A2(_17882_),
    .ZN(_17883_)
  );
  INV_X1 _53545_ (
    .A(_17883_),
    .ZN(_17884_)
  );
  AND2_X1 _53546_ (
    .A1(_17880_),
    .A2(_17884_),
    .ZN(_01520_)
  );
  AND2_X1 _53547_ (
    .A1(_21980_),
    .A2(_02901_),
    .ZN(_17885_)
  );
  INV_X1 _53548_ (
    .A(_17885_),
    .ZN(_17886_)
  );
  AND2_X1 _53549_ (
    .A1(mem_rdata_q[29]),
    .A2(_22523_),
    .ZN(_17887_)
  );
  INV_X1 _53550_ (
    .A(_17887_),
    .ZN(_17888_)
  );
  AND2_X1 _53551_ (
    .A1(_17876_),
    .A2(_17888_),
    .ZN(_17889_)
  );
  INV_X1 _53552_ (
    .A(_17889_),
    .ZN(_17890_)
  );
  AND2_X1 _53553_ (
    .A1(_17886_),
    .A2(_17890_),
    .ZN(_01521_)
  );
  AND2_X1 _53554_ (
    .A1(_21981_),
    .A2(_02901_),
    .ZN(_17891_)
  );
  INV_X1 _53555_ (
    .A(_17891_),
    .ZN(_17892_)
  );
  AND2_X1 _53556_ (
    .A1(mem_rdata_q[28]),
    .A2(_22523_),
    .ZN(_17893_)
  );
  INV_X1 _53557_ (
    .A(_17893_),
    .ZN(_17894_)
  );
  AND2_X1 _53558_ (
    .A1(_17876_),
    .A2(_17894_),
    .ZN(_17895_)
  );
  INV_X1 _53559_ (
    .A(_17895_),
    .ZN(_17896_)
  );
  AND2_X1 _53560_ (
    .A1(_17892_),
    .A2(_17896_),
    .ZN(_01522_)
  );
  AND2_X1 _53561_ (
    .A1(_21982_),
    .A2(_02901_),
    .ZN(_17897_)
  );
  INV_X1 _53562_ (
    .A(_17897_),
    .ZN(_17898_)
  );
  AND2_X1 _53563_ (
    .A1(mem_rdata_q[27]),
    .A2(_22523_),
    .ZN(_17899_)
  );
  INV_X1 _53564_ (
    .A(_17899_),
    .ZN(_17900_)
  );
  AND2_X1 _53565_ (
    .A1(_17876_),
    .A2(_17900_),
    .ZN(_17901_)
  );
  INV_X1 _53566_ (
    .A(_17901_),
    .ZN(_17902_)
  );
  AND2_X1 _53567_ (
    .A1(_17898_),
    .A2(_17902_),
    .ZN(_01523_)
  );
  AND2_X1 _53568_ (
    .A1(_21983_),
    .A2(_02901_),
    .ZN(_17903_)
  );
  INV_X1 _53569_ (
    .A(_17903_),
    .ZN(_17904_)
  );
  AND2_X1 _53570_ (
    .A1(mem_rdata_q[26]),
    .A2(_22523_),
    .ZN(_17905_)
  );
  INV_X1 _53571_ (
    .A(_17905_),
    .ZN(_17906_)
  );
  AND2_X1 _53572_ (
    .A1(_17876_),
    .A2(_17906_),
    .ZN(_17907_)
  );
  INV_X1 _53573_ (
    .A(_17907_),
    .ZN(_17908_)
  );
  AND2_X1 _53574_ (
    .A1(_17904_),
    .A2(_17908_),
    .ZN(_01524_)
  );
  AND2_X1 _53575_ (
    .A1(_21984_),
    .A2(_02901_),
    .ZN(_17909_)
  );
  INV_X1 _53576_ (
    .A(_17909_),
    .ZN(_17910_)
  );
  AND2_X1 _53577_ (
    .A1(mem_rdata_q[25]),
    .A2(_22523_),
    .ZN(_17911_)
  );
  INV_X1 _53578_ (
    .A(_17911_),
    .ZN(_17912_)
  );
  AND2_X1 _53579_ (
    .A1(_17876_),
    .A2(_17912_),
    .ZN(_17913_)
  );
  INV_X1 _53580_ (
    .A(_17913_),
    .ZN(_17914_)
  );
  AND2_X1 _53581_ (
    .A1(_17910_),
    .A2(_17914_),
    .ZN(_01525_)
  );
  AND2_X1 _53582_ (
    .A1(_21985_),
    .A2(_02901_),
    .ZN(_17915_)
  );
  INV_X1 _53583_ (
    .A(_17915_),
    .ZN(_17916_)
  );
  AND2_X1 _53584_ (
    .A1(mem_rdata_q[24]),
    .A2(_22523_),
    .ZN(_17917_)
  );
  INV_X1 _53585_ (
    .A(_17917_),
    .ZN(_17918_)
  );
  AND2_X1 _53586_ (
    .A1(_17876_),
    .A2(_17918_),
    .ZN(_17919_)
  );
  INV_X1 _53587_ (
    .A(_17919_),
    .ZN(_17920_)
  );
  AND2_X1 _53588_ (
    .A1(_17916_),
    .A2(_17920_),
    .ZN(_01526_)
  );
  AND2_X1 _53589_ (
    .A1(_21986_),
    .A2(_02901_),
    .ZN(_17921_)
  );
  INV_X1 _53590_ (
    .A(_17921_),
    .ZN(_17922_)
  );
  AND2_X1 _53591_ (
    .A1(mem_rdata_q[23]),
    .A2(_22523_),
    .ZN(_17923_)
  );
  INV_X1 _53592_ (
    .A(_17923_),
    .ZN(_17924_)
  );
  AND2_X1 _53593_ (
    .A1(_17876_),
    .A2(_17924_),
    .ZN(_17925_)
  );
  INV_X1 _53594_ (
    .A(_17925_),
    .ZN(_17926_)
  );
  AND2_X1 _53595_ (
    .A1(_17922_),
    .A2(_17926_),
    .ZN(_01527_)
  );
  AND2_X1 _53596_ (
    .A1(_21987_),
    .A2(_02901_),
    .ZN(_17927_)
  );
  INV_X1 _53597_ (
    .A(_17927_),
    .ZN(_17928_)
  );
  AND2_X1 _53598_ (
    .A1(mem_rdata_q[22]),
    .A2(_22523_),
    .ZN(_17929_)
  );
  INV_X1 _53599_ (
    .A(_17929_),
    .ZN(_17930_)
  );
  AND2_X1 _53600_ (
    .A1(_17876_),
    .A2(_17930_),
    .ZN(_17931_)
  );
  INV_X1 _53601_ (
    .A(_17931_),
    .ZN(_17932_)
  );
  AND2_X1 _53602_ (
    .A1(_17928_),
    .A2(_17932_),
    .ZN(_01528_)
  );
  AND2_X1 _53603_ (
    .A1(_21988_),
    .A2(_02901_),
    .ZN(_17933_)
  );
  INV_X1 _53604_ (
    .A(_17933_),
    .ZN(_17934_)
  );
  AND2_X1 _53605_ (
    .A1(mem_rdata_q[21]),
    .A2(_22523_),
    .ZN(_17935_)
  );
  INV_X1 _53606_ (
    .A(_17935_),
    .ZN(_17936_)
  );
  AND2_X1 _53607_ (
    .A1(_17876_),
    .A2(_17936_),
    .ZN(_17937_)
  );
  INV_X1 _53608_ (
    .A(_17937_),
    .ZN(_17938_)
  );
  AND2_X1 _53609_ (
    .A1(_17934_),
    .A2(_17938_),
    .ZN(_01529_)
  );
  AND2_X1 _53610_ (
    .A1(_21989_),
    .A2(_02901_),
    .ZN(_17939_)
  );
  INV_X1 _53611_ (
    .A(_17939_),
    .ZN(_17940_)
  );
  AND2_X1 _53612_ (
    .A1(mem_rdata_q[20]),
    .A2(_22523_),
    .ZN(_17941_)
  );
  INV_X1 _53613_ (
    .A(_17941_),
    .ZN(_17942_)
  );
  AND2_X1 _53614_ (
    .A1(_17876_),
    .A2(_17942_),
    .ZN(_17943_)
  );
  INV_X1 _53615_ (
    .A(_17943_),
    .ZN(_17944_)
  );
  AND2_X1 _53616_ (
    .A1(_17940_),
    .A2(_17944_),
    .ZN(_01530_)
  );
  AND2_X1 _53617_ (
    .A1(_21990_),
    .A2(_02901_),
    .ZN(_17945_)
  );
  INV_X1 _53618_ (
    .A(_17945_),
    .ZN(_17946_)
  );
  AND2_X1 _53619_ (
    .A1(_17868_),
    .A2(_17874_),
    .ZN(_17947_)
  );
  AND2_X1 _53620_ (
    .A1(mem_rdata_q[19]),
    .A2(_22523_),
    .ZN(_17948_)
  );
  INV_X1 _53621_ (
    .A(_17948_),
    .ZN(_17949_)
  );
  AND2_X1 _53622_ (
    .A1(instr_jal),
    .A2(decoded_imm_j[19]),
    .ZN(_17950_)
  );
  INV_X1 _53623_ (
    .A(_17950_),
    .ZN(_17951_)
  );
  AND2_X1 _53624_ (
    .A1(_17949_),
    .A2(_17951_),
    .ZN(_17952_)
  );
  AND2_X1 _53625_ (
    .A1(_17947_),
    .A2(_17952_),
    .ZN(_17953_)
  );
  INV_X1 _53626_ (
    .A(_17953_),
    .ZN(_17954_)
  );
  AND2_X1 _53627_ (
    .A1(_17946_),
    .A2(_17954_),
    .ZN(_01531_)
  );
  AND2_X1 _53628_ (
    .A1(_21991_),
    .A2(_02901_),
    .ZN(_17955_)
  );
  INV_X1 _53629_ (
    .A(_17955_),
    .ZN(_17956_)
  );
  AND2_X1 _53630_ (
    .A1(mem_rdata_q[18]),
    .A2(_22523_),
    .ZN(_17957_)
  );
  INV_X1 _53631_ (
    .A(_17957_),
    .ZN(_17958_)
  );
  AND2_X1 _53632_ (
    .A1(instr_jal),
    .A2(decoded_imm_j[18]),
    .ZN(_17959_)
  );
  INV_X1 _53633_ (
    .A(_17959_),
    .ZN(_17960_)
  );
  AND2_X1 _53634_ (
    .A1(_17958_),
    .A2(_17960_),
    .ZN(_17961_)
  );
  AND2_X1 _53635_ (
    .A1(_17947_),
    .A2(_17961_),
    .ZN(_17962_)
  );
  INV_X1 _53636_ (
    .A(_17962_),
    .ZN(_17963_)
  );
  AND2_X1 _53637_ (
    .A1(_17956_),
    .A2(_17963_),
    .ZN(_01532_)
  );
  AND2_X1 _53638_ (
    .A1(_21992_),
    .A2(_02901_),
    .ZN(_17964_)
  );
  INV_X1 _53639_ (
    .A(_17964_),
    .ZN(_17965_)
  );
  AND2_X1 _53640_ (
    .A1(instr_jal),
    .A2(decoded_rs1[2]),
    .ZN(_17966_)
  );
  INV_X1 _53641_ (
    .A(_17966_),
    .ZN(_17967_)
  );
  AND2_X1 _53642_ (
    .A1(mem_rdata_q[17]),
    .A2(_22523_),
    .ZN(_17968_)
  );
  INV_X1 _53643_ (
    .A(_17968_),
    .ZN(_17969_)
  );
  AND2_X1 _53644_ (
    .A1(_17967_),
    .A2(_17969_),
    .ZN(_17970_)
  );
  AND2_X1 _53645_ (
    .A1(_17947_),
    .A2(_17970_),
    .ZN(_17971_)
  );
  INV_X1 _53646_ (
    .A(_17971_),
    .ZN(_17972_)
  );
  AND2_X1 _53647_ (
    .A1(_17965_),
    .A2(_17972_),
    .ZN(_01533_)
  );
  AND2_X1 _53648_ (
    .A1(_21993_),
    .A2(_02901_),
    .ZN(_17973_)
  );
  INV_X1 _53649_ (
    .A(_17973_),
    .ZN(_17974_)
  );
  AND2_X1 _53650_ (
    .A1(mem_rdata_q[16]),
    .A2(_22523_),
    .ZN(_17975_)
  );
  INV_X1 _53651_ (
    .A(_17975_),
    .ZN(_17976_)
  );
  AND2_X1 _53652_ (
    .A1(instr_jal),
    .A2(decoded_rs1[1]),
    .ZN(_17977_)
  );
  INV_X1 _53653_ (
    .A(_17977_),
    .ZN(_17978_)
  );
  AND2_X1 _53654_ (
    .A1(_17976_),
    .A2(_17978_),
    .ZN(_17979_)
  );
  AND2_X1 _53655_ (
    .A1(_17947_),
    .A2(_17979_),
    .ZN(_17980_)
  );
  INV_X1 _53656_ (
    .A(_17980_),
    .ZN(_17981_)
  );
  AND2_X1 _53657_ (
    .A1(_17974_),
    .A2(_17981_),
    .ZN(_01534_)
  );
  AND2_X1 _53658_ (
    .A1(_21994_),
    .A2(_02901_),
    .ZN(_17982_)
  );
  INV_X1 _53659_ (
    .A(_17982_),
    .ZN(_17983_)
  );
  AND2_X1 _53660_ (
    .A1(mem_rdata_q[15]),
    .A2(_22523_),
    .ZN(_17984_)
  );
  INV_X1 _53661_ (
    .A(_17984_),
    .ZN(_17985_)
  );
  AND2_X1 _53662_ (
    .A1(instr_jal),
    .A2(decoded_rs1[0]),
    .ZN(_17986_)
  );
  INV_X1 _53663_ (
    .A(_17986_),
    .ZN(_17987_)
  );
  AND2_X1 _53664_ (
    .A1(_17985_),
    .A2(_17987_),
    .ZN(_17988_)
  );
  AND2_X1 _53665_ (
    .A1(_17947_),
    .A2(_17988_),
    .ZN(_17989_)
  );
  INV_X1 _53666_ (
    .A(_17989_),
    .ZN(_17990_)
  );
  AND2_X1 _53667_ (
    .A1(_17983_),
    .A2(_17990_),
    .ZN(_01535_)
  );
  AND2_X1 _53668_ (
    .A1(_21995_),
    .A2(_02901_),
    .ZN(_17991_)
  );
  INV_X1 _53669_ (
    .A(_17991_),
    .ZN(_17992_)
  );
  AND2_X1 _53670_ (
    .A1(mem_rdata_q[14]),
    .A2(_22523_),
    .ZN(_17993_)
  );
  INV_X1 _53671_ (
    .A(_17993_),
    .ZN(_17994_)
  );
  AND2_X1 _53672_ (
    .A1(instr_jal),
    .A2(decoded_imm_j[14]),
    .ZN(_17995_)
  );
  INV_X1 _53673_ (
    .A(_17995_),
    .ZN(_17996_)
  );
  AND2_X1 _53674_ (
    .A1(_17994_),
    .A2(_17996_),
    .ZN(_17997_)
  );
  AND2_X1 _53675_ (
    .A1(_17947_),
    .A2(_17997_),
    .ZN(_17998_)
  );
  INV_X1 _53676_ (
    .A(_17998_),
    .ZN(_17999_)
  );
  AND2_X1 _53677_ (
    .A1(_17992_),
    .A2(_17999_),
    .ZN(_01536_)
  );
  AND2_X1 _53678_ (
    .A1(_21996_),
    .A2(_02901_),
    .ZN(_18000_)
  );
  INV_X1 _53679_ (
    .A(_18000_),
    .ZN(_18001_)
  );
  AND2_X1 _53680_ (
    .A1(mem_rdata_q[13]),
    .A2(_22523_),
    .ZN(_18002_)
  );
  INV_X1 _53681_ (
    .A(_18002_),
    .ZN(_18003_)
  );
  AND2_X1 _53682_ (
    .A1(instr_jal),
    .A2(decoded_imm_j[13]),
    .ZN(_18004_)
  );
  INV_X1 _53683_ (
    .A(_18004_),
    .ZN(_18005_)
  );
  AND2_X1 _53684_ (
    .A1(_18003_),
    .A2(_18005_),
    .ZN(_18006_)
  );
  AND2_X1 _53685_ (
    .A1(_17947_),
    .A2(_18006_),
    .ZN(_18007_)
  );
  INV_X1 _53686_ (
    .A(_18007_),
    .ZN(_18008_)
  );
  AND2_X1 _53687_ (
    .A1(_18001_),
    .A2(_18008_),
    .ZN(_01537_)
  );
  AND2_X1 _53688_ (
    .A1(_21997_),
    .A2(_02901_),
    .ZN(_18009_)
  );
  INV_X1 _53689_ (
    .A(_18009_),
    .ZN(_18010_)
  );
  AND2_X1 _53690_ (
    .A1(mem_rdata_q[12]),
    .A2(_22523_),
    .ZN(_18011_)
  );
  INV_X1 _53691_ (
    .A(_18011_),
    .ZN(_18012_)
  );
  AND2_X1 _53692_ (
    .A1(instr_jal),
    .A2(decoded_imm_j[12]),
    .ZN(_18013_)
  );
  INV_X1 _53693_ (
    .A(_18013_),
    .ZN(_18014_)
  );
  AND2_X1 _53694_ (
    .A1(_18012_),
    .A2(_18014_),
    .ZN(_18015_)
  );
  AND2_X1 _53695_ (
    .A1(_17947_),
    .A2(_18015_),
    .ZN(_18016_)
  );
  INV_X1 _53696_ (
    .A(_18016_),
    .ZN(_18017_)
  );
  AND2_X1 _53697_ (
    .A1(_18010_),
    .A2(_18017_),
    .ZN(_01538_)
  );
  AND2_X1 _53698_ (
    .A1(_21998_),
    .A2(_02901_),
    .ZN(_18018_)
  );
  INV_X1 _53699_ (
    .A(_18018_),
    .ZN(_18019_)
  );
  AND2_X1 _53700_ (
    .A1(is_beq_bne_blt_bge_bltu_bgeu),
    .A2(mem_rdata_q[7]),
    .ZN(_18020_)
  );
  INV_X1 _53701_ (
    .A(_18020_),
    .ZN(_18021_)
  );
  AND2_X1 _53702_ (
    .A1(mem_rdata_q[31]),
    .A2(is_sb_sh_sw),
    .ZN(_18022_)
  );
  INV_X1 _53703_ (
    .A(_18022_),
    .ZN(_18023_)
  );
  AND2_X1 _53704_ (
    .A1(instr_jal),
    .A2(decoded_rs2[0]),
    .ZN(_18024_)
  );
  INV_X1 _53705_ (
    .A(_18024_),
    .ZN(_18025_)
  );
  AND2_X1 _53706_ (
    .A1(_18023_),
    .A2(_18025_),
    .ZN(_18026_)
  );
  AND2_X1 _53707_ (
    .A1(_18021_),
    .A2(_18026_),
    .ZN(_18027_)
  );
  AND2_X1 _53708_ (
    .A1(_17868_),
    .A2(_18027_),
    .ZN(_18028_)
  );
  INV_X1 _53709_ (
    .A(_18028_),
    .ZN(_18029_)
  );
  AND2_X1 _53710_ (
    .A1(_18019_),
    .A2(_18029_),
    .ZN(_01539_)
  );
  AND2_X1 _53711_ (
    .A1(_11683_),
    .A2(_17871_),
    .ZN(_18030_)
  );
  INV_X1 _53712_ (
    .A(_18030_),
    .ZN(_18031_)
  );
  AND2_X1 _53713_ (
    .A1(mem_rdata_q[30]),
    .A2(_18031_),
    .ZN(_18032_)
  );
  INV_X1 _53714_ (
    .A(_18032_),
    .ZN(_18033_)
  );
  AND2_X1 _53715_ (
    .A1(instr_jal),
    .A2(decoded_imm_j[10]),
    .ZN(_18034_)
  );
  INV_X1 _53716_ (
    .A(_18034_),
    .ZN(_18035_)
  );
  AND2_X1 _53717_ (
    .A1(_21999_),
    .A2(_02901_),
    .ZN(_18036_)
  );
  INV_X1 _53718_ (
    .A(_18036_),
    .ZN(_18037_)
  );
  AND2_X1 _53719_ (
    .A1(_02900_),
    .A2(_18035_),
    .ZN(_18038_)
  );
  AND2_X1 _53720_ (
    .A1(_18033_),
    .A2(_18038_),
    .ZN(_18039_)
  );
  INV_X1 _53721_ (
    .A(_18039_),
    .ZN(_18040_)
  );
  AND2_X1 _53722_ (
    .A1(_18037_),
    .A2(_18040_),
    .ZN(_01540_)
  );
  AND2_X1 _53723_ (
    .A1(mem_rdata_q[29]),
    .A2(_18031_),
    .ZN(_18041_)
  );
  INV_X1 _53724_ (
    .A(_18041_),
    .ZN(_18042_)
  );
  AND2_X1 _53725_ (
    .A1(instr_jal),
    .A2(decoded_imm_j[9]),
    .ZN(_18043_)
  );
  INV_X1 _53726_ (
    .A(_18043_),
    .ZN(_18044_)
  );
  AND2_X1 _53727_ (
    .A1(_22000_),
    .A2(_02901_),
    .ZN(_18045_)
  );
  INV_X1 _53728_ (
    .A(_18045_),
    .ZN(_18046_)
  );
  AND2_X1 _53729_ (
    .A1(_02900_),
    .A2(_18044_),
    .ZN(_18047_)
  );
  AND2_X1 _53730_ (
    .A1(_18042_),
    .A2(_18047_),
    .ZN(_18048_)
  );
  INV_X1 _53731_ (
    .A(_18048_),
    .ZN(_18049_)
  );
  AND2_X1 _53732_ (
    .A1(_18046_),
    .A2(_18049_),
    .ZN(_01541_)
  );
  AND2_X1 _53733_ (
    .A1(mem_rdata_q[28]),
    .A2(_18031_),
    .ZN(_18050_)
  );
  INV_X1 _53734_ (
    .A(_18050_),
    .ZN(_18051_)
  );
  AND2_X1 _53735_ (
    .A1(instr_jal),
    .A2(decoded_imm_j[8]),
    .ZN(_18052_)
  );
  INV_X1 _53736_ (
    .A(_18052_),
    .ZN(_18053_)
  );
  AND2_X1 _53737_ (
    .A1(_22001_),
    .A2(_02901_),
    .ZN(_18054_)
  );
  INV_X1 _53738_ (
    .A(_18054_),
    .ZN(_18055_)
  );
  AND2_X1 _53739_ (
    .A1(_02900_),
    .A2(_18053_),
    .ZN(_18056_)
  );
  AND2_X1 _53740_ (
    .A1(_18051_),
    .A2(_18056_),
    .ZN(_18057_)
  );
  INV_X1 _53741_ (
    .A(_18057_),
    .ZN(_18058_)
  );
  AND2_X1 _53742_ (
    .A1(_18055_),
    .A2(_18058_),
    .ZN(_01542_)
  );
  AND2_X1 _53743_ (
    .A1(mem_rdata_q[27]),
    .A2(_18031_),
    .ZN(_18059_)
  );
  INV_X1 _53744_ (
    .A(_18059_),
    .ZN(_18060_)
  );
  AND2_X1 _53745_ (
    .A1(instr_jal),
    .A2(decoded_imm_j[7]),
    .ZN(_18061_)
  );
  INV_X1 _53746_ (
    .A(_18061_),
    .ZN(_18062_)
  );
  AND2_X1 _53747_ (
    .A1(_22002_),
    .A2(_02901_),
    .ZN(_18063_)
  );
  INV_X1 _53748_ (
    .A(_18063_),
    .ZN(_18064_)
  );
  AND2_X1 _53749_ (
    .A1(_02900_),
    .A2(_18062_),
    .ZN(_18065_)
  );
  AND2_X1 _53750_ (
    .A1(_18060_),
    .A2(_18065_),
    .ZN(_18066_)
  );
  INV_X1 _53751_ (
    .A(_18066_),
    .ZN(_18067_)
  );
  AND2_X1 _53752_ (
    .A1(_18064_),
    .A2(_18067_),
    .ZN(_01543_)
  );
  AND2_X1 _53753_ (
    .A1(mem_rdata_q[26]),
    .A2(_18031_),
    .ZN(_18068_)
  );
  INV_X1 _53754_ (
    .A(_18068_),
    .ZN(_18069_)
  );
  AND2_X1 _53755_ (
    .A1(instr_jal),
    .A2(decoded_imm_j[6]),
    .ZN(_18070_)
  );
  INV_X1 _53756_ (
    .A(_18070_),
    .ZN(_18071_)
  );
  AND2_X1 _53757_ (
    .A1(_22003_),
    .A2(_02901_),
    .ZN(_18072_)
  );
  INV_X1 _53758_ (
    .A(_18072_),
    .ZN(_18073_)
  );
  AND2_X1 _53759_ (
    .A1(_02900_),
    .A2(_18071_),
    .ZN(_18074_)
  );
  AND2_X1 _53760_ (
    .A1(_18069_),
    .A2(_18074_),
    .ZN(_18075_)
  );
  INV_X1 _53761_ (
    .A(_18075_),
    .ZN(_18076_)
  );
  AND2_X1 _53762_ (
    .A1(_18073_),
    .A2(_18076_),
    .ZN(_01544_)
  );
  AND2_X1 _53763_ (
    .A1(mem_rdata_q[25]),
    .A2(_18031_),
    .ZN(_18077_)
  );
  INV_X1 _53764_ (
    .A(_18077_),
    .ZN(_18078_)
  );
  AND2_X1 _53765_ (
    .A1(instr_jal),
    .A2(decoded_imm_j[5]),
    .ZN(_18079_)
  );
  INV_X1 _53766_ (
    .A(_18079_),
    .ZN(_18080_)
  );
  AND2_X1 _53767_ (
    .A1(_22004_),
    .A2(_02901_),
    .ZN(_18081_)
  );
  INV_X1 _53768_ (
    .A(_18081_),
    .ZN(_18082_)
  );
  AND2_X1 _53769_ (
    .A1(_02900_),
    .A2(_18080_),
    .ZN(_18083_)
  );
  AND2_X1 _53770_ (
    .A1(_18078_),
    .A2(_18083_),
    .ZN(_18084_)
  );
  INV_X1 _53771_ (
    .A(_18084_),
    .ZN(_18085_)
  );
  AND2_X1 _53772_ (
    .A1(_18082_),
    .A2(_18085_),
    .ZN(_01545_)
  );
  AND2_X1 _53773_ (
    .A1(mem_rdata_q[24]),
    .A2(_11684_),
    .ZN(_18086_)
  );
  INV_X1 _53774_ (
    .A(_18086_),
    .ZN(_18087_)
  );
  AND2_X1 _53775_ (
    .A1(instr_jal),
    .A2(decoded_imm_j[4]),
    .ZN(_18088_)
  );
  INV_X1 _53776_ (
    .A(_18088_),
    .ZN(_18089_)
  );
  AND2_X1 _53777_ (
    .A1(mem_rdata_q[11]),
    .A2(_17872_),
    .ZN(_18090_)
  );
  INV_X1 _53778_ (
    .A(_18090_),
    .ZN(_18091_)
  );
  AND2_X1 _53779_ (
    .A1(_22005_),
    .A2(_02901_),
    .ZN(_18092_)
  );
  INV_X1 _53780_ (
    .A(_18092_),
    .ZN(_18093_)
  );
  AND2_X1 _53781_ (
    .A1(_02900_),
    .A2(_18089_),
    .ZN(_18094_)
  );
  AND2_X1 _53782_ (
    .A1(_18087_),
    .A2(_18094_),
    .ZN(_18095_)
  );
  AND2_X1 _53783_ (
    .A1(_18091_),
    .A2(_18095_),
    .ZN(_18096_)
  );
  INV_X1 _53784_ (
    .A(_18096_),
    .ZN(_18097_)
  );
  AND2_X1 _53785_ (
    .A1(_18093_),
    .A2(_18097_),
    .ZN(_01546_)
  );
  AND2_X1 _53786_ (
    .A1(mem_rdata_q[23]),
    .A2(_11684_),
    .ZN(_18098_)
  );
  INV_X1 _53787_ (
    .A(_18098_),
    .ZN(_18099_)
  );
  AND2_X1 _53788_ (
    .A1(mem_rdata_q[10]),
    .A2(_17872_),
    .ZN(_18100_)
  );
  INV_X1 _53789_ (
    .A(_18100_),
    .ZN(_18101_)
  );
  AND2_X1 _53790_ (
    .A1(instr_jal),
    .A2(decoded_rs2[3]),
    .ZN(_18102_)
  );
  INV_X1 _53791_ (
    .A(_18102_),
    .ZN(_18103_)
  );
  AND2_X1 _53792_ (
    .A1(_02900_),
    .A2(_18103_),
    .ZN(_18104_)
  );
  AND2_X1 _53793_ (
    .A1(_18101_),
    .A2(_18104_),
    .ZN(_18105_)
  );
  AND2_X1 _53794_ (
    .A1(_18099_),
    .A2(_18105_),
    .ZN(_18106_)
  );
  INV_X1 _53795_ (
    .A(_18106_),
    .ZN(_18107_)
  );
  AND2_X1 _53796_ (
    .A1(_22006_),
    .A2(_02901_),
    .ZN(_18108_)
  );
  INV_X1 _53797_ (
    .A(_18108_),
    .ZN(_18109_)
  );
  AND2_X1 _53798_ (
    .A1(_18107_),
    .A2(_18109_),
    .ZN(_01547_)
  );
  AND2_X1 _53799_ (
    .A1(mem_rdata_q[22]),
    .A2(_11684_),
    .ZN(_18110_)
  );
  INV_X1 _53800_ (
    .A(_18110_),
    .ZN(_18111_)
  );
  AND2_X1 _53801_ (
    .A1(mem_rdata_q[9]),
    .A2(_17872_),
    .ZN(_18112_)
  );
  INV_X1 _53802_ (
    .A(_18112_),
    .ZN(_18113_)
  );
  AND2_X1 _53803_ (
    .A1(instr_jal),
    .A2(decoded_rs2[2]),
    .ZN(_18114_)
  );
  INV_X1 _53804_ (
    .A(_18114_),
    .ZN(_18115_)
  );
  AND2_X1 _53805_ (
    .A1(_02900_),
    .A2(_18115_),
    .ZN(_18116_)
  );
  AND2_X1 _53806_ (
    .A1(_18113_),
    .A2(_18116_),
    .ZN(_18117_)
  );
  AND2_X1 _53807_ (
    .A1(_18111_),
    .A2(_18117_),
    .ZN(_18118_)
  );
  INV_X1 _53808_ (
    .A(_18118_),
    .ZN(_18119_)
  );
  AND2_X1 _53809_ (
    .A1(_22007_),
    .A2(_02901_),
    .ZN(_18120_)
  );
  INV_X1 _53810_ (
    .A(_18120_),
    .ZN(_18121_)
  );
  AND2_X1 _53811_ (
    .A1(_18119_),
    .A2(_18121_),
    .ZN(_01548_)
  );
  AND2_X1 _53812_ (
    .A1(mem_rdata_q[21]),
    .A2(_11684_),
    .ZN(_18122_)
  );
  INV_X1 _53813_ (
    .A(_18122_),
    .ZN(_18123_)
  );
  AND2_X1 _53814_ (
    .A1(mem_rdata_q[8]),
    .A2(_17872_),
    .ZN(_18124_)
  );
  INV_X1 _53815_ (
    .A(_18124_),
    .ZN(_18125_)
  );
  AND2_X1 _53816_ (
    .A1(_02900_),
    .A2(_03413_),
    .ZN(_18126_)
  );
  AND2_X1 _53817_ (
    .A1(_18125_),
    .A2(_18126_),
    .ZN(_18127_)
  );
  AND2_X1 _53818_ (
    .A1(_18123_),
    .A2(_18127_),
    .ZN(_18128_)
  );
  INV_X1 _53819_ (
    .A(_18128_),
    .ZN(_18129_)
  );
  AND2_X1 _53820_ (
    .A1(_22008_),
    .A2(_02901_),
    .ZN(_18130_)
  );
  INV_X1 _53821_ (
    .A(_18130_),
    .ZN(_18131_)
  );
  AND2_X1 _53822_ (
    .A1(_18129_),
    .A2(_18131_),
    .ZN(_01549_)
  );
  AND2_X1 _53823_ (
    .A1(_00035_),
    .A2(_22317_),
    .ZN(_18132_)
  );
  INV_X1 _53824_ (
    .A(_18132_),
    .ZN(_18133_)
  );
  AND2_X1 _53825_ (
    .A1(_22327_),
    .A2(_18132_),
    .ZN(_01550_)
  );
  INV_X1 _53826_ (
    .A(_01550_),
    .ZN(_18134_)
  );
  AND2_X1 _53827_ (
    .A1(_02464_),
    .A2(_02913_),
    .ZN(_18135_)
  );
  INV_X1 _53828_ (
    .A(_18135_),
    .ZN(_18136_)
  );
  AND2_X1 _53829_ (
    .A1(reg_next_pc[0]),
    .A2(resetn),
    .ZN(_18137_)
  );
  AND2_X1 _53830_ (
    .A1(_18136_),
    .A2(_18137_),
    .ZN(_01551_)
  );
  AND2_X1 _53831_ (
    .A1(_22009_),
    .A2(_11307_),
    .ZN(_18138_)
  );
  INV_X1 _53832_ (
    .A(_18138_),
    .ZN(_18139_)
  );
  AND2_X1 _53833_ (
    .A1(_10496_),
    .A2(_11306_),
    .ZN(_18140_)
  );
  INV_X1 _53834_ (
    .A(_18140_),
    .ZN(_18141_)
  );
  AND2_X1 _53835_ (
    .A1(_18139_),
    .A2(_18141_),
    .ZN(_01552_)
  );
  AND2_X1 _53836_ (
    .A1(_22010_),
    .A2(_11307_),
    .ZN(_18142_)
  );
  INV_X1 _53837_ (
    .A(_18142_),
    .ZN(_18143_)
  );
  AND2_X1 _53838_ (
    .A1(_10491_),
    .A2(_11306_),
    .ZN(_18144_)
  );
  INV_X1 _53839_ (
    .A(_18144_),
    .ZN(_18145_)
  );
  AND2_X1 _53840_ (
    .A1(_18143_),
    .A2(_18145_),
    .ZN(_01553_)
  );
  AND2_X1 _53841_ (
    .A1(_22011_),
    .A2(_11307_),
    .ZN(_18146_)
  );
  INV_X1 _53842_ (
    .A(_18146_),
    .ZN(_18147_)
  );
  AND2_X1 _53843_ (
    .A1(_10486_),
    .A2(_11306_),
    .ZN(_18148_)
  );
  INV_X1 _53844_ (
    .A(_18148_),
    .ZN(_18149_)
  );
  AND2_X1 _53845_ (
    .A1(_18147_),
    .A2(_18149_),
    .ZN(_01554_)
  );
  AND2_X1 _53846_ (
    .A1(_22012_),
    .A2(_11307_),
    .ZN(_18150_)
  );
  INV_X1 _53847_ (
    .A(_18150_),
    .ZN(_18151_)
  );
  AND2_X1 _53848_ (
    .A1(_10501_),
    .A2(_11306_),
    .ZN(_18152_)
  );
  INV_X1 _53849_ (
    .A(_18152_),
    .ZN(_18153_)
  );
  AND2_X1 _53850_ (
    .A1(_18151_),
    .A2(_18153_),
    .ZN(_01555_)
  );
  AND2_X1 _53851_ (
    .A1(_22013_),
    .A2(_11307_),
    .ZN(_18154_)
  );
  INV_X1 _53852_ (
    .A(_18154_),
    .ZN(_18155_)
  );
  AND2_X1 _53853_ (
    .A1(_10506_),
    .A2(_11306_),
    .ZN(_18156_)
  );
  INV_X1 _53854_ (
    .A(_18156_),
    .ZN(_18157_)
  );
  AND2_X1 _53855_ (
    .A1(_18155_),
    .A2(_18157_),
    .ZN(_01556_)
  );
  AND2_X1 _53856_ (
    .A1(_22014_),
    .A2(_11307_),
    .ZN(_18158_)
  );
  INV_X1 _53857_ (
    .A(_18158_),
    .ZN(_18159_)
  );
  AND2_X1 _53858_ (
    .A1(_10516_),
    .A2(_11306_),
    .ZN(_18160_)
  );
  INV_X1 _53859_ (
    .A(_18160_),
    .ZN(_18161_)
  );
  AND2_X1 _53860_ (
    .A1(_18159_),
    .A2(_18161_),
    .ZN(_01557_)
  );
  AND2_X1 _53861_ (
    .A1(_22015_),
    .A2(_11307_),
    .ZN(_18162_)
  );
  INV_X1 _53862_ (
    .A(_18162_),
    .ZN(_18163_)
  );
  AND2_X1 _53863_ (
    .A1(_10481_),
    .A2(_11306_),
    .ZN(_18164_)
  );
  INV_X1 _53864_ (
    .A(_18164_),
    .ZN(_18165_)
  );
  AND2_X1 _53865_ (
    .A1(_18163_),
    .A2(_18165_),
    .ZN(_01558_)
  );
  AND2_X1 _53866_ (
    .A1(_22016_),
    .A2(_11307_),
    .ZN(_18166_)
  );
  INV_X1 _53867_ (
    .A(_18166_),
    .ZN(_18167_)
  );
  AND2_X1 _53868_ (
    .A1(_11417_),
    .A2(_18167_),
    .ZN(_01559_)
  );
  AND2_X1 _53869_ (
    .A1(_22017_),
    .A2(_11307_),
    .ZN(_18168_)
  );
  INV_X1 _53870_ (
    .A(_18168_),
    .ZN(_18169_)
  );
  AND2_X1 _53871_ (
    .A1(_10426_),
    .A2(_11306_),
    .ZN(_18170_)
  );
  INV_X1 _53872_ (
    .A(_18170_),
    .ZN(_18171_)
  );
  AND2_X1 _53873_ (
    .A1(_18169_),
    .A2(_18171_),
    .ZN(_01560_)
  );
  AND2_X1 _53874_ (
    .A1(_10431_),
    .A2(_11306_),
    .ZN(_18172_)
  );
  INV_X1 _53875_ (
    .A(_18172_),
    .ZN(_18173_)
  );
  AND2_X1 _53876_ (
    .A1(_22018_),
    .A2(_11307_),
    .ZN(_18174_)
  );
  INV_X1 _53877_ (
    .A(_18174_),
    .ZN(_18175_)
  );
  AND2_X1 _53878_ (
    .A1(_18173_),
    .A2(_18175_),
    .ZN(_01561_)
  );
  AND2_X1 _53879_ (
    .A1(_22019_),
    .A2(_11307_),
    .ZN(_18176_)
  );
  INV_X1 _53880_ (
    .A(_18176_),
    .ZN(_18177_)
  );
  AND2_X1 _53881_ (
    .A1(_10451_),
    .A2(_11306_),
    .ZN(_18178_)
  );
  INV_X1 _53882_ (
    .A(_18178_),
    .ZN(_18179_)
  );
  AND2_X1 _53883_ (
    .A1(_18177_),
    .A2(_18179_),
    .ZN(_01562_)
  );
  AND2_X1 _53884_ (
    .A1(_22020_),
    .A2(_11307_),
    .ZN(_18180_)
  );
  INV_X1 _53885_ (
    .A(_18180_),
    .ZN(_18181_)
  );
  AND2_X1 _53886_ (
    .A1(_10456_),
    .A2(_11306_),
    .ZN(_18182_)
  );
  INV_X1 _53887_ (
    .A(_18182_),
    .ZN(_18183_)
  );
  AND2_X1 _53888_ (
    .A1(_18181_),
    .A2(_18183_),
    .ZN(_01563_)
  );
  AND2_X1 _53889_ (
    .A1(_22021_),
    .A2(_11307_),
    .ZN(_18184_)
  );
  INV_X1 _53890_ (
    .A(_18184_),
    .ZN(_18185_)
  );
  AND2_X1 _53891_ (
    .A1(_10436_),
    .A2(_11306_),
    .ZN(_18186_)
  );
  INV_X1 _53892_ (
    .A(_18186_),
    .ZN(_18187_)
  );
  AND2_X1 _53893_ (
    .A1(_18185_),
    .A2(_18187_),
    .ZN(_01564_)
  );
  AND2_X1 _53894_ (
    .A1(_22022_),
    .A2(_11307_),
    .ZN(_18188_)
  );
  INV_X1 _53895_ (
    .A(_18188_),
    .ZN(_18189_)
  );
  AND2_X1 _53896_ (
    .A1(_10441_),
    .A2(_11306_),
    .ZN(_18190_)
  );
  INV_X1 _53897_ (
    .A(_18190_),
    .ZN(_18191_)
  );
  AND2_X1 _53898_ (
    .A1(_18189_),
    .A2(_18191_),
    .ZN(_01565_)
  );
  AND2_X1 _53899_ (
    .A1(_22023_),
    .A2(_11307_),
    .ZN(_18192_)
  );
  INV_X1 _53900_ (
    .A(_18192_),
    .ZN(_18193_)
  );
  AND2_X1 _53901_ (
    .A1(_10446_),
    .A2(_11306_),
    .ZN(_18194_)
  );
  INV_X1 _53902_ (
    .A(_18194_),
    .ZN(_18195_)
  );
  AND2_X1 _53903_ (
    .A1(_18193_),
    .A2(_18195_),
    .ZN(_01566_)
  );
  AND2_X1 _53904_ (
    .A1(_22326_),
    .A2(_11107_),
    .ZN(_18196_)
  );
  INV_X1 _53905_ (
    .A(_18196_),
    .ZN(_18197_)
  );
  AND2_X1 _53906_ (
    .A1(_22256_),
    .A2(_18133_),
    .ZN(_18198_)
  );
  INV_X1 _53907_ (
    .A(_18198_),
    .ZN(_18199_)
  );
  AND2_X1 _53908_ (
    .A1(_18197_),
    .A2(_18199_),
    .ZN(_18200_)
  );
  INV_X1 _53909_ (
    .A(_18200_),
    .ZN(_18201_)
  );
  AND2_X1 _53910_ (
    .A1(cpu_state[0]),
    .A2(_18201_),
    .ZN(_18202_)
  );
  INV_X1 _53911_ (
    .A(_18202_),
    .ZN(_18203_)
  );
  AND2_X1 _53912_ (
    .A1(_11141_),
    .A2(_18203_),
    .ZN(_18204_)
  );
  INV_X1 _53913_ (
    .A(_18204_),
    .ZN(_18205_)
  );
  AND2_X1 _53914_ (
    .A1(_21037_),
    .A2(_21103_),
    .ZN(_18206_)
  );
  INV_X1 _53915_ (
    .A(_18206_),
    .ZN(_18207_)
  );
  AND2_X1 _53916_ (
    .A1(_22298_),
    .A2(_18207_),
    .ZN(_18208_)
  );
  INV_X1 _53917_ (
    .A(_18208_),
    .ZN(_18209_)
  );
  AND2_X1 _53918_ (
    .A1(reg_op1[0]),
    .A2(_12198_),
    .ZN(_18210_)
  );
  INV_X1 _53919_ (
    .A(_18210_),
    .ZN(_18211_)
  );
  AND2_X1 _53920_ (
    .A1(_12195_),
    .A2(_18211_),
    .ZN(_18212_)
  );
  INV_X1 _53921_ (
    .A(_18212_),
    .ZN(_18213_)
  );
  AND2_X1 _53922_ (
    .A1(_21168_),
    .A2(_22024_),
    .ZN(_18214_)
  );
  INV_X1 _53923_ (
    .A(_18214_),
    .ZN(_18215_)
  );
  AND2_X1 _53924_ (
    .A1(_22301_),
    .A2(_18215_),
    .ZN(_18216_)
  );
  AND2_X1 _53925_ (
    .A1(_18213_),
    .A2(_18216_),
    .ZN(_18217_)
  );
  INV_X1 _53926_ (
    .A(_18217_),
    .ZN(_18218_)
  );
  AND2_X1 _53927_ (
    .A1(_18209_),
    .A2(_18218_),
    .ZN(_18219_)
  );
  AND2_X1 _53928_ (
    .A1(resetn),
    .A2(_18219_),
    .ZN(_18220_)
  );
  AND2_X1 _53929_ (
    .A1(_18205_),
    .A2(_18220_),
    .ZN(_01567_)
  );
  AND2_X1 _53930_ (
    .A1(_22266_),
    .A2(_18133_),
    .ZN(_18221_)
  );
  INV_X1 _53931_ (
    .A(_18221_),
    .ZN(_18222_)
  );
  AND2_X1 _53932_ (
    .A1(_18197_),
    .A2(_18222_),
    .ZN(_18223_)
  );
  INV_X1 _53933_ (
    .A(_18223_),
    .ZN(_18224_)
  );
  AND2_X1 _53934_ (
    .A1(cpu_state[1]),
    .A2(_18224_),
    .ZN(_18225_)
  );
  INV_X1 _53935_ (
    .A(_18225_),
    .ZN(_18226_)
  );
  AND2_X1 _53936_ (
    .A1(_11144_),
    .A2(_18226_),
    .ZN(_18227_)
  );
  INV_X1 _53937_ (
    .A(_18227_),
    .ZN(_18228_)
  );
  AND2_X1 _53938_ (
    .A1(_18220_),
    .A2(_18228_),
    .ZN(_01568_)
  );
  AND2_X1 _53939_ (
    .A1(is_sll_srl_sra),
    .A2(_05841_),
    .ZN(_18229_)
  );
  INV_X1 _53940_ (
    .A(_18229_),
    .ZN(_18230_)
  );
  AND2_X1 _53941_ (
    .A1(_22296_),
    .A2(_18197_),
    .ZN(_18231_)
  );
  INV_X1 _53942_ (
    .A(_18231_),
    .ZN(_18232_)
  );
  AND2_X1 _53943_ (
    .A1(cpu_state[2]),
    .A2(_18232_),
    .ZN(_18233_)
  );
  INV_X1 _53944_ (
    .A(_18233_),
    .ZN(_18234_)
  );
  AND2_X1 _53945_ (
    .A1(is_slli_srli_srai),
    .A2(_22271_),
    .ZN(_18235_)
  );
  INV_X1 _53946_ (
    .A(_18235_),
    .ZN(_18236_)
  );
  AND2_X1 _53947_ (
    .A1(_18234_),
    .A2(_18236_),
    .ZN(_18237_)
  );
  AND2_X1 _53948_ (
    .A1(_18230_),
    .A2(_18237_),
    .ZN(_18238_)
  );
  INV_X1 _53949_ (
    .A(_18238_),
    .ZN(_18239_)
  );
  AND2_X1 _53950_ (
    .A1(_18220_),
    .A2(_18239_),
    .ZN(_01569_)
  );
  AND2_X1 _53951_ (
    .A1(_21290_),
    .A2(_21291_),
    .ZN(_18240_)
  );
  AND2_X1 _53952_ (
    .A1(_05841_),
    .A2(_18240_),
    .ZN(_18241_)
  );
  INV_X1 _53953_ (
    .A(_18241_),
    .ZN(_18242_)
  );
  AND2_X1 _53954_ (
    .A1(cpu_state[3]),
    .A2(_18196_),
    .ZN(_18243_)
  );
  INV_X1 _53955_ (
    .A(_18243_),
    .ZN(_18244_)
  );
  AND2_X1 _53956_ (
    .A1(cpu_state[3]),
    .A2(_11092_),
    .ZN(_18245_)
  );
  AND2_X1 _53957_ (
    .A1(_22316_),
    .A2(_18245_),
    .ZN(_18246_)
  );
  INV_X1 _53958_ (
    .A(_18246_),
    .ZN(_18247_)
  );
  AND2_X1 _53959_ (
    .A1(_18244_),
    .A2(_18247_),
    .ZN(_18248_)
  );
  AND2_X1 _53960_ (
    .A1(_04967_),
    .A2(_18248_),
    .ZN(_18249_)
  );
  AND2_X1 _53961_ (
    .A1(_18242_),
    .A2(_18249_),
    .ZN(_18250_)
  );
  INV_X1 _53962_ (
    .A(_18250_),
    .ZN(_18251_)
  );
  AND2_X1 _53963_ (
    .A1(_18220_),
    .A2(_18251_),
    .ZN(_01570_)
  );
  AND2_X1 _53964_ (
    .A1(cpu_state[4]),
    .A2(_18220_),
    .ZN(_18252_)
  );
  AND2_X1 _53965_ (
    .A1(_18196_),
    .A2(_18252_),
    .ZN(_01571_)
  );
  AND2_X1 _53966_ (
    .A1(_02464_),
    .A2(_11131_),
    .ZN(_18253_)
  );
  INV_X1 _53967_ (
    .A(_18253_),
    .ZN(_18254_)
  );
  AND2_X1 _53968_ (
    .A1(cpu_state[5]),
    .A2(_18196_),
    .ZN(_18255_)
  );
  INV_X1 _53969_ (
    .A(_18255_),
    .ZN(_18256_)
  );
  AND2_X1 _53970_ (
    .A1(_18254_),
    .A2(_18256_),
    .ZN(_18257_)
  );
  INV_X1 _53971_ (
    .A(_18257_),
    .ZN(_18258_)
  );
  AND2_X1 _53972_ (
    .A1(_18220_),
    .A2(_18258_),
    .ZN(_01572_)
  );
  AND2_X1 _53973_ (
    .A1(_11134_),
    .A2(_18197_),
    .ZN(_18259_)
  );
  INV_X1 _53974_ (
    .A(_18259_),
    .ZN(_18260_)
  );
  AND2_X1 _53975_ (
    .A1(cpu_state[6]),
    .A2(_18260_),
    .ZN(_18261_)
  );
  INV_X1 _53976_ (
    .A(_18261_),
    .ZN(_18262_)
  );
  AND2_X1 _53977_ (
    .A1(is_beq_bne_blt_bge_bltu_bgeu),
    .A2(_22316_),
    .ZN(_18263_)
  );
  INV_X1 _53978_ (
    .A(_18263_),
    .ZN(_18264_)
  );
  AND2_X1 _53979_ (
    .A1(_11090_),
    .A2(_18264_),
    .ZN(_18265_)
  );
  INV_X1 _53980_ (
    .A(_18265_),
    .ZN(_18266_)
  );
  AND2_X1 _53981_ (
    .A1(resetn),
    .A2(_22283_),
    .ZN(_18267_)
  );
  AND2_X1 _53982_ (
    .A1(_11120_),
    .A2(_18267_),
    .ZN(_18268_)
  );
  AND2_X1 _53983_ (
    .A1(_18266_),
    .A2(_18268_),
    .ZN(_18269_)
  );
  AND2_X1 _53984_ (
    .A1(_18134_),
    .A2(_18269_),
    .ZN(_18270_)
  );
  AND2_X1 _53985_ (
    .A1(_18262_),
    .A2(_18270_),
    .ZN(_18271_)
  );
  INV_X1 _53986_ (
    .A(_18271_),
    .ZN(_18272_)
  );
  AND2_X1 _53987_ (
    .A1(_18219_),
    .A2(_18272_),
    .ZN(_01573_)
  );
  AND2_X1 _53988_ (
    .A1(_22035_),
    .A2(_11103_),
    .ZN(_18273_)
  );
  INV_X1 _53989_ (
    .A(_18273_),
    .ZN(_18274_)
  );
  AND2_X1 _53990_ (
    .A1(resetn),
    .A2(_18274_),
    .ZN(_18275_)
  );
  INV_X1 _53991_ (
    .A(_18275_),
    .ZN(_18276_)
  );
  AND2_X1 _53992_ (
    .A1(_18219_),
    .A2(_18276_),
    .ZN(_18277_)
  );
  INV_X1 _53993_ (
    .A(_18277_),
    .ZN(_01574_)
  );
  AND2_X1 _53994_ (
    .A1(reg_pc[1]),
    .A2(_22335_),
    .ZN(_18278_)
  );
  INV_X1 _53995_ (
    .A(_18278_),
    .ZN(_18279_)
  );
  AND2_X1 _53996_ (
    .A1(\cpuregs[26] [1]),
    .A2(_22149_),
    .ZN(_18280_)
  );
  INV_X1 _53997_ (
    .A(_18280_),
    .ZN(_18281_)
  );
  AND2_X1 _53998_ (
    .A1(\cpuregs[30] [1]),
    .A2(_00008_[2]),
    .ZN(_18282_)
  );
  INV_X1 _53999_ (
    .A(_18282_),
    .ZN(_18283_)
  );
  AND2_X1 _54000_ (
    .A1(_22147_),
    .A2(_18283_),
    .ZN(_18284_)
  );
  AND2_X1 _54001_ (
    .A1(_18281_),
    .A2(_18284_),
    .ZN(_18285_)
  );
  INV_X1 _54002_ (
    .A(_18285_),
    .ZN(_18286_)
  );
  AND2_X1 _54003_ (
    .A1(\cpuregs[31] [1]),
    .A2(_00008_[2]),
    .ZN(_18287_)
  );
  INV_X1 _54004_ (
    .A(_18287_),
    .ZN(_18288_)
  );
  AND2_X1 _54005_ (
    .A1(\cpuregs[27] [1]),
    .A2(_22149_),
    .ZN(_18289_)
  );
  INV_X1 _54006_ (
    .A(_18289_),
    .ZN(_18290_)
  );
  AND2_X1 _54007_ (
    .A1(_00008_[0]),
    .A2(_18290_),
    .ZN(_18291_)
  );
  AND2_X1 _54008_ (
    .A1(_18288_),
    .A2(_18291_),
    .ZN(_18292_)
  );
  INV_X1 _54009_ (
    .A(_18292_),
    .ZN(_18293_)
  );
  AND2_X1 _54010_ (
    .A1(_18286_),
    .A2(_18293_),
    .ZN(_18294_)
  );
  AND2_X1 _54011_ (
    .A1(\cpuregs[18] [1]),
    .A2(_22149_),
    .ZN(_18295_)
  );
  INV_X1 _54012_ (
    .A(_18295_),
    .ZN(_18296_)
  );
  AND2_X1 _54013_ (
    .A1(\cpuregs[22] [1]),
    .A2(_00008_[2]),
    .ZN(_18297_)
  );
  INV_X1 _54014_ (
    .A(_18297_),
    .ZN(_18298_)
  );
  AND2_X1 _54015_ (
    .A1(_22147_),
    .A2(_18298_),
    .ZN(_18299_)
  );
  AND2_X1 _54016_ (
    .A1(_18296_),
    .A2(_18299_),
    .ZN(_18300_)
  );
  INV_X1 _54017_ (
    .A(_18300_),
    .ZN(_18301_)
  );
  AND2_X1 _54018_ (
    .A1(\cpuregs[19] [1]),
    .A2(_22149_),
    .ZN(_18302_)
  );
  INV_X1 _54019_ (
    .A(_18302_),
    .ZN(_18303_)
  );
  AND2_X1 _54020_ (
    .A1(\cpuregs[23] [1]),
    .A2(_00008_[2]),
    .ZN(_18304_)
  );
  INV_X1 _54021_ (
    .A(_18304_),
    .ZN(_18305_)
  );
  AND2_X1 _54022_ (
    .A1(_00008_[0]),
    .A2(_18305_),
    .ZN(_18306_)
  );
  AND2_X1 _54023_ (
    .A1(_18303_),
    .A2(_18306_),
    .ZN(_18307_)
  );
  INV_X1 _54024_ (
    .A(_18307_),
    .ZN(_18308_)
  );
  AND2_X1 _54025_ (
    .A1(_00008_[3]),
    .A2(_18294_),
    .ZN(_18309_)
  );
  INV_X1 _54026_ (
    .A(_18309_),
    .ZN(_18310_)
  );
  AND2_X1 _54027_ (
    .A1(_22150_),
    .A2(_18308_),
    .ZN(_18311_)
  );
  AND2_X1 _54028_ (
    .A1(_18301_),
    .A2(_18311_),
    .ZN(_18312_)
  );
  INV_X1 _54029_ (
    .A(_18312_),
    .ZN(_18313_)
  );
  AND2_X1 _54030_ (
    .A1(_18310_),
    .A2(_18313_),
    .ZN(_18314_)
  );
  INV_X1 _54031_ (
    .A(_18314_),
    .ZN(_18315_)
  );
  AND2_X1 _54032_ (
    .A1(_21834_),
    .A2(_22149_),
    .ZN(_18316_)
  );
  INV_X1 _54033_ (
    .A(_18316_),
    .ZN(_18317_)
  );
  AND2_X1 _54034_ (
    .A1(_21890_),
    .A2(_00008_[2]),
    .ZN(_18318_)
  );
  INV_X1 _54035_ (
    .A(_18318_),
    .ZN(_18319_)
  );
  AND2_X1 _54036_ (
    .A1(_21568_),
    .A2(_22149_),
    .ZN(_18320_)
  );
  INV_X1 _54037_ (
    .A(_18320_),
    .ZN(_18321_)
  );
  AND2_X1 _54038_ (
    .A1(_21906_),
    .A2(_00008_[2]),
    .ZN(_18322_)
  );
  INV_X1 _54039_ (
    .A(_18322_),
    .ZN(_18323_)
  );
  AND2_X1 _54040_ (
    .A1(_18321_),
    .A2(_18323_),
    .ZN(_18324_)
  );
  AND2_X1 _54041_ (
    .A1(_00008_[0]),
    .A2(_18319_),
    .ZN(_18325_)
  );
  AND2_X1 _54042_ (
    .A1(_18317_),
    .A2(_18325_),
    .ZN(_18326_)
  );
  INV_X1 _54043_ (
    .A(_18326_),
    .ZN(_18327_)
  );
  AND2_X1 _54044_ (
    .A1(_22147_),
    .A2(_18324_),
    .ZN(_18328_)
  );
  INV_X1 _54045_ (
    .A(_18328_),
    .ZN(_18329_)
  );
  AND2_X1 _54046_ (
    .A1(_18327_),
    .A2(_18329_),
    .ZN(_18330_)
  );
  AND2_X1 _54047_ (
    .A1(_00008_[3]),
    .A2(_18330_),
    .ZN(_18331_)
  );
  INV_X1 _54048_ (
    .A(_18331_),
    .ZN(_18332_)
  );
  AND2_X1 _54049_ (
    .A1(\cpuregs[20] [1]),
    .A2(_00008_[2]),
    .ZN(_18333_)
  );
  INV_X1 _54050_ (
    .A(_18333_),
    .ZN(_18334_)
  );
  AND2_X1 _54051_ (
    .A1(\cpuregs[16] [1]),
    .A2(_22149_),
    .ZN(_18335_)
  );
  INV_X1 _54052_ (
    .A(_18335_),
    .ZN(_18336_)
  );
  AND2_X1 _54053_ (
    .A1(_18334_),
    .A2(_18336_),
    .ZN(_18337_)
  );
  AND2_X1 _54054_ (
    .A1(_22147_),
    .A2(_18337_),
    .ZN(_18338_)
  );
  INV_X1 _54055_ (
    .A(_18338_),
    .ZN(_18339_)
  );
  AND2_X1 _54056_ (
    .A1(\cpuregs[21] [1]),
    .A2(_00008_[2]),
    .ZN(_18340_)
  );
  INV_X1 _54057_ (
    .A(_18340_),
    .ZN(_18341_)
  );
  AND2_X1 _54058_ (
    .A1(\cpuregs[17] [1]),
    .A2(_22149_),
    .ZN(_18342_)
  );
  INV_X1 _54059_ (
    .A(_18342_),
    .ZN(_18343_)
  );
  AND2_X1 _54060_ (
    .A1(_00008_[0]),
    .A2(_18343_),
    .ZN(_18344_)
  );
  AND2_X1 _54061_ (
    .A1(_18341_),
    .A2(_18344_),
    .ZN(_18345_)
  );
  INV_X1 _54062_ (
    .A(_18345_),
    .ZN(_18346_)
  );
  AND2_X1 _54063_ (
    .A1(_18339_),
    .A2(_18346_),
    .ZN(_18347_)
  );
  INV_X1 _54064_ (
    .A(_18347_),
    .ZN(_18348_)
  );
  AND2_X1 _54065_ (
    .A1(_22150_),
    .A2(_18348_),
    .ZN(_18349_)
  );
  INV_X1 _54066_ (
    .A(_18349_),
    .ZN(_18350_)
  );
  AND2_X1 _54067_ (
    .A1(_22148_),
    .A2(_18332_),
    .ZN(_18351_)
  );
  AND2_X1 _54068_ (
    .A1(_18350_),
    .A2(_18351_),
    .ZN(_18352_)
  );
  INV_X1 _54069_ (
    .A(_18352_),
    .ZN(_18353_)
  );
  AND2_X1 _54070_ (
    .A1(_00008_[1]),
    .A2(_18315_),
    .ZN(_18354_)
  );
  INV_X1 _54071_ (
    .A(_18354_),
    .ZN(_18355_)
  );
  AND2_X1 _54072_ (
    .A1(_00008_[4]),
    .A2(_18355_),
    .ZN(_18356_)
  );
  AND2_X1 _54073_ (
    .A1(_18353_),
    .A2(_18356_),
    .ZN(_18357_)
  );
  INV_X1 _54074_ (
    .A(_18357_),
    .ZN(_18358_)
  );
  AND2_X1 _54075_ (
    .A1(_21780_),
    .A2(_00008_[2]),
    .ZN(_18359_)
  );
  INV_X1 _54076_ (
    .A(_18359_),
    .ZN(_18360_)
  );
  AND2_X1 _54077_ (
    .A1(_21488_),
    .A2(_22149_),
    .ZN(_18361_)
  );
  INV_X1 _54078_ (
    .A(_18361_),
    .ZN(_18362_)
  );
  AND2_X1 _54079_ (
    .A1(_21538_),
    .A2(_22149_),
    .ZN(_18363_)
  );
  INV_X1 _54080_ (
    .A(_18363_),
    .ZN(_18364_)
  );
  AND2_X1 _54081_ (
    .A1(_21805_),
    .A2(_00008_[2]),
    .ZN(_18365_)
  );
  INV_X1 _54082_ (
    .A(_18365_),
    .ZN(_18366_)
  );
  AND2_X1 _54083_ (
    .A1(_18364_),
    .A2(_18366_),
    .ZN(_18367_)
  );
  AND2_X1 _54084_ (
    .A1(_00008_[0]),
    .A2(_18362_),
    .ZN(_18368_)
  );
  AND2_X1 _54085_ (
    .A1(_18360_),
    .A2(_18368_),
    .ZN(_18369_)
  );
  INV_X1 _54086_ (
    .A(_18369_),
    .ZN(_18370_)
  );
  AND2_X1 _54087_ (
    .A1(_22147_),
    .A2(_18367_),
    .ZN(_18371_)
  );
  INV_X1 _54088_ (
    .A(_18371_),
    .ZN(_18372_)
  );
  AND2_X1 _54089_ (
    .A1(_18370_),
    .A2(_18372_),
    .ZN(_18373_)
  );
  AND2_X1 _54090_ (
    .A1(_00008_[1]),
    .A2(_18373_),
    .ZN(_18374_)
  );
  INV_X1 _54091_ (
    .A(_18374_),
    .ZN(_18375_)
  );
  AND2_X1 _54092_ (
    .A1(_21513_),
    .A2(_22149_),
    .ZN(_18376_)
  );
  INV_X1 _54093_ (
    .A(_18376_),
    .ZN(_18377_)
  );
  AND2_X1 _54094_ (
    .A1(_21733_),
    .A2(_00008_[2]),
    .ZN(_18378_)
  );
  INV_X1 _54095_ (
    .A(_18378_),
    .ZN(_18379_)
  );
  AND2_X1 _54096_ (
    .A1(_21954_),
    .A2(_22149_),
    .ZN(_18380_)
  );
  INV_X1 _54097_ (
    .A(_18380_),
    .ZN(_18381_)
  );
  AND2_X1 _54098_ (
    .A1(_21670_),
    .A2(_00008_[2]),
    .ZN(_18382_)
  );
  INV_X1 _54099_ (
    .A(_18382_),
    .ZN(_18383_)
  );
  AND2_X1 _54100_ (
    .A1(_18381_),
    .A2(_18383_),
    .ZN(_18384_)
  );
  AND2_X1 _54101_ (
    .A1(_00008_[0]),
    .A2(_18377_),
    .ZN(_18385_)
  );
  AND2_X1 _54102_ (
    .A1(_18379_),
    .A2(_18385_),
    .ZN(_18386_)
  );
  INV_X1 _54103_ (
    .A(_18386_),
    .ZN(_18387_)
  );
  AND2_X1 _54104_ (
    .A1(_22147_),
    .A2(_18384_),
    .ZN(_18388_)
  );
  INV_X1 _54105_ (
    .A(_18388_),
    .ZN(_18389_)
  );
  AND2_X1 _54106_ (
    .A1(_18387_),
    .A2(_18389_),
    .ZN(_18390_)
  );
  AND2_X1 _54107_ (
    .A1(_22148_),
    .A2(_18390_),
    .ZN(_18391_)
  );
  INV_X1 _54108_ (
    .A(_18391_),
    .ZN(_18392_)
  );
  AND2_X1 _54109_ (
    .A1(_18375_),
    .A2(_18392_),
    .ZN(_18393_)
  );
  INV_X1 _54110_ (
    .A(_18393_),
    .ZN(_18394_)
  );
  AND2_X1 _54111_ (
    .A1(_22150_),
    .A2(_18394_),
    .ZN(_18395_)
  );
  INV_X1 _54112_ (
    .A(_18395_),
    .ZN(_18396_)
  );
  AND2_X1 _54113_ (
    .A1(\cpuregs[9] [1]),
    .A2(_22148_),
    .ZN(_18397_)
  );
  INV_X1 _54114_ (
    .A(_18397_),
    .ZN(_18398_)
  );
  AND2_X1 _54115_ (
    .A1(\cpuregs[11] [1]),
    .A2(_00008_[1]),
    .ZN(_18399_)
  );
  INV_X1 _54116_ (
    .A(_18399_),
    .ZN(_18400_)
  );
  AND2_X1 _54117_ (
    .A1(_22149_),
    .A2(_18400_),
    .ZN(_18401_)
  );
  AND2_X1 _54118_ (
    .A1(_18398_),
    .A2(_18401_),
    .ZN(_18402_)
  );
  INV_X1 _54119_ (
    .A(_18402_),
    .ZN(_18403_)
  );
  AND2_X1 _54120_ (
    .A1(\cpuregs[13] [1]),
    .A2(_22148_),
    .ZN(_18404_)
  );
  INV_X1 _54121_ (
    .A(_18404_),
    .ZN(_18405_)
  );
  AND2_X1 _54122_ (
    .A1(\cpuregs[15] [1]),
    .A2(_00008_[1]),
    .ZN(_18406_)
  );
  INV_X1 _54123_ (
    .A(_18406_),
    .ZN(_18407_)
  );
  AND2_X1 _54124_ (
    .A1(_00008_[2]),
    .A2(_18407_),
    .ZN(_18408_)
  );
  AND2_X1 _54125_ (
    .A1(_18405_),
    .A2(_18408_),
    .ZN(_18409_)
  );
  INV_X1 _54126_ (
    .A(_18409_),
    .ZN(_18410_)
  );
  AND2_X1 _54127_ (
    .A1(_18403_),
    .A2(_18410_),
    .ZN(_18411_)
  );
  INV_X1 _54128_ (
    .A(_18411_),
    .ZN(_18412_)
  );
  AND2_X1 _54129_ (
    .A1(_00008_[0]),
    .A2(_18412_),
    .ZN(_18413_)
  );
  INV_X1 _54130_ (
    .A(_18413_),
    .ZN(_18414_)
  );
  AND2_X1 _54131_ (
    .A1(\cpuregs[8] [1]),
    .A2(_22148_),
    .ZN(_18415_)
  );
  INV_X1 _54132_ (
    .A(_18415_),
    .ZN(_18416_)
  );
  AND2_X1 _54133_ (
    .A1(\cpuregs[10] [1]),
    .A2(_00008_[1]),
    .ZN(_18417_)
  );
  INV_X1 _54134_ (
    .A(_18417_),
    .ZN(_18418_)
  );
  AND2_X1 _54135_ (
    .A1(_22149_),
    .A2(_18418_),
    .ZN(_18419_)
  );
  AND2_X1 _54136_ (
    .A1(_18416_),
    .A2(_18419_),
    .ZN(_18420_)
  );
  INV_X1 _54137_ (
    .A(_18420_),
    .ZN(_18421_)
  );
  AND2_X1 _54138_ (
    .A1(\cpuregs[12] [1]),
    .A2(_22148_),
    .ZN(_18422_)
  );
  INV_X1 _54139_ (
    .A(_18422_),
    .ZN(_18423_)
  );
  AND2_X1 _54140_ (
    .A1(\cpuregs[14] [1]),
    .A2(_00008_[1]),
    .ZN(_18424_)
  );
  INV_X1 _54141_ (
    .A(_18424_),
    .ZN(_18425_)
  );
  AND2_X1 _54142_ (
    .A1(_00008_[2]),
    .A2(_18425_),
    .ZN(_18426_)
  );
  AND2_X1 _54143_ (
    .A1(_18423_),
    .A2(_18426_),
    .ZN(_18427_)
  );
  INV_X1 _54144_ (
    .A(_18427_),
    .ZN(_18428_)
  );
  AND2_X1 _54145_ (
    .A1(_18421_),
    .A2(_18428_),
    .ZN(_18429_)
  );
  INV_X1 _54146_ (
    .A(_18429_),
    .ZN(_18430_)
  );
  AND2_X1 _54147_ (
    .A1(_22147_),
    .A2(_18430_),
    .ZN(_18431_)
  );
  INV_X1 _54148_ (
    .A(_18431_),
    .ZN(_18432_)
  );
  AND2_X1 _54149_ (
    .A1(_18414_),
    .A2(_18432_),
    .ZN(_18433_)
  );
  INV_X1 _54150_ (
    .A(_18433_),
    .ZN(_18434_)
  );
  AND2_X1 _54151_ (
    .A1(_00008_[3]),
    .A2(_18434_),
    .ZN(_18435_)
  );
  INV_X1 _54152_ (
    .A(_18435_),
    .ZN(_18436_)
  );
  AND2_X1 _54153_ (
    .A1(_18396_),
    .A2(_18436_),
    .ZN(_18437_)
  );
  INV_X1 _54154_ (
    .A(_18437_),
    .ZN(_18438_)
  );
  AND2_X1 _54155_ (
    .A1(_22151_),
    .A2(_18438_),
    .ZN(_18439_)
  );
  INV_X1 _54156_ (
    .A(_18439_),
    .ZN(_18440_)
  );
  AND2_X1 _54157_ (
    .A1(_22546_),
    .A2(_18358_),
    .ZN(_18441_)
  );
  AND2_X1 _54158_ (
    .A1(_18440_),
    .A2(_18441_),
    .ZN(_18442_)
  );
  INV_X1 _54159_ (
    .A(_18442_),
    .ZN(_18443_)
  );
  AND2_X1 _54160_ (
    .A1(_18279_),
    .A2(_18443_),
    .ZN(_18444_)
  );
  INV_X1 _54161_ (
    .A(_18444_),
    .ZN(_18445_)
  );
  AND2_X1 _54162_ (
    .A1(_22271_),
    .A2(_18445_),
    .ZN(_18446_)
  );
  INV_X1 _54163_ (
    .A(_18446_),
    .ZN(_18447_)
  );
  AND2_X1 _54164_ (
    .A1(_22561_),
    .A2(_22766_),
    .ZN(_18448_)
  );
  INV_X1 _54165_ (
    .A(_18448_),
    .ZN(_18449_)
  );
  AND2_X1 _54166_ (
    .A1(reg_op1[2]),
    .A2(_22290_),
    .ZN(_18450_)
  );
  INV_X1 _54167_ (
    .A(_18450_),
    .ZN(_18451_)
  );
  AND2_X1 _54168_ (
    .A1(_23202_),
    .A2(_18451_),
    .ZN(_18452_)
  );
  AND2_X1 _54169_ (
    .A1(_22024_),
    .A2(_22334_),
    .ZN(_18453_)
  );
  INV_X1 _54170_ (
    .A(_18453_),
    .ZN(_18454_)
  );
  AND2_X1 _54171_ (
    .A1(_22572_),
    .A2(_18452_),
    .ZN(_18455_)
  );
  INV_X1 _54172_ (
    .A(_18455_),
    .ZN(_18456_)
  );
  AND2_X1 _54173_ (
    .A1(_22573_),
    .A2(_23197_),
    .ZN(_18457_)
  );
  INV_X1 _54174_ (
    .A(_18457_),
    .ZN(_18458_)
  );
  AND2_X1 _54175_ (
    .A1(_22295_),
    .A2(_18458_),
    .ZN(_18459_)
  );
  AND2_X1 _54176_ (
    .A1(_18456_),
    .A2(_18459_),
    .ZN(_18460_)
  );
  INV_X1 _54177_ (
    .A(_18460_),
    .ZN(_18461_)
  );
  AND2_X1 _54178_ (
    .A1(_22559_),
    .A2(_18449_),
    .ZN(_18462_)
  );
  AND2_X1 _54179_ (
    .A1(_22768_),
    .A2(_18462_),
    .ZN(_18463_)
  );
  INV_X1 _54180_ (
    .A(_18463_),
    .ZN(_18464_)
  );
  AND2_X1 _54181_ (
    .A1(_18461_),
    .A2(_18464_),
    .ZN(_18465_)
  );
  AND2_X1 _54182_ (
    .A1(_22333_),
    .A2(_18465_),
    .ZN(_18466_)
  );
  AND2_X1 _54183_ (
    .A1(_18447_),
    .A2(_18466_),
    .ZN(_18467_)
  );
  INV_X1 _54184_ (
    .A(_18467_),
    .ZN(_18468_)
  );
  AND2_X1 _54185_ (
    .A1(_18454_),
    .A2(_18468_),
    .ZN(_01575_)
  );
  AND2_X1 _54186_ (
    .A1(_21060_),
    .A2(_22504_),
    .ZN(_18469_)
  );
  INV_X1 _54187_ (
    .A(_18469_),
    .ZN(_00003_)
  );
  AND2_X1 _54188_ (
    .A1(_21058_),
    .A2(_22505_),
    .ZN(_18470_)
  );
  INV_X1 _54189_ (
    .A(_18470_),
    .ZN(_00004_)
  );
  AND2_X1 _54190_ (
    .A1(_11763_),
    .A2(_11766_),
    .ZN(mem_la_read)
  );
  AND2_X1 _54191_ (
    .A1(_22326_),
    .A2(_11093_),
    .ZN(_18471_)
  );
  INV_X1 _54192_ (
    .A(_18471_),
    .ZN(_18472_)
  );
  AND2_X1 _54193_ (
    .A1(_11307_),
    .A2(_18134_),
    .ZN(_18473_)
  );
  INV_X1 _54194_ (
    .A(_18473_),
    .ZN(_18474_)
  );
  AND2_X1 _54195_ (
    .A1(_18472_),
    .A2(_18474_),
    .ZN(_00000_)
  );
  AND2_X1 _54196_ (
    .A1(_21064_),
    .A2(_21065_),
    .ZN(_18475_)
  );
  INV_X1 _54197_ (
    .A(_18475_),
    .ZN(_18476_)
  );
  AND2_X1 _54198_ (
    .A1(_21063_),
    .A2(_18475_),
    .ZN(_18477_)
  );
  INV_X1 _54199_ (
    .A(_18477_),
    .ZN(_18478_)
  );
  AND2_X1 _54200_ (
    .A1(_22256_),
    .A2(_18132_),
    .ZN(_18479_)
  );
  AND2_X1 _54201_ (
    .A1(_18478_),
    .A2(_18479_),
    .ZN(_18480_)
  );
  AND2_X1 _54202_ (
    .A1(_12196_),
    .A2(_18214_),
    .ZN(_18481_)
  );
  INV_X1 _54203_ (
    .A(_18481_),
    .ZN(_18482_)
  );
  AND2_X1 _54204_ (
    .A1(_12474_),
    .A2(_18482_),
    .ZN(_18483_)
  );
  INV_X1 _54205_ (
    .A(_18483_),
    .ZN(_18484_)
  );
  AND2_X1 _54206_ (
    .A1(mem_rdata[0]),
    .A2(_18484_),
    .ZN(_18485_)
  );
  INV_X1 _54207_ (
    .A(_18485_),
    .ZN(_18486_)
  );
  AND2_X1 _54208_ (
    .A1(_21168_),
    .A2(_22064_),
    .ZN(_18487_)
  );
  AND2_X1 _54209_ (
    .A1(_12196_),
    .A2(_18487_),
    .ZN(_18488_)
  );
  INV_X1 _54210_ (
    .A(_18488_),
    .ZN(_18489_)
  );
  AND2_X1 _54211_ (
    .A1(_12495_),
    .A2(_18489_),
    .ZN(_18490_)
  );
  INV_X1 _54212_ (
    .A(_18490_),
    .ZN(_18491_)
  );
  AND2_X1 _54213_ (
    .A1(mem_rdata[16]),
    .A2(_18491_),
    .ZN(_18492_)
  );
  INV_X1 _54214_ (
    .A(_18492_),
    .ZN(_18493_)
  );
  AND2_X1 _54215_ (
    .A1(_22063_),
    .A2(_22064_),
    .ZN(_18494_)
  );
  AND2_X1 _54216_ (
    .A1(mem_rdata[24]),
    .A2(_18494_),
    .ZN(_18495_)
  );
  INV_X1 _54217_ (
    .A(_18495_),
    .ZN(_18496_)
  );
  AND2_X1 _54218_ (
    .A1(_22024_),
    .A2(_22063_),
    .ZN(_18497_)
  );
  AND2_X1 _54219_ (
    .A1(mem_rdata[8]),
    .A2(_18497_),
    .ZN(_18498_)
  );
  INV_X1 _54220_ (
    .A(_18498_),
    .ZN(_18499_)
  );
  AND2_X1 _54221_ (
    .A1(_18496_),
    .A2(_18499_),
    .ZN(_18500_)
  );
  INV_X1 _54222_ (
    .A(_18500_),
    .ZN(_18501_)
  );
  AND2_X1 _54223_ (
    .A1(_12196_),
    .A2(_18501_),
    .ZN(_18502_)
  );
  INV_X1 _54224_ (
    .A(_18502_),
    .ZN(_18503_)
  );
  AND2_X1 _54225_ (
    .A1(_18493_),
    .A2(_18503_),
    .ZN(_18504_)
  );
  AND2_X1 _54226_ (
    .A1(_18486_),
    .A2(_18504_),
    .ZN(_18505_)
  );
  INV_X1 _54227_ (
    .A(_18505_),
    .ZN(_18506_)
  );
  AND2_X1 _54228_ (
    .A1(_18480_),
    .A2(_18506_),
    .ZN(_18507_)
  );
  INV_X1 _54229_ (
    .A(_18507_),
    .ZN(_18508_)
  );
  AND2_X1 _54230_ (
    .A1(reg_op1[0]),
    .A2(_22282_),
    .ZN(_18509_)
  );
  INV_X1 _54231_ (
    .A(_18509_),
    .ZN(_18510_)
  );
  AND2_X1 _54232_ (
    .A1(count_instr[32]),
    .A2(instr_rdinstrh),
    .ZN(_18511_)
  );
  INV_X1 _54233_ (
    .A(_18511_),
    .ZN(_18512_)
  );
  AND2_X1 _54234_ (
    .A1(count_instr[0]),
    .A2(instr_rdinstr),
    .ZN(_18513_)
  );
  INV_X1 _54235_ (
    .A(_18513_),
    .ZN(_18514_)
  );
  AND2_X1 _54236_ (
    .A1(_18512_),
    .A2(_18514_),
    .ZN(_18515_)
  );
  AND2_X1 _54237_ (
    .A1(instr_rdcycle),
    .A2(count_cycle[0]),
    .ZN(_18516_)
  );
  INV_X1 _54238_ (
    .A(_18516_),
    .ZN(_18517_)
  );
  AND2_X1 _54239_ (
    .A1(instr_rdcycleh),
    .A2(count_cycle[32]),
    .ZN(_18518_)
  );
  INV_X1 _54240_ (
    .A(_18518_),
    .ZN(_18519_)
  );
  AND2_X1 _54241_ (
    .A1(_18517_),
    .A2(_18519_),
    .ZN(_18520_)
  );
  AND2_X1 _54242_ (
    .A1(_18515_),
    .A2(_18520_),
    .ZN(_18521_)
  );
  INV_X1 _54243_ (
    .A(_18521_),
    .ZN(_18522_)
  );
  AND2_X1 _54244_ (
    .A1(_22271_),
    .A2(_18522_),
    .ZN(_18523_)
  );
  INV_X1 _54245_ (
    .A(_18523_),
    .ZN(_18524_)
  );
  AND2_X1 _54246_ (
    .A1(reg_next_pc[0]),
    .A2(decoded_imm[0]),
    .ZN(_18525_)
  );
  INV_X1 _54247_ (
    .A(_18525_),
    .ZN(_18526_)
  );
  AND2_X1 _54248_ (
    .A1(_21037_),
    .A2(_21286_),
    .ZN(_18527_)
  );
  INV_X1 _54249_ (
    .A(_18527_),
    .ZN(_18528_)
  );
  AND2_X1 _54250_ (
    .A1(_18526_),
    .A2(_18528_),
    .ZN(_18529_)
  );
  AND2_X1 _54251_ (
    .A1(_11090_),
    .A2(_18529_),
    .ZN(_18530_)
  );
  INV_X1 _54252_ (
    .A(_18530_),
    .ZN(_18531_)
  );
  AND2_X1 _54253_ (
    .A1(_18524_),
    .A2(_18531_),
    .ZN(_18532_)
  );
  AND2_X1 _54254_ (
    .A1(_18510_),
    .A2(_18532_),
    .ZN(_18533_)
  );
  AND2_X1 _54255_ (
    .A1(_18508_),
    .A2(_18533_),
    .ZN(_18534_)
  );
  INV_X1 _54256_ (
    .A(_18534_),
    .ZN(_18535_)
  );
  AND2_X1 _54257_ (
    .A1(resetn),
    .A2(_18535_),
    .ZN(_00005_[0])
  );
  AND2_X1 _54258_ (
    .A1(mem_rdata[1]),
    .A2(_18484_),
    .ZN(_18536_)
  );
  INV_X1 _54259_ (
    .A(_18536_),
    .ZN(_18537_)
  );
  AND2_X1 _54260_ (
    .A1(mem_rdata[17]),
    .A2(_18491_),
    .ZN(_18538_)
  );
  INV_X1 _54261_ (
    .A(_18538_),
    .ZN(_18539_)
  );
  AND2_X1 _54262_ (
    .A1(mem_rdata[25]),
    .A2(_18494_),
    .ZN(_18540_)
  );
  INV_X1 _54263_ (
    .A(_18540_),
    .ZN(_18541_)
  );
  AND2_X1 _54264_ (
    .A1(mem_rdata[9]),
    .A2(_18497_),
    .ZN(_18542_)
  );
  INV_X1 _54265_ (
    .A(_18542_),
    .ZN(_18543_)
  );
  AND2_X1 _54266_ (
    .A1(_18541_),
    .A2(_18543_),
    .ZN(_18544_)
  );
  INV_X1 _54267_ (
    .A(_18544_),
    .ZN(_18545_)
  );
  AND2_X1 _54268_ (
    .A1(_12196_),
    .A2(_18545_),
    .ZN(_18546_)
  );
  INV_X1 _54269_ (
    .A(_18546_),
    .ZN(_18547_)
  );
  AND2_X1 _54270_ (
    .A1(_18539_),
    .A2(_18547_),
    .ZN(_18548_)
  );
  AND2_X1 _54271_ (
    .A1(_18537_),
    .A2(_18548_),
    .ZN(_18549_)
  );
  INV_X1 _54272_ (
    .A(_18549_),
    .ZN(_18550_)
  );
  AND2_X1 _54273_ (
    .A1(_18480_),
    .A2(_18550_),
    .ZN(_18551_)
  );
  INV_X1 _54274_ (
    .A(_18551_),
    .ZN(_18552_)
  );
  AND2_X1 _54275_ (
    .A1(reg_pc[1]),
    .A2(decoded_imm[1]),
    .ZN(_18553_)
  );
  INV_X1 _54276_ (
    .A(_18553_),
    .ZN(_18554_)
  );
  AND2_X1 _54277_ (
    .A1(_21103_),
    .A2(_22008_),
    .ZN(_18555_)
  );
  INV_X1 _54278_ (
    .A(_18555_),
    .ZN(_18556_)
  );
  AND2_X1 _54279_ (
    .A1(_18554_),
    .A2(_18556_),
    .ZN(_18557_)
  );
  INV_X1 _54280_ (
    .A(_18557_),
    .ZN(_18558_)
  );
  AND2_X1 _54281_ (
    .A1(_18526_),
    .A2(_18558_),
    .ZN(_18559_)
  );
  INV_X1 _54282_ (
    .A(_18559_),
    .ZN(_18560_)
  );
  AND2_X1 _54283_ (
    .A1(_18525_),
    .A2(_18557_),
    .ZN(_18561_)
  );
  INV_X1 _54284_ (
    .A(_18561_),
    .ZN(_18562_)
  );
  AND2_X1 _54285_ (
    .A1(_11090_),
    .A2(_18562_),
    .ZN(_18563_)
  );
  AND2_X1 _54286_ (
    .A1(_18560_),
    .A2(_18563_),
    .ZN(_18564_)
  );
  INV_X1 _54287_ (
    .A(_18564_),
    .ZN(_18565_)
  );
  AND2_X1 _54288_ (
    .A1(reg_op1[1]),
    .A2(_22282_),
    .ZN(_18566_)
  );
  INV_X1 _54289_ (
    .A(_18566_),
    .ZN(_18567_)
  );
  AND2_X1 _54290_ (
    .A1(instr_rdcycle),
    .A2(count_cycle[1]),
    .ZN(_18568_)
  );
  INV_X1 _54291_ (
    .A(_18568_),
    .ZN(_18569_)
  );
  AND2_X1 _54292_ (
    .A1(count_instr[33]),
    .A2(instr_rdinstrh),
    .ZN(_18570_)
  );
  INV_X1 _54293_ (
    .A(_18570_),
    .ZN(_18571_)
  );
  AND2_X1 _54294_ (
    .A1(_18569_),
    .A2(_18571_),
    .ZN(_18572_)
  );
  AND2_X1 _54295_ (
    .A1(count_instr[1]),
    .A2(instr_rdinstr),
    .ZN(_18573_)
  );
  INV_X1 _54296_ (
    .A(_18573_),
    .ZN(_18574_)
  );
  AND2_X1 _54297_ (
    .A1(instr_rdcycleh),
    .A2(count_cycle[33]),
    .ZN(_18575_)
  );
  INV_X1 _54298_ (
    .A(_18575_),
    .ZN(_18576_)
  );
  AND2_X1 _54299_ (
    .A1(_18574_),
    .A2(_18576_),
    .ZN(_18577_)
  );
  AND2_X1 _54300_ (
    .A1(_18572_),
    .A2(_18577_),
    .ZN(_18578_)
  );
  INV_X1 _54301_ (
    .A(_18578_),
    .ZN(_18579_)
  );
  AND2_X1 _54302_ (
    .A1(_22271_),
    .A2(_18579_),
    .ZN(_18580_)
  );
  INV_X1 _54303_ (
    .A(_18580_),
    .ZN(_18581_)
  );
  AND2_X1 _54304_ (
    .A1(_18567_),
    .A2(_18581_),
    .ZN(_18582_)
  );
  AND2_X1 _54305_ (
    .A1(_18565_),
    .A2(_18582_),
    .ZN(_18583_)
  );
  AND2_X1 _54306_ (
    .A1(_18552_),
    .A2(_18583_),
    .ZN(_18584_)
  );
  INV_X1 _54307_ (
    .A(_18584_),
    .ZN(_18585_)
  );
  AND2_X1 _54308_ (
    .A1(resetn),
    .A2(_18585_),
    .ZN(_00005_[1])
  );
  AND2_X1 _54309_ (
    .A1(mem_rdata[2]),
    .A2(_18484_),
    .ZN(_18586_)
  );
  INV_X1 _54310_ (
    .A(_18586_),
    .ZN(_18587_)
  );
  AND2_X1 _54311_ (
    .A1(mem_rdata[18]),
    .A2(_18491_),
    .ZN(_18588_)
  );
  INV_X1 _54312_ (
    .A(_18588_),
    .ZN(_18589_)
  );
  AND2_X1 _54313_ (
    .A1(mem_rdata[26]),
    .A2(_18494_),
    .ZN(_18590_)
  );
  INV_X1 _54314_ (
    .A(_18590_),
    .ZN(_18591_)
  );
  AND2_X1 _54315_ (
    .A1(mem_rdata[10]),
    .A2(_18497_),
    .ZN(_18592_)
  );
  INV_X1 _54316_ (
    .A(_18592_),
    .ZN(_18593_)
  );
  AND2_X1 _54317_ (
    .A1(_18591_),
    .A2(_18593_),
    .ZN(_18594_)
  );
  INV_X1 _54318_ (
    .A(_18594_),
    .ZN(_18595_)
  );
  AND2_X1 _54319_ (
    .A1(_12196_),
    .A2(_18595_),
    .ZN(_18596_)
  );
  INV_X1 _54320_ (
    .A(_18596_),
    .ZN(_18597_)
  );
  AND2_X1 _54321_ (
    .A1(_18589_),
    .A2(_18597_),
    .ZN(_18598_)
  );
  AND2_X1 _54322_ (
    .A1(_18587_),
    .A2(_18598_),
    .ZN(_18599_)
  );
  INV_X1 _54323_ (
    .A(_18599_),
    .ZN(_18600_)
  );
  AND2_X1 _54324_ (
    .A1(_18480_),
    .A2(_18600_),
    .ZN(_18601_)
  );
  INV_X1 _54325_ (
    .A(_18601_),
    .ZN(_18602_)
  );
  AND2_X1 _54326_ (
    .A1(_18554_),
    .A2(_18562_),
    .ZN(_18603_)
  );
  INV_X1 _54327_ (
    .A(_18603_),
    .ZN(_18604_)
  );
  AND2_X1 _54328_ (
    .A1(reg_pc[2]),
    .A2(decoded_imm[2]),
    .ZN(_18605_)
  );
  INV_X1 _54329_ (
    .A(_18605_),
    .ZN(_18606_)
  );
  AND2_X1 _54330_ (
    .A1(_21102_),
    .A2(_22007_),
    .ZN(_18607_)
  );
  INV_X1 _54331_ (
    .A(_18607_),
    .ZN(_18608_)
  );
  AND2_X1 _54332_ (
    .A1(_18606_),
    .A2(_18608_),
    .ZN(_18609_)
  );
  INV_X1 _54333_ (
    .A(_18609_),
    .ZN(_18610_)
  );
  AND2_X1 _54334_ (
    .A1(_18604_),
    .A2(_18609_),
    .ZN(_18611_)
  );
  INV_X1 _54335_ (
    .A(_18611_),
    .ZN(_18612_)
  );
  AND2_X1 _54336_ (
    .A1(_18603_),
    .A2(_18610_),
    .ZN(_18613_)
  );
  INV_X1 _54337_ (
    .A(_18613_),
    .ZN(_18614_)
  );
  AND2_X1 _54338_ (
    .A1(_11090_),
    .A2(_18614_),
    .ZN(_18615_)
  );
  AND2_X1 _54339_ (
    .A1(_18612_),
    .A2(_18615_),
    .ZN(_18616_)
  );
  INV_X1 _54340_ (
    .A(_18616_),
    .ZN(_18617_)
  );
  AND2_X1 _54341_ (
    .A1(reg_op1[2]),
    .A2(_22282_),
    .ZN(_18618_)
  );
  INV_X1 _54342_ (
    .A(_18618_),
    .ZN(_18619_)
  );
  AND2_X1 _54343_ (
    .A1(instr_rdcycle),
    .A2(count_cycle[2]),
    .ZN(_18620_)
  );
  INV_X1 _54344_ (
    .A(_18620_),
    .ZN(_18621_)
  );
  AND2_X1 _54345_ (
    .A1(instr_rdcycleh),
    .A2(count_cycle[34]),
    .ZN(_18622_)
  );
  INV_X1 _54346_ (
    .A(_18622_),
    .ZN(_18623_)
  );
  AND2_X1 _54347_ (
    .A1(_18621_),
    .A2(_18623_),
    .ZN(_18624_)
  );
  AND2_X1 _54348_ (
    .A1(count_instr[2]),
    .A2(instr_rdinstr),
    .ZN(_18625_)
  );
  INV_X1 _54349_ (
    .A(_18625_),
    .ZN(_18626_)
  );
  AND2_X1 _54350_ (
    .A1(count_instr[34]),
    .A2(instr_rdinstrh),
    .ZN(_18627_)
  );
  INV_X1 _54351_ (
    .A(_18627_),
    .ZN(_18628_)
  );
  AND2_X1 _54352_ (
    .A1(_18626_),
    .A2(_18628_),
    .ZN(_18629_)
  );
  AND2_X1 _54353_ (
    .A1(_18624_),
    .A2(_18629_),
    .ZN(_18630_)
  );
  INV_X1 _54354_ (
    .A(_18630_),
    .ZN(_18631_)
  );
  AND2_X1 _54355_ (
    .A1(_22271_),
    .A2(_18631_),
    .ZN(_18632_)
  );
  INV_X1 _54356_ (
    .A(_18632_),
    .ZN(_18633_)
  );
  AND2_X1 _54357_ (
    .A1(_18619_),
    .A2(_18633_),
    .ZN(_18634_)
  );
  AND2_X1 _54358_ (
    .A1(_18617_),
    .A2(_18634_),
    .ZN(_18635_)
  );
  AND2_X1 _54359_ (
    .A1(_18602_),
    .A2(_18635_),
    .ZN(_18636_)
  );
  INV_X1 _54360_ (
    .A(_18636_),
    .ZN(_18637_)
  );
  AND2_X1 _54361_ (
    .A1(resetn),
    .A2(_18637_),
    .ZN(_00005_[2])
  );
  AND2_X1 _54362_ (
    .A1(_18606_),
    .A2(_18612_),
    .ZN(_18638_)
  );
  INV_X1 _54363_ (
    .A(_18638_),
    .ZN(_18639_)
  );
  AND2_X1 _54364_ (
    .A1(reg_pc[3]),
    .A2(decoded_imm[3]),
    .ZN(_18640_)
  );
  INV_X1 _54365_ (
    .A(_18640_),
    .ZN(_18641_)
  );
  AND2_X1 _54366_ (
    .A1(_21101_),
    .A2(_22006_),
    .ZN(_18642_)
  );
  INV_X1 _54367_ (
    .A(_18642_),
    .ZN(_18643_)
  );
  AND2_X1 _54368_ (
    .A1(_18641_),
    .A2(_18643_),
    .ZN(_18644_)
  );
  INV_X1 _54369_ (
    .A(_18644_),
    .ZN(_18645_)
  );
  AND2_X1 _54370_ (
    .A1(_18639_),
    .A2(_18644_),
    .ZN(_18646_)
  );
  INV_X1 _54371_ (
    .A(_18646_),
    .ZN(_18647_)
  );
  AND2_X1 _54372_ (
    .A1(_18638_),
    .A2(_18645_),
    .ZN(_18648_)
  );
  INV_X1 _54373_ (
    .A(_18648_),
    .ZN(_18649_)
  );
  AND2_X1 _54374_ (
    .A1(_11090_),
    .A2(_18649_),
    .ZN(_18650_)
  );
  AND2_X1 _54375_ (
    .A1(_18647_),
    .A2(_18650_),
    .ZN(_18651_)
  );
  INV_X1 _54376_ (
    .A(_18651_),
    .ZN(_18652_)
  );
  AND2_X1 _54377_ (
    .A1(mem_rdata[3]),
    .A2(_18484_),
    .ZN(_18653_)
  );
  INV_X1 _54378_ (
    .A(_18653_),
    .ZN(_18654_)
  );
  AND2_X1 _54379_ (
    .A1(mem_rdata[27]),
    .A2(_18494_),
    .ZN(_18655_)
  );
  INV_X1 _54380_ (
    .A(_18655_),
    .ZN(_18656_)
  );
  AND2_X1 _54381_ (
    .A1(mem_rdata[11]),
    .A2(_18497_),
    .ZN(_18657_)
  );
  INV_X1 _54382_ (
    .A(_18657_),
    .ZN(_18658_)
  );
  AND2_X1 _54383_ (
    .A1(_18656_),
    .A2(_18658_),
    .ZN(_18659_)
  );
  INV_X1 _54384_ (
    .A(_18659_),
    .ZN(_18660_)
  );
  AND2_X1 _54385_ (
    .A1(_12196_),
    .A2(_18660_),
    .ZN(_18661_)
  );
  INV_X1 _54386_ (
    .A(_18661_),
    .ZN(_18662_)
  );
  AND2_X1 _54387_ (
    .A1(mem_rdata[19]),
    .A2(_18491_),
    .ZN(_18663_)
  );
  INV_X1 _54388_ (
    .A(_18663_),
    .ZN(_18664_)
  );
  AND2_X1 _54389_ (
    .A1(_18662_),
    .A2(_18664_),
    .ZN(_18665_)
  );
  AND2_X1 _54390_ (
    .A1(_18654_),
    .A2(_18665_),
    .ZN(_18666_)
  );
  INV_X1 _54391_ (
    .A(_18666_),
    .ZN(_18667_)
  );
  AND2_X1 _54392_ (
    .A1(_18480_),
    .A2(_18667_),
    .ZN(_18668_)
  );
  INV_X1 _54393_ (
    .A(_18668_),
    .ZN(_18669_)
  );
  AND2_X1 _54394_ (
    .A1(reg_op1[3]),
    .A2(_22282_),
    .ZN(_18670_)
  );
  INV_X1 _54395_ (
    .A(_18670_),
    .ZN(_18671_)
  );
  AND2_X1 _54396_ (
    .A1(instr_rdcycle),
    .A2(count_cycle[3]),
    .ZN(_18672_)
  );
  INV_X1 _54397_ (
    .A(_18672_),
    .ZN(_18673_)
  );
  AND2_X1 _54398_ (
    .A1(instr_rdcycleh),
    .A2(count_cycle[35]),
    .ZN(_18674_)
  );
  INV_X1 _54399_ (
    .A(_18674_),
    .ZN(_18675_)
  );
  AND2_X1 _54400_ (
    .A1(_18673_),
    .A2(_18675_),
    .ZN(_18676_)
  );
  AND2_X1 _54401_ (
    .A1(count_instr[35]),
    .A2(instr_rdinstrh),
    .ZN(_18677_)
  );
  INV_X1 _54402_ (
    .A(_18677_),
    .ZN(_18678_)
  );
  AND2_X1 _54403_ (
    .A1(count_instr[3]),
    .A2(instr_rdinstr),
    .ZN(_18679_)
  );
  INV_X1 _54404_ (
    .A(_18679_),
    .ZN(_18680_)
  );
  AND2_X1 _54405_ (
    .A1(_18678_),
    .A2(_18680_),
    .ZN(_18681_)
  );
  AND2_X1 _54406_ (
    .A1(_18676_),
    .A2(_18681_),
    .ZN(_18682_)
  );
  INV_X1 _54407_ (
    .A(_18682_),
    .ZN(_18683_)
  );
  AND2_X1 _54408_ (
    .A1(_22271_),
    .A2(_18683_),
    .ZN(_18684_)
  );
  INV_X1 _54409_ (
    .A(_18684_),
    .ZN(_18685_)
  );
  AND2_X1 _54410_ (
    .A1(_18671_),
    .A2(_18685_),
    .ZN(_18686_)
  );
  AND2_X1 _54411_ (
    .A1(_18669_),
    .A2(_18686_),
    .ZN(_18687_)
  );
  AND2_X1 _54412_ (
    .A1(_18652_),
    .A2(_18687_),
    .ZN(_18688_)
  );
  INV_X1 _54413_ (
    .A(_18688_),
    .ZN(_18689_)
  );
  AND2_X1 _54414_ (
    .A1(resetn),
    .A2(_18689_),
    .ZN(_00005_[3])
  );
  AND2_X1 _54415_ (
    .A1(_18641_),
    .A2(_18647_),
    .ZN(_18690_)
  );
  INV_X1 _54416_ (
    .A(_18690_),
    .ZN(_18691_)
  );
  AND2_X1 _54417_ (
    .A1(reg_pc[4]),
    .A2(decoded_imm[4]),
    .ZN(_18692_)
  );
  INV_X1 _54418_ (
    .A(_18692_),
    .ZN(_18693_)
  );
  AND2_X1 _54419_ (
    .A1(_21100_),
    .A2(_22005_),
    .ZN(_18694_)
  );
  INV_X1 _54420_ (
    .A(_18694_),
    .ZN(_18695_)
  );
  AND2_X1 _54421_ (
    .A1(_18693_),
    .A2(_18695_),
    .ZN(_18696_)
  );
  INV_X1 _54422_ (
    .A(_18696_),
    .ZN(_18697_)
  );
  AND2_X1 _54423_ (
    .A1(_18691_),
    .A2(_18696_),
    .ZN(_18698_)
  );
  INV_X1 _54424_ (
    .A(_18698_),
    .ZN(_18699_)
  );
  AND2_X1 _54425_ (
    .A1(_18690_),
    .A2(_18697_),
    .ZN(_18700_)
  );
  INV_X1 _54426_ (
    .A(_18700_),
    .ZN(_18701_)
  );
  AND2_X1 _54427_ (
    .A1(_11090_),
    .A2(_18701_),
    .ZN(_18702_)
  );
  AND2_X1 _54428_ (
    .A1(_18699_),
    .A2(_18702_),
    .ZN(_18703_)
  );
  INV_X1 _54429_ (
    .A(_18703_),
    .ZN(_18704_)
  );
  AND2_X1 _54430_ (
    .A1(mem_rdata[4]),
    .A2(_18484_),
    .ZN(_18705_)
  );
  INV_X1 _54431_ (
    .A(_18705_),
    .ZN(_18706_)
  );
  AND2_X1 _54432_ (
    .A1(mem_rdata[28]),
    .A2(_18494_),
    .ZN(_18707_)
  );
  INV_X1 _54433_ (
    .A(_18707_),
    .ZN(_18708_)
  );
  AND2_X1 _54434_ (
    .A1(mem_rdata[12]),
    .A2(_18497_),
    .ZN(_18709_)
  );
  INV_X1 _54435_ (
    .A(_18709_),
    .ZN(_18710_)
  );
  AND2_X1 _54436_ (
    .A1(_18708_),
    .A2(_18710_),
    .ZN(_18711_)
  );
  INV_X1 _54437_ (
    .A(_18711_),
    .ZN(_18712_)
  );
  AND2_X1 _54438_ (
    .A1(_12196_),
    .A2(_18712_),
    .ZN(_18713_)
  );
  INV_X1 _54439_ (
    .A(_18713_),
    .ZN(_18714_)
  );
  AND2_X1 _54440_ (
    .A1(mem_rdata[20]),
    .A2(_18491_),
    .ZN(_18715_)
  );
  INV_X1 _54441_ (
    .A(_18715_),
    .ZN(_18716_)
  );
  AND2_X1 _54442_ (
    .A1(_18714_),
    .A2(_18716_),
    .ZN(_18717_)
  );
  AND2_X1 _54443_ (
    .A1(_18706_),
    .A2(_18717_),
    .ZN(_18718_)
  );
  INV_X1 _54444_ (
    .A(_18718_),
    .ZN(_18719_)
  );
  AND2_X1 _54445_ (
    .A1(_18480_),
    .A2(_18719_),
    .ZN(_18720_)
  );
  INV_X1 _54446_ (
    .A(_18720_),
    .ZN(_18721_)
  );
  AND2_X1 _54447_ (
    .A1(count_instr[36]),
    .A2(instr_rdinstrh),
    .ZN(_18722_)
  );
  INV_X1 _54448_ (
    .A(_18722_),
    .ZN(_18723_)
  );
  AND2_X1 _54449_ (
    .A1(count_instr[4]),
    .A2(instr_rdinstr),
    .ZN(_18724_)
  );
  INV_X1 _54450_ (
    .A(_18724_),
    .ZN(_18725_)
  );
  AND2_X1 _54451_ (
    .A1(_18723_),
    .A2(_18725_),
    .ZN(_18726_)
  );
  AND2_X1 _54452_ (
    .A1(instr_rdcycle),
    .A2(count_cycle[4]),
    .ZN(_18727_)
  );
  INV_X1 _54453_ (
    .A(_18727_),
    .ZN(_18728_)
  );
  AND2_X1 _54454_ (
    .A1(instr_rdcycleh),
    .A2(count_cycle[36]),
    .ZN(_18729_)
  );
  INV_X1 _54455_ (
    .A(_18729_),
    .ZN(_18730_)
  );
  AND2_X1 _54456_ (
    .A1(_18728_),
    .A2(_18730_),
    .ZN(_18731_)
  );
  AND2_X1 _54457_ (
    .A1(_18726_),
    .A2(_18731_),
    .ZN(_18732_)
  );
  INV_X1 _54458_ (
    .A(_18732_),
    .ZN(_18733_)
  );
  AND2_X1 _54459_ (
    .A1(_22271_),
    .A2(_18733_),
    .ZN(_18734_)
  );
  INV_X1 _54460_ (
    .A(_18734_),
    .ZN(_18735_)
  );
  AND2_X1 _54461_ (
    .A1(reg_op1[4]),
    .A2(_22282_),
    .ZN(_18736_)
  );
  INV_X1 _54462_ (
    .A(_18736_),
    .ZN(_18737_)
  );
  AND2_X1 _54463_ (
    .A1(_18735_),
    .A2(_18737_),
    .ZN(_18738_)
  );
  AND2_X1 _54464_ (
    .A1(_18721_),
    .A2(_18738_),
    .ZN(_18739_)
  );
  AND2_X1 _54465_ (
    .A1(_18704_),
    .A2(_18739_),
    .ZN(_18740_)
  );
  INV_X1 _54466_ (
    .A(_18740_),
    .ZN(_18741_)
  );
  AND2_X1 _54467_ (
    .A1(resetn),
    .A2(_18741_),
    .ZN(_00005_[4])
  );
  AND2_X1 _54468_ (
    .A1(_18693_),
    .A2(_18699_),
    .ZN(_18742_)
  );
  INV_X1 _54469_ (
    .A(_18742_),
    .ZN(_18743_)
  );
  AND2_X1 _54470_ (
    .A1(reg_pc[5]),
    .A2(decoded_imm[5]),
    .ZN(_18744_)
  );
  INV_X1 _54471_ (
    .A(_18744_),
    .ZN(_18745_)
  );
  AND2_X1 _54472_ (
    .A1(_21099_),
    .A2(_22004_),
    .ZN(_18746_)
  );
  INV_X1 _54473_ (
    .A(_18746_),
    .ZN(_18747_)
  );
  AND2_X1 _54474_ (
    .A1(_18745_),
    .A2(_18747_),
    .ZN(_18748_)
  );
  INV_X1 _54475_ (
    .A(_18748_),
    .ZN(_18749_)
  );
  AND2_X1 _54476_ (
    .A1(_18742_),
    .A2(_18749_),
    .ZN(_18750_)
  );
  INV_X1 _54477_ (
    .A(_18750_),
    .ZN(_18751_)
  );
  AND2_X1 _54478_ (
    .A1(_18743_),
    .A2(_18748_),
    .ZN(_18752_)
  );
  INV_X1 _54479_ (
    .A(_18752_),
    .ZN(_18753_)
  );
  AND2_X1 _54480_ (
    .A1(_11090_),
    .A2(_18751_),
    .ZN(_18754_)
  );
  AND2_X1 _54481_ (
    .A1(_18753_),
    .A2(_18754_),
    .ZN(_18755_)
  );
  INV_X1 _54482_ (
    .A(_18755_),
    .ZN(_18756_)
  );
  AND2_X1 _54483_ (
    .A1(mem_rdata[5]),
    .A2(_18484_),
    .ZN(_18757_)
  );
  INV_X1 _54484_ (
    .A(_18757_),
    .ZN(_18758_)
  );
  AND2_X1 _54485_ (
    .A1(mem_rdata[29]),
    .A2(_18494_),
    .ZN(_18759_)
  );
  INV_X1 _54486_ (
    .A(_18759_),
    .ZN(_18760_)
  );
  AND2_X1 _54487_ (
    .A1(mem_rdata[13]),
    .A2(_18497_),
    .ZN(_18761_)
  );
  INV_X1 _54488_ (
    .A(_18761_),
    .ZN(_18762_)
  );
  AND2_X1 _54489_ (
    .A1(_18760_),
    .A2(_18762_),
    .ZN(_18763_)
  );
  INV_X1 _54490_ (
    .A(_18763_),
    .ZN(_18764_)
  );
  AND2_X1 _54491_ (
    .A1(_12196_),
    .A2(_18764_),
    .ZN(_18765_)
  );
  INV_X1 _54492_ (
    .A(_18765_),
    .ZN(_18766_)
  );
  AND2_X1 _54493_ (
    .A1(mem_rdata[21]),
    .A2(_18491_),
    .ZN(_18767_)
  );
  INV_X1 _54494_ (
    .A(_18767_),
    .ZN(_18768_)
  );
  AND2_X1 _54495_ (
    .A1(_18766_),
    .A2(_18768_),
    .ZN(_18769_)
  );
  AND2_X1 _54496_ (
    .A1(_18758_),
    .A2(_18769_),
    .ZN(_18770_)
  );
  INV_X1 _54497_ (
    .A(_18770_),
    .ZN(_18771_)
  );
  AND2_X1 _54498_ (
    .A1(_18480_),
    .A2(_18771_),
    .ZN(_18772_)
  );
  INV_X1 _54499_ (
    .A(_18772_),
    .ZN(_18773_)
  );
  AND2_X1 _54500_ (
    .A1(instr_rdcycleh),
    .A2(count_cycle[37]),
    .ZN(_18774_)
  );
  INV_X1 _54501_ (
    .A(_18774_),
    .ZN(_18775_)
  );
  AND2_X1 _54502_ (
    .A1(count_instr[5]),
    .A2(instr_rdinstr),
    .ZN(_18776_)
  );
  INV_X1 _54503_ (
    .A(_18776_),
    .ZN(_18777_)
  );
  AND2_X1 _54504_ (
    .A1(_18775_),
    .A2(_18777_),
    .ZN(_18778_)
  );
  AND2_X1 _54505_ (
    .A1(instr_rdcycle),
    .A2(count_cycle[5]),
    .ZN(_18779_)
  );
  INV_X1 _54506_ (
    .A(_18779_),
    .ZN(_18780_)
  );
  AND2_X1 _54507_ (
    .A1(count_instr[37]),
    .A2(instr_rdinstrh),
    .ZN(_18781_)
  );
  INV_X1 _54508_ (
    .A(_18781_),
    .ZN(_18782_)
  );
  AND2_X1 _54509_ (
    .A1(_18780_),
    .A2(_18782_),
    .ZN(_18783_)
  );
  AND2_X1 _54510_ (
    .A1(_18778_),
    .A2(_18783_),
    .ZN(_18784_)
  );
  INV_X1 _54511_ (
    .A(_18784_),
    .ZN(_18785_)
  );
  AND2_X1 _54512_ (
    .A1(_22271_),
    .A2(_18785_),
    .ZN(_18786_)
  );
  INV_X1 _54513_ (
    .A(_18786_),
    .ZN(_18787_)
  );
  AND2_X1 _54514_ (
    .A1(reg_op1[5]),
    .A2(_22282_),
    .ZN(_18788_)
  );
  INV_X1 _54515_ (
    .A(_18788_),
    .ZN(_18789_)
  );
  AND2_X1 _54516_ (
    .A1(_18773_),
    .A2(_18787_),
    .ZN(_18790_)
  );
  AND2_X1 _54517_ (
    .A1(_18789_),
    .A2(_18790_),
    .ZN(_18791_)
  );
  AND2_X1 _54518_ (
    .A1(_18756_),
    .A2(_18791_),
    .ZN(_18792_)
  );
  INV_X1 _54519_ (
    .A(_18792_),
    .ZN(_18793_)
  );
  AND2_X1 _54520_ (
    .A1(resetn),
    .A2(_18793_),
    .ZN(_00005_[5])
  );
  AND2_X1 _54521_ (
    .A1(_18745_),
    .A2(_18753_),
    .ZN(_18794_)
  );
  INV_X1 _54522_ (
    .A(_18794_),
    .ZN(_18795_)
  );
  AND2_X1 _54523_ (
    .A1(reg_pc[6]),
    .A2(decoded_imm[6]),
    .ZN(_18796_)
  );
  INV_X1 _54524_ (
    .A(_18796_),
    .ZN(_18797_)
  );
  AND2_X1 _54525_ (
    .A1(_21098_),
    .A2(_22003_),
    .ZN(_18798_)
  );
  INV_X1 _54526_ (
    .A(_18798_),
    .ZN(_18799_)
  );
  AND2_X1 _54527_ (
    .A1(_18797_),
    .A2(_18799_),
    .ZN(_18800_)
  );
  INV_X1 _54528_ (
    .A(_18800_),
    .ZN(_18801_)
  );
  AND2_X1 _54529_ (
    .A1(_18795_),
    .A2(_18800_),
    .ZN(_18802_)
  );
  INV_X1 _54530_ (
    .A(_18802_),
    .ZN(_18803_)
  );
  AND2_X1 _54531_ (
    .A1(_18794_),
    .A2(_18801_),
    .ZN(_18804_)
  );
  INV_X1 _54532_ (
    .A(_18804_),
    .ZN(_18805_)
  );
  AND2_X1 _54533_ (
    .A1(_11090_),
    .A2(_18805_),
    .ZN(_18806_)
  );
  AND2_X1 _54534_ (
    .A1(_18803_),
    .A2(_18806_),
    .ZN(_18807_)
  );
  INV_X1 _54535_ (
    .A(_18807_),
    .ZN(_18808_)
  );
  AND2_X1 _54536_ (
    .A1(mem_rdata[6]),
    .A2(_18484_),
    .ZN(_18809_)
  );
  INV_X1 _54537_ (
    .A(_18809_),
    .ZN(_18810_)
  );
  AND2_X1 _54538_ (
    .A1(mem_rdata[30]),
    .A2(_18494_),
    .ZN(_18811_)
  );
  INV_X1 _54539_ (
    .A(_18811_),
    .ZN(_18812_)
  );
  AND2_X1 _54540_ (
    .A1(mem_rdata[14]),
    .A2(_18497_),
    .ZN(_18813_)
  );
  INV_X1 _54541_ (
    .A(_18813_),
    .ZN(_18814_)
  );
  AND2_X1 _54542_ (
    .A1(_18812_),
    .A2(_18814_),
    .ZN(_18815_)
  );
  INV_X1 _54543_ (
    .A(_18815_),
    .ZN(_18816_)
  );
  AND2_X1 _54544_ (
    .A1(_12196_),
    .A2(_18816_),
    .ZN(_18817_)
  );
  INV_X1 _54545_ (
    .A(_18817_),
    .ZN(_18818_)
  );
  AND2_X1 _54546_ (
    .A1(mem_rdata[22]),
    .A2(_18491_),
    .ZN(_18819_)
  );
  INV_X1 _54547_ (
    .A(_18819_),
    .ZN(_18820_)
  );
  AND2_X1 _54548_ (
    .A1(_18818_),
    .A2(_18820_),
    .ZN(_18821_)
  );
  AND2_X1 _54549_ (
    .A1(_18810_),
    .A2(_18821_),
    .ZN(_18822_)
  );
  INV_X1 _54550_ (
    .A(_18822_),
    .ZN(_18823_)
  );
  AND2_X1 _54551_ (
    .A1(_18480_),
    .A2(_18823_),
    .ZN(_18824_)
  );
  INV_X1 _54552_ (
    .A(_18824_),
    .ZN(_18825_)
  );
  AND2_X1 _54553_ (
    .A1(reg_op1[6]),
    .A2(_22282_),
    .ZN(_18826_)
  );
  INV_X1 _54554_ (
    .A(_18826_),
    .ZN(_18827_)
  );
  AND2_X1 _54555_ (
    .A1(instr_rdcycleh),
    .A2(count_cycle[38]),
    .ZN(_18828_)
  );
  INV_X1 _54556_ (
    .A(_18828_),
    .ZN(_18829_)
  );
  AND2_X1 _54557_ (
    .A1(count_instr[6]),
    .A2(instr_rdinstr),
    .ZN(_18830_)
  );
  INV_X1 _54558_ (
    .A(_18830_),
    .ZN(_18831_)
  );
  AND2_X1 _54559_ (
    .A1(_18829_),
    .A2(_18831_),
    .ZN(_18832_)
  );
  AND2_X1 _54560_ (
    .A1(instr_rdcycle),
    .A2(count_cycle[6]),
    .ZN(_18833_)
  );
  INV_X1 _54561_ (
    .A(_18833_),
    .ZN(_18834_)
  );
  AND2_X1 _54562_ (
    .A1(count_instr[38]),
    .A2(instr_rdinstrh),
    .ZN(_18835_)
  );
  INV_X1 _54563_ (
    .A(_18835_),
    .ZN(_18836_)
  );
  AND2_X1 _54564_ (
    .A1(_18834_),
    .A2(_18836_),
    .ZN(_18837_)
  );
  AND2_X1 _54565_ (
    .A1(_18832_),
    .A2(_18837_),
    .ZN(_18838_)
  );
  INV_X1 _54566_ (
    .A(_18838_),
    .ZN(_18839_)
  );
  AND2_X1 _54567_ (
    .A1(_22271_),
    .A2(_18839_),
    .ZN(_18840_)
  );
  INV_X1 _54568_ (
    .A(_18840_),
    .ZN(_18841_)
  );
  AND2_X1 _54569_ (
    .A1(_18827_),
    .A2(_18841_),
    .ZN(_18842_)
  );
  AND2_X1 _54570_ (
    .A1(_18825_),
    .A2(_18842_),
    .ZN(_18843_)
  );
  AND2_X1 _54571_ (
    .A1(_18808_),
    .A2(_18843_),
    .ZN(_18844_)
  );
  INV_X1 _54572_ (
    .A(_18844_),
    .ZN(_18845_)
  );
  AND2_X1 _54573_ (
    .A1(resetn),
    .A2(_18845_),
    .ZN(_00005_[6])
  );
  AND2_X1 _54574_ (
    .A1(mem_rdata[7]),
    .A2(_18484_),
    .ZN(_18846_)
  );
  INV_X1 _54575_ (
    .A(_18846_),
    .ZN(_18847_)
  );
  AND2_X1 _54576_ (
    .A1(mem_rdata[31]),
    .A2(_18494_),
    .ZN(_18848_)
  );
  INV_X1 _54577_ (
    .A(_18848_),
    .ZN(_18849_)
  );
  AND2_X1 _54578_ (
    .A1(mem_rdata[15]),
    .A2(_18497_),
    .ZN(_18850_)
  );
  INV_X1 _54579_ (
    .A(_18850_),
    .ZN(_18851_)
  );
  AND2_X1 _54580_ (
    .A1(_18849_),
    .A2(_18851_),
    .ZN(_18852_)
  );
  INV_X1 _54581_ (
    .A(_18852_),
    .ZN(_18853_)
  );
  AND2_X1 _54582_ (
    .A1(_12196_),
    .A2(_18853_),
    .ZN(_18854_)
  );
  INV_X1 _54583_ (
    .A(_18854_),
    .ZN(_18855_)
  );
  AND2_X1 _54584_ (
    .A1(mem_rdata[23]),
    .A2(_18491_),
    .ZN(_18856_)
  );
  INV_X1 _54585_ (
    .A(_18856_),
    .ZN(_18857_)
  );
  AND2_X1 _54586_ (
    .A1(_18855_),
    .A2(_18857_),
    .ZN(_18858_)
  );
  AND2_X1 _54587_ (
    .A1(_18847_),
    .A2(_18858_),
    .ZN(_18859_)
  );
  INV_X1 _54588_ (
    .A(_18859_),
    .ZN(_18860_)
  );
  AND2_X1 _54589_ (
    .A1(_18480_),
    .A2(_18860_),
    .ZN(_18861_)
  );
  INV_X1 _54590_ (
    .A(_18861_),
    .ZN(_18862_)
  );
  AND2_X1 _54591_ (
    .A1(reg_op1[7]),
    .A2(_22282_),
    .ZN(_18863_)
  );
  INV_X1 _54592_ (
    .A(_18863_),
    .ZN(_18864_)
  );
  AND2_X1 _54593_ (
    .A1(count_instr[39]),
    .A2(instr_rdinstrh),
    .ZN(_18865_)
  );
  INV_X1 _54594_ (
    .A(_18865_),
    .ZN(_18866_)
  );
  AND2_X1 _54595_ (
    .A1(count_instr[7]),
    .A2(instr_rdinstr),
    .ZN(_18867_)
  );
  INV_X1 _54596_ (
    .A(_18867_),
    .ZN(_18868_)
  );
  AND2_X1 _54597_ (
    .A1(_18866_),
    .A2(_18868_),
    .ZN(_18869_)
  );
  AND2_X1 _54598_ (
    .A1(instr_rdcycle),
    .A2(count_cycle[7]),
    .ZN(_18870_)
  );
  INV_X1 _54599_ (
    .A(_18870_),
    .ZN(_18871_)
  );
  AND2_X1 _54600_ (
    .A1(instr_rdcycleh),
    .A2(count_cycle[39]),
    .ZN(_18872_)
  );
  INV_X1 _54601_ (
    .A(_18872_),
    .ZN(_18873_)
  );
  AND2_X1 _54602_ (
    .A1(_18871_),
    .A2(_18873_),
    .ZN(_18874_)
  );
  AND2_X1 _54603_ (
    .A1(_18869_),
    .A2(_18874_),
    .ZN(_18875_)
  );
  INV_X1 _54604_ (
    .A(_18875_),
    .ZN(_18876_)
  );
  AND2_X1 _54605_ (
    .A1(_22271_),
    .A2(_18876_),
    .ZN(_18877_)
  );
  INV_X1 _54606_ (
    .A(_18877_),
    .ZN(_18878_)
  );
  AND2_X1 _54607_ (
    .A1(_18864_),
    .A2(_18878_),
    .ZN(_18879_)
  );
  AND2_X1 _54608_ (
    .A1(_18862_),
    .A2(_18879_),
    .ZN(_18880_)
  );
  AND2_X1 _54609_ (
    .A1(_18797_),
    .A2(_18803_),
    .ZN(_18881_)
  );
  INV_X1 _54610_ (
    .A(_18881_),
    .ZN(_18882_)
  );
  AND2_X1 _54611_ (
    .A1(reg_pc[7]),
    .A2(decoded_imm[7]),
    .ZN(_18883_)
  );
  INV_X1 _54612_ (
    .A(_18883_),
    .ZN(_18884_)
  );
  AND2_X1 _54613_ (
    .A1(_21097_),
    .A2(_22002_),
    .ZN(_18885_)
  );
  INV_X1 _54614_ (
    .A(_18885_),
    .ZN(_18886_)
  );
  AND2_X1 _54615_ (
    .A1(_18884_),
    .A2(_18886_),
    .ZN(_18887_)
  );
  INV_X1 _54616_ (
    .A(_18887_),
    .ZN(_18888_)
  );
  AND2_X1 _54617_ (
    .A1(_18881_),
    .A2(_18888_),
    .ZN(_18889_)
  );
  INV_X1 _54618_ (
    .A(_18889_),
    .ZN(_18890_)
  );
  AND2_X1 _54619_ (
    .A1(_18882_),
    .A2(_18887_),
    .ZN(_18891_)
  );
  INV_X1 _54620_ (
    .A(_18891_),
    .ZN(_18892_)
  );
  AND2_X1 _54621_ (
    .A1(_18890_),
    .A2(_18892_),
    .ZN(_18893_)
  );
  AND2_X1 _54622_ (
    .A1(_11090_),
    .A2(_18893_),
    .ZN(_18894_)
  );
  INV_X1 _54623_ (
    .A(_18894_),
    .ZN(_18895_)
  );
  AND2_X1 _54624_ (
    .A1(_18880_),
    .A2(_18895_),
    .ZN(_18896_)
  );
  INV_X1 _54625_ (
    .A(_18896_),
    .ZN(_18897_)
  );
  AND2_X1 _54626_ (
    .A1(resetn),
    .A2(_18897_),
    .ZN(_00005_[7])
  );
  AND2_X1 _54627_ (
    .A1(latched_is_lb),
    .A2(_18860_),
    .ZN(_18898_)
  );
  INV_X1 _54628_ (
    .A(_18898_),
    .ZN(_18899_)
  );
  AND2_X1 _54629_ (
    .A1(mem_rdata[8]),
    .A2(_12475_),
    .ZN(_18900_)
  );
  INV_X1 _54630_ (
    .A(_18900_),
    .ZN(_18901_)
  );
  AND2_X1 _54631_ (
    .A1(mem_rdata[24]),
    .A2(_12494_),
    .ZN(_18902_)
  );
  INV_X1 _54632_ (
    .A(_18902_),
    .ZN(_18903_)
  );
  AND2_X1 _54633_ (
    .A1(_18901_),
    .A2(_18903_),
    .ZN(_18904_)
  );
  INV_X1 _54634_ (
    .A(_18904_),
    .ZN(_18905_)
  );
  AND2_X1 _54635_ (
    .A1(_18476_),
    .A2(_18905_),
    .ZN(_18906_)
  );
  INV_X1 _54636_ (
    .A(_18906_),
    .ZN(_18907_)
  );
  AND2_X1 _54637_ (
    .A1(_18899_),
    .A2(_18907_),
    .ZN(_18908_)
  );
  INV_X1 _54638_ (
    .A(_18908_),
    .ZN(_18909_)
  );
  AND2_X1 _54639_ (
    .A1(_18479_),
    .A2(_18909_),
    .ZN(_18910_)
  );
  INV_X1 _54640_ (
    .A(_18910_),
    .ZN(_18911_)
  );
  AND2_X1 _54641_ (
    .A1(reg_op1[8]),
    .A2(_22282_),
    .ZN(_18912_)
  );
  INV_X1 _54642_ (
    .A(_18912_),
    .ZN(_18913_)
  );
  AND2_X1 _54643_ (
    .A1(count_instr[8]),
    .A2(instr_rdinstr),
    .ZN(_18914_)
  );
  INV_X1 _54644_ (
    .A(_18914_),
    .ZN(_18915_)
  );
  AND2_X1 _54645_ (
    .A1(instr_rdcycleh),
    .A2(count_cycle[40]),
    .ZN(_18916_)
  );
  INV_X1 _54646_ (
    .A(_18916_),
    .ZN(_18917_)
  );
  AND2_X1 _54647_ (
    .A1(_18915_),
    .A2(_18917_),
    .ZN(_18918_)
  );
  AND2_X1 _54648_ (
    .A1(count_instr[40]),
    .A2(instr_rdinstrh),
    .ZN(_18919_)
  );
  INV_X1 _54649_ (
    .A(_18919_),
    .ZN(_18920_)
  );
  AND2_X1 _54650_ (
    .A1(instr_rdcycle),
    .A2(count_cycle[8]),
    .ZN(_18921_)
  );
  INV_X1 _54651_ (
    .A(_18921_),
    .ZN(_18922_)
  );
  AND2_X1 _54652_ (
    .A1(_18920_),
    .A2(_18922_),
    .ZN(_18923_)
  );
  AND2_X1 _54653_ (
    .A1(_18918_),
    .A2(_18923_),
    .ZN(_18924_)
  );
  INV_X1 _54654_ (
    .A(_18924_),
    .ZN(_18925_)
  );
  AND2_X1 _54655_ (
    .A1(_22271_),
    .A2(_18925_),
    .ZN(_18926_)
  );
  INV_X1 _54656_ (
    .A(_18926_),
    .ZN(_18927_)
  );
  AND2_X1 _54657_ (
    .A1(_18913_),
    .A2(_18927_),
    .ZN(_18928_)
  );
  AND2_X1 _54658_ (
    .A1(_18911_),
    .A2(_18928_),
    .ZN(_18929_)
  );
  AND2_X1 _54659_ (
    .A1(reg_pc[8]),
    .A2(decoded_imm[8]),
    .ZN(_18930_)
  );
  INV_X1 _54660_ (
    .A(_18930_),
    .ZN(_18931_)
  );
  AND2_X1 _54661_ (
    .A1(_21096_),
    .A2(_22001_),
    .ZN(_18932_)
  );
  INV_X1 _54662_ (
    .A(_18932_),
    .ZN(_18933_)
  );
  AND2_X1 _54663_ (
    .A1(_18931_),
    .A2(_18933_),
    .ZN(_18934_)
  );
  INV_X1 _54664_ (
    .A(_18934_),
    .ZN(_18935_)
  );
  AND2_X1 _54665_ (
    .A1(_18882_),
    .A2(_18886_),
    .ZN(_18936_)
  );
  INV_X1 _54666_ (
    .A(_18936_),
    .ZN(_18937_)
  );
  AND2_X1 _54667_ (
    .A1(_18881_),
    .A2(_18884_),
    .ZN(_18938_)
  );
  INV_X1 _54668_ (
    .A(_18938_),
    .ZN(_18939_)
  );
  AND2_X1 _54669_ (
    .A1(_18884_),
    .A2(_18937_),
    .ZN(_18940_)
  );
  AND2_X1 _54670_ (
    .A1(_18886_),
    .A2(_18939_),
    .ZN(_18941_)
  );
  AND2_X1 _54671_ (
    .A1(_18935_),
    .A2(_18940_),
    .ZN(_18942_)
  );
  INV_X1 _54672_ (
    .A(_18942_),
    .ZN(_18943_)
  );
  AND2_X1 _54673_ (
    .A1(_18934_),
    .A2(_18941_),
    .ZN(_18944_)
  );
  INV_X1 _54674_ (
    .A(_18944_),
    .ZN(_18945_)
  );
  AND2_X1 _54675_ (
    .A1(_11090_),
    .A2(_18943_),
    .ZN(_18946_)
  );
  AND2_X1 _54676_ (
    .A1(_18945_),
    .A2(_18946_),
    .ZN(_18947_)
  );
  INV_X1 _54677_ (
    .A(_18947_),
    .ZN(_18948_)
  );
  AND2_X1 _54678_ (
    .A1(_18929_),
    .A2(_18948_),
    .ZN(_18949_)
  );
  INV_X1 _54679_ (
    .A(_18949_),
    .ZN(_18950_)
  );
  AND2_X1 _54680_ (
    .A1(resetn),
    .A2(_18950_),
    .ZN(_00005_[8])
  );
  AND2_X1 _54681_ (
    .A1(_18931_),
    .A2(_18945_),
    .ZN(_18951_)
  );
  INV_X1 _54682_ (
    .A(_18951_),
    .ZN(_18952_)
  );
  AND2_X1 _54683_ (
    .A1(reg_pc[9]),
    .A2(decoded_imm[9]),
    .ZN(_18953_)
  );
  INV_X1 _54684_ (
    .A(_18953_),
    .ZN(_18954_)
  );
  AND2_X1 _54685_ (
    .A1(_21095_),
    .A2(_22000_),
    .ZN(_18955_)
  );
  INV_X1 _54686_ (
    .A(_18955_),
    .ZN(_18956_)
  );
  AND2_X1 _54687_ (
    .A1(_18954_),
    .A2(_18956_),
    .ZN(_18957_)
  );
  INV_X1 _54688_ (
    .A(_18957_),
    .ZN(_18958_)
  );
  AND2_X1 _54689_ (
    .A1(_18952_),
    .A2(_18957_),
    .ZN(_18959_)
  );
  INV_X1 _54690_ (
    .A(_18959_),
    .ZN(_18960_)
  );
  AND2_X1 _54691_ (
    .A1(_18951_),
    .A2(_18958_),
    .ZN(_18961_)
  );
  INV_X1 _54692_ (
    .A(_18961_),
    .ZN(_18962_)
  );
  AND2_X1 _54693_ (
    .A1(_11090_),
    .A2(_18962_),
    .ZN(_18963_)
  );
  AND2_X1 _54694_ (
    .A1(_18960_),
    .A2(_18963_),
    .ZN(_18964_)
  );
  INV_X1 _54695_ (
    .A(_18964_),
    .ZN(_18965_)
  );
  AND2_X1 _54696_ (
    .A1(mem_rdata[9]),
    .A2(_12475_),
    .ZN(_18966_)
  );
  INV_X1 _54697_ (
    .A(_18966_),
    .ZN(_18967_)
  );
  AND2_X1 _54698_ (
    .A1(mem_rdata[25]),
    .A2(_12494_),
    .ZN(_18968_)
  );
  INV_X1 _54699_ (
    .A(_18968_),
    .ZN(_18969_)
  );
  AND2_X1 _54700_ (
    .A1(_18967_),
    .A2(_18969_),
    .ZN(_18970_)
  );
  INV_X1 _54701_ (
    .A(_18970_),
    .ZN(_18971_)
  );
  AND2_X1 _54702_ (
    .A1(_18476_),
    .A2(_18971_),
    .ZN(_18972_)
  );
  INV_X1 _54703_ (
    .A(_18972_),
    .ZN(_18973_)
  );
  AND2_X1 _54704_ (
    .A1(_18899_),
    .A2(_18973_),
    .ZN(_18974_)
  );
  INV_X1 _54705_ (
    .A(_18974_),
    .ZN(_18975_)
  );
  AND2_X1 _54706_ (
    .A1(_18479_),
    .A2(_18975_),
    .ZN(_18976_)
  );
  INV_X1 _54707_ (
    .A(_18976_),
    .ZN(_18977_)
  );
  AND2_X1 _54708_ (
    .A1(count_instr[41]),
    .A2(instr_rdinstrh),
    .ZN(_18978_)
  );
  INV_X1 _54709_ (
    .A(_18978_),
    .ZN(_18979_)
  );
  AND2_X1 _54710_ (
    .A1(count_instr[9]),
    .A2(instr_rdinstr),
    .ZN(_18980_)
  );
  INV_X1 _54711_ (
    .A(_18980_),
    .ZN(_18981_)
  );
  AND2_X1 _54712_ (
    .A1(_18979_),
    .A2(_18981_),
    .ZN(_18982_)
  );
  AND2_X1 _54713_ (
    .A1(instr_rdcycle),
    .A2(count_cycle[9]),
    .ZN(_18983_)
  );
  INV_X1 _54714_ (
    .A(_18983_),
    .ZN(_18984_)
  );
  AND2_X1 _54715_ (
    .A1(instr_rdcycleh),
    .A2(count_cycle[41]),
    .ZN(_18985_)
  );
  INV_X1 _54716_ (
    .A(_18985_),
    .ZN(_18986_)
  );
  AND2_X1 _54717_ (
    .A1(_18984_),
    .A2(_18986_),
    .ZN(_18987_)
  );
  AND2_X1 _54718_ (
    .A1(_18982_),
    .A2(_18987_),
    .ZN(_18988_)
  );
  INV_X1 _54719_ (
    .A(_18988_),
    .ZN(_18989_)
  );
  AND2_X1 _54720_ (
    .A1(_22271_),
    .A2(_18989_),
    .ZN(_18990_)
  );
  INV_X1 _54721_ (
    .A(_18990_),
    .ZN(_18991_)
  );
  AND2_X1 _54722_ (
    .A1(reg_op1[9]),
    .A2(_22282_),
    .ZN(_18992_)
  );
  INV_X1 _54723_ (
    .A(_18992_),
    .ZN(_18993_)
  );
  AND2_X1 _54724_ (
    .A1(_18991_),
    .A2(_18993_),
    .ZN(_18994_)
  );
  AND2_X1 _54725_ (
    .A1(_18977_),
    .A2(_18994_),
    .ZN(_18995_)
  );
  AND2_X1 _54726_ (
    .A1(_18965_),
    .A2(_18995_),
    .ZN(_18996_)
  );
  INV_X1 _54727_ (
    .A(_18996_),
    .ZN(_18997_)
  );
  AND2_X1 _54728_ (
    .A1(resetn),
    .A2(_18997_),
    .ZN(_00005_[9])
  );
  AND2_X1 _54729_ (
    .A1(mem_rdata[10]),
    .A2(_12475_),
    .ZN(_18998_)
  );
  INV_X1 _54730_ (
    .A(_18998_),
    .ZN(_18999_)
  );
  AND2_X1 _54731_ (
    .A1(mem_rdata[26]),
    .A2(_12494_),
    .ZN(_19000_)
  );
  INV_X1 _54732_ (
    .A(_19000_),
    .ZN(_19001_)
  );
  AND2_X1 _54733_ (
    .A1(_18999_),
    .A2(_19001_),
    .ZN(_19002_)
  );
  INV_X1 _54734_ (
    .A(_19002_),
    .ZN(_19003_)
  );
  AND2_X1 _54735_ (
    .A1(_18476_),
    .A2(_19003_),
    .ZN(_19004_)
  );
  INV_X1 _54736_ (
    .A(_19004_),
    .ZN(_19005_)
  );
  AND2_X1 _54737_ (
    .A1(_18899_),
    .A2(_19005_),
    .ZN(_19006_)
  );
  INV_X1 _54738_ (
    .A(_19006_),
    .ZN(_19007_)
  );
  AND2_X1 _54739_ (
    .A1(_18479_),
    .A2(_19007_),
    .ZN(_19008_)
  );
  INV_X1 _54740_ (
    .A(_19008_),
    .ZN(_19009_)
  );
  AND2_X1 _54741_ (
    .A1(reg_op1[10]),
    .A2(_22282_),
    .ZN(_19010_)
  );
  INV_X1 _54742_ (
    .A(_19010_),
    .ZN(_19011_)
  );
  AND2_X1 _54743_ (
    .A1(count_instr[10]),
    .A2(instr_rdinstr),
    .ZN(_19012_)
  );
  INV_X1 _54744_ (
    .A(_19012_),
    .ZN(_19013_)
  );
  AND2_X1 _54745_ (
    .A1(instr_rdcycleh),
    .A2(count_cycle[42]),
    .ZN(_19014_)
  );
  INV_X1 _54746_ (
    .A(_19014_),
    .ZN(_19015_)
  );
  AND2_X1 _54747_ (
    .A1(_19013_),
    .A2(_19015_),
    .ZN(_19016_)
  );
  AND2_X1 _54748_ (
    .A1(count_instr[42]),
    .A2(instr_rdinstrh),
    .ZN(_19017_)
  );
  INV_X1 _54749_ (
    .A(_19017_),
    .ZN(_19018_)
  );
  AND2_X1 _54750_ (
    .A1(instr_rdcycle),
    .A2(count_cycle[10]),
    .ZN(_19019_)
  );
  INV_X1 _54751_ (
    .A(_19019_),
    .ZN(_19020_)
  );
  AND2_X1 _54752_ (
    .A1(_19018_),
    .A2(_19020_),
    .ZN(_19021_)
  );
  AND2_X1 _54753_ (
    .A1(_19016_),
    .A2(_19021_),
    .ZN(_19022_)
  );
  INV_X1 _54754_ (
    .A(_19022_),
    .ZN(_19023_)
  );
  AND2_X1 _54755_ (
    .A1(_22271_),
    .A2(_19023_),
    .ZN(_19024_)
  );
  INV_X1 _54756_ (
    .A(_19024_),
    .ZN(_19025_)
  );
  AND2_X1 _54757_ (
    .A1(_19011_),
    .A2(_19025_),
    .ZN(_19026_)
  );
  AND2_X1 _54758_ (
    .A1(_19009_),
    .A2(_19026_),
    .ZN(_19027_)
  );
  AND2_X1 _54759_ (
    .A1(reg_pc[10]),
    .A2(decoded_imm[10]),
    .ZN(_19028_)
  );
  INV_X1 _54760_ (
    .A(_19028_),
    .ZN(_19029_)
  );
  AND2_X1 _54761_ (
    .A1(_21094_),
    .A2(_21999_),
    .ZN(_19030_)
  );
  INV_X1 _54762_ (
    .A(_19030_),
    .ZN(_19031_)
  );
  AND2_X1 _54763_ (
    .A1(_19029_),
    .A2(_19031_),
    .ZN(_19032_)
  );
  INV_X1 _54764_ (
    .A(_19032_),
    .ZN(_19033_)
  );
  AND2_X1 _54765_ (
    .A1(_18951_),
    .A2(_18954_),
    .ZN(_19034_)
  );
  INV_X1 _54766_ (
    .A(_19034_),
    .ZN(_19035_)
  );
  AND2_X1 _54767_ (
    .A1(_18952_),
    .A2(_18956_),
    .ZN(_19036_)
  );
  INV_X1 _54768_ (
    .A(_19036_),
    .ZN(_19037_)
  );
  AND2_X1 _54769_ (
    .A1(_18956_),
    .A2(_19035_),
    .ZN(_19038_)
  );
  AND2_X1 _54770_ (
    .A1(_18954_),
    .A2(_19037_),
    .ZN(_19039_)
  );
  AND2_X1 _54771_ (
    .A1(_19032_),
    .A2(_19038_),
    .ZN(_19040_)
  );
  INV_X1 _54772_ (
    .A(_19040_),
    .ZN(_19041_)
  );
  AND2_X1 _54773_ (
    .A1(_19033_),
    .A2(_19039_),
    .ZN(_19042_)
  );
  INV_X1 _54774_ (
    .A(_19042_),
    .ZN(_19043_)
  );
  AND2_X1 _54775_ (
    .A1(_11090_),
    .A2(_19041_),
    .ZN(_19044_)
  );
  AND2_X1 _54776_ (
    .A1(_19043_),
    .A2(_19044_),
    .ZN(_19045_)
  );
  INV_X1 _54777_ (
    .A(_19045_),
    .ZN(_19046_)
  );
  AND2_X1 _54778_ (
    .A1(_19027_),
    .A2(_19046_),
    .ZN(_19047_)
  );
  INV_X1 _54779_ (
    .A(_19047_),
    .ZN(_19048_)
  );
  AND2_X1 _54780_ (
    .A1(resetn),
    .A2(_19048_),
    .ZN(_00005_[10])
  );
  AND2_X1 _54781_ (
    .A1(mem_rdata[11]),
    .A2(_12475_),
    .ZN(_19049_)
  );
  INV_X1 _54782_ (
    .A(_19049_),
    .ZN(_19050_)
  );
  AND2_X1 _54783_ (
    .A1(mem_rdata[27]),
    .A2(_12494_),
    .ZN(_19051_)
  );
  INV_X1 _54784_ (
    .A(_19051_),
    .ZN(_19052_)
  );
  AND2_X1 _54785_ (
    .A1(_19050_),
    .A2(_19052_),
    .ZN(_19053_)
  );
  INV_X1 _54786_ (
    .A(_19053_),
    .ZN(_19054_)
  );
  AND2_X1 _54787_ (
    .A1(_18476_),
    .A2(_19054_),
    .ZN(_19055_)
  );
  INV_X1 _54788_ (
    .A(_19055_),
    .ZN(_19056_)
  );
  AND2_X1 _54789_ (
    .A1(_18899_),
    .A2(_19056_),
    .ZN(_19057_)
  );
  INV_X1 _54790_ (
    .A(_19057_),
    .ZN(_19058_)
  );
  AND2_X1 _54791_ (
    .A1(_18479_),
    .A2(_19058_),
    .ZN(_19059_)
  );
  INV_X1 _54792_ (
    .A(_19059_),
    .ZN(_19060_)
  );
  AND2_X1 _54793_ (
    .A1(count_instr[11]),
    .A2(instr_rdinstr),
    .ZN(_19061_)
  );
  INV_X1 _54794_ (
    .A(_19061_),
    .ZN(_19062_)
  );
  AND2_X1 _54795_ (
    .A1(instr_rdcycleh),
    .A2(count_cycle[43]),
    .ZN(_19063_)
  );
  INV_X1 _54796_ (
    .A(_19063_),
    .ZN(_19064_)
  );
  AND2_X1 _54797_ (
    .A1(_19062_),
    .A2(_19064_),
    .ZN(_19065_)
  );
  AND2_X1 _54798_ (
    .A1(count_instr[43]),
    .A2(instr_rdinstrh),
    .ZN(_19066_)
  );
  INV_X1 _54799_ (
    .A(_19066_),
    .ZN(_19067_)
  );
  AND2_X1 _54800_ (
    .A1(instr_rdcycle),
    .A2(count_cycle[11]),
    .ZN(_19068_)
  );
  INV_X1 _54801_ (
    .A(_19068_),
    .ZN(_19069_)
  );
  AND2_X1 _54802_ (
    .A1(_19067_),
    .A2(_19069_),
    .ZN(_19070_)
  );
  AND2_X1 _54803_ (
    .A1(_19065_),
    .A2(_19070_),
    .ZN(_19071_)
  );
  INV_X1 _54804_ (
    .A(_19071_),
    .ZN(_19072_)
  );
  AND2_X1 _54805_ (
    .A1(_22271_),
    .A2(_19072_),
    .ZN(_19073_)
  );
  INV_X1 _54806_ (
    .A(_19073_),
    .ZN(_19074_)
  );
  AND2_X1 _54807_ (
    .A1(reg_op1[11]),
    .A2(_22282_),
    .ZN(_19075_)
  );
  INV_X1 _54808_ (
    .A(_19075_),
    .ZN(_19076_)
  );
  AND2_X1 _54809_ (
    .A1(_19074_),
    .A2(_19076_),
    .ZN(_19077_)
  );
  AND2_X1 _54810_ (
    .A1(_19029_),
    .A2(_19041_),
    .ZN(_19078_)
  );
  INV_X1 _54811_ (
    .A(_19078_),
    .ZN(_19079_)
  );
  AND2_X1 _54812_ (
    .A1(reg_pc[11]),
    .A2(decoded_imm[11]),
    .ZN(_19080_)
  );
  INV_X1 _54813_ (
    .A(_19080_),
    .ZN(_19081_)
  );
  AND2_X1 _54814_ (
    .A1(_21093_),
    .A2(_21998_),
    .ZN(_19082_)
  );
  INV_X1 _54815_ (
    .A(_19082_),
    .ZN(_19083_)
  );
  AND2_X1 _54816_ (
    .A1(_19081_),
    .A2(_19083_),
    .ZN(_19084_)
  );
  INV_X1 _54817_ (
    .A(_19084_),
    .ZN(_19085_)
  );
  AND2_X1 _54818_ (
    .A1(_19079_),
    .A2(_19084_),
    .ZN(_19086_)
  );
  INV_X1 _54819_ (
    .A(_19086_),
    .ZN(_19087_)
  );
  AND2_X1 _54820_ (
    .A1(_19078_),
    .A2(_19085_),
    .ZN(_19088_)
  );
  INV_X1 _54821_ (
    .A(_19088_),
    .ZN(_19089_)
  );
  AND2_X1 _54822_ (
    .A1(_11090_),
    .A2(_19087_),
    .ZN(_19090_)
  );
  AND2_X1 _54823_ (
    .A1(_19089_),
    .A2(_19090_),
    .ZN(_19091_)
  );
  INV_X1 _54824_ (
    .A(_19091_),
    .ZN(_19092_)
  );
  AND2_X1 _54825_ (
    .A1(_19077_),
    .A2(_19092_),
    .ZN(_19093_)
  );
  AND2_X1 _54826_ (
    .A1(_19060_),
    .A2(_19093_),
    .ZN(_19094_)
  );
  INV_X1 _54827_ (
    .A(_19094_),
    .ZN(_19095_)
  );
  AND2_X1 _54828_ (
    .A1(resetn),
    .A2(_19095_),
    .ZN(_00005_[11])
  );
  AND2_X1 _54829_ (
    .A1(reg_pc[12]),
    .A2(decoded_imm[12]),
    .ZN(_19096_)
  );
  INV_X1 _54830_ (
    .A(_19096_),
    .ZN(_19097_)
  );
  AND2_X1 _54831_ (
    .A1(_21092_),
    .A2(_21997_),
    .ZN(_19098_)
  );
  INV_X1 _54832_ (
    .A(_19098_),
    .ZN(_19099_)
  );
  AND2_X1 _54833_ (
    .A1(_19097_),
    .A2(_19099_),
    .ZN(_19100_)
  );
  INV_X1 _54834_ (
    .A(_19100_),
    .ZN(_19101_)
  );
  AND2_X1 _54835_ (
    .A1(_19078_),
    .A2(_19081_),
    .ZN(_19102_)
  );
  INV_X1 _54836_ (
    .A(_19102_),
    .ZN(_19103_)
  );
  AND2_X1 _54837_ (
    .A1(_19079_),
    .A2(_19083_),
    .ZN(_19104_)
  );
  INV_X1 _54838_ (
    .A(_19104_),
    .ZN(_19105_)
  );
  AND2_X1 _54839_ (
    .A1(_19083_),
    .A2(_19103_),
    .ZN(_19106_)
  );
  AND2_X1 _54840_ (
    .A1(_19081_),
    .A2(_19105_),
    .ZN(_19107_)
  );
  AND2_X1 _54841_ (
    .A1(_19100_),
    .A2(_19106_),
    .ZN(_19108_)
  );
  INV_X1 _54842_ (
    .A(_19108_),
    .ZN(_19109_)
  );
  AND2_X1 _54843_ (
    .A1(_19101_),
    .A2(_19107_),
    .ZN(_19110_)
  );
  INV_X1 _54844_ (
    .A(_19110_),
    .ZN(_19111_)
  );
  AND2_X1 _54845_ (
    .A1(_19109_),
    .A2(_19111_),
    .ZN(_19112_)
  );
  AND2_X1 _54846_ (
    .A1(_11090_),
    .A2(_19112_),
    .ZN(_19113_)
  );
  INV_X1 _54847_ (
    .A(_19113_),
    .ZN(_19114_)
  );
  AND2_X1 _54848_ (
    .A1(mem_rdata[12]),
    .A2(_12475_),
    .ZN(_19115_)
  );
  INV_X1 _54849_ (
    .A(_19115_),
    .ZN(_19116_)
  );
  AND2_X1 _54850_ (
    .A1(mem_rdata[28]),
    .A2(_12494_),
    .ZN(_19117_)
  );
  INV_X1 _54851_ (
    .A(_19117_),
    .ZN(_19118_)
  );
  AND2_X1 _54852_ (
    .A1(_19116_),
    .A2(_19118_),
    .ZN(_19119_)
  );
  INV_X1 _54853_ (
    .A(_19119_),
    .ZN(_19120_)
  );
  AND2_X1 _54854_ (
    .A1(_18476_),
    .A2(_19120_),
    .ZN(_19121_)
  );
  INV_X1 _54855_ (
    .A(_19121_),
    .ZN(_19122_)
  );
  AND2_X1 _54856_ (
    .A1(_18899_),
    .A2(_19122_),
    .ZN(_19123_)
  );
  INV_X1 _54857_ (
    .A(_19123_),
    .ZN(_19124_)
  );
  AND2_X1 _54858_ (
    .A1(_18479_),
    .A2(_19124_),
    .ZN(_19125_)
  );
  INV_X1 _54859_ (
    .A(_19125_),
    .ZN(_19126_)
  );
  AND2_X1 _54860_ (
    .A1(reg_op1[12]),
    .A2(_22282_),
    .ZN(_19127_)
  );
  INV_X1 _54861_ (
    .A(_19127_),
    .ZN(_19128_)
  );
  AND2_X1 _54862_ (
    .A1(count_instr[12]),
    .A2(instr_rdinstr),
    .ZN(_19129_)
  );
  INV_X1 _54863_ (
    .A(_19129_),
    .ZN(_19130_)
  );
  AND2_X1 _54864_ (
    .A1(instr_rdcycleh),
    .A2(count_cycle[44]),
    .ZN(_19131_)
  );
  INV_X1 _54865_ (
    .A(_19131_),
    .ZN(_19132_)
  );
  AND2_X1 _54866_ (
    .A1(_19130_),
    .A2(_19132_),
    .ZN(_19133_)
  );
  AND2_X1 _54867_ (
    .A1(count_instr[44]),
    .A2(instr_rdinstrh),
    .ZN(_19134_)
  );
  INV_X1 _54868_ (
    .A(_19134_),
    .ZN(_19135_)
  );
  AND2_X1 _54869_ (
    .A1(instr_rdcycle),
    .A2(count_cycle[12]),
    .ZN(_19136_)
  );
  INV_X1 _54870_ (
    .A(_19136_),
    .ZN(_19137_)
  );
  AND2_X1 _54871_ (
    .A1(_19135_),
    .A2(_19137_),
    .ZN(_19138_)
  );
  AND2_X1 _54872_ (
    .A1(_19133_),
    .A2(_19138_),
    .ZN(_19139_)
  );
  INV_X1 _54873_ (
    .A(_19139_),
    .ZN(_19140_)
  );
  AND2_X1 _54874_ (
    .A1(_22271_),
    .A2(_19140_),
    .ZN(_19141_)
  );
  INV_X1 _54875_ (
    .A(_19141_),
    .ZN(_19142_)
  );
  AND2_X1 _54876_ (
    .A1(_19128_),
    .A2(_19142_),
    .ZN(_19143_)
  );
  AND2_X1 _54877_ (
    .A1(_19126_),
    .A2(_19143_),
    .ZN(_19144_)
  );
  AND2_X1 _54878_ (
    .A1(_19114_),
    .A2(_19144_),
    .ZN(_19145_)
  );
  INV_X1 _54879_ (
    .A(_19145_),
    .ZN(_19146_)
  );
  AND2_X1 _54880_ (
    .A1(resetn),
    .A2(_19146_),
    .ZN(_00005_[12])
  );
  AND2_X1 _54881_ (
    .A1(mem_rdata[13]),
    .A2(_12475_),
    .ZN(_19147_)
  );
  INV_X1 _54882_ (
    .A(_19147_),
    .ZN(_19148_)
  );
  AND2_X1 _54883_ (
    .A1(mem_rdata[29]),
    .A2(_12494_),
    .ZN(_19149_)
  );
  INV_X1 _54884_ (
    .A(_19149_),
    .ZN(_19150_)
  );
  AND2_X1 _54885_ (
    .A1(_19148_),
    .A2(_19150_),
    .ZN(_19151_)
  );
  INV_X1 _54886_ (
    .A(_19151_),
    .ZN(_19152_)
  );
  AND2_X1 _54887_ (
    .A1(_18476_),
    .A2(_19152_),
    .ZN(_19153_)
  );
  INV_X1 _54888_ (
    .A(_19153_),
    .ZN(_19154_)
  );
  AND2_X1 _54889_ (
    .A1(_18899_),
    .A2(_19154_),
    .ZN(_19155_)
  );
  INV_X1 _54890_ (
    .A(_19155_),
    .ZN(_19156_)
  );
  AND2_X1 _54891_ (
    .A1(_18479_),
    .A2(_19156_),
    .ZN(_19157_)
  );
  INV_X1 _54892_ (
    .A(_19157_),
    .ZN(_19158_)
  );
  AND2_X1 _54893_ (
    .A1(reg_op1[13]),
    .A2(_22282_),
    .ZN(_19159_)
  );
  INV_X1 _54894_ (
    .A(_19159_),
    .ZN(_19160_)
  );
  AND2_X1 _54895_ (
    .A1(count_instr[13]),
    .A2(instr_rdinstr),
    .ZN(_19161_)
  );
  INV_X1 _54896_ (
    .A(_19161_),
    .ZN(_19162_)
  );
  AND2_X1 _54897_ (
    .A1(instr_rdcycleh),
    .A2(count_cycle[45]),
    .ZN(_19163_)
  );
  INV_X1 _54898_ (
    .A(_19163_),
    .ZN(_19164_)
  );
  AND2_X1 _54899_ (
    .A1(_19162_),
    .A2(_19164_),
    .ZN(_19165_)
  );
  AND2_X1 _54900_ (
    .A1(count_instr[45]),
    .A2(instr_rdinstrh),
    .ZN(_19166_)
  );
  INV_X1 _54901_ (
    .A(_19166_),
    .ZN(_19167_)
  );
  AND2_X1 _54902_ (
    .A1(instr_rdcycle),
    .A2(count_cycle[13]),
    .ZN(_19168_)
  );
  INV_X1 _54903_ (
    .A(_19168_),
    .ZN(_19169_)
  );
  AND2_X1 _54904_ (
    .A1(_19167_),
    .A2(_19169_),
    .ZN(_19170_)
  );
  AND2_X1 _54905_ (
    .A1(_19165_),
    .A2(_19170_),
    .ZN(_19171_)
  );
  INV_X1 _54906_ (
    .A(_19171_),
    .ZN(_19172_)
  );
  AND2_X1 _54907_ (
    .A1(_22271_),
    .A2(_19172_),
    .ZN(_19173_)
  );
  INV_X1 _54908_ (
    .A(_19173_),
    .ZN(_19174_)
  );
  AND2_X1 _54909_ (
    .A1(_19160_),
    .A2(_19174_),
    .ZN(_19175_)
  );
  AND2_X1 _54910_ (
    .A1(_19158_),
    .A2(_19175_),
    .ZN(_19176_)
  );
  AND2_X1 _54911_ (
    .A1(_19097_),
    .A2(_19109_),
    .ZN(_19177_)
  );
  INV_X1 _54912_ (
    .A(_19177_),
    .ZN(_19178_)
  );
  AND2_X1 _54913_ (
    .A1(reg_pc[13]),
    .A2(decoded_imm[13]),
    .ZN(_19179_)
  );
  INV_X1 _54914_ (
    .A(_19179_),
    .ZN(_19180_)
  );
  AND2_X1 _54915_ (
    .A1(_21091_),
    .A2(_21996_),
    .ZN(_19181_)
  );
  INV_X1 _54916_ (
    .A(_19181_),
    .ZN(_19182_)
  );
  AND2_X1 _54917_ (
    .A1(_19180_),
    .A2(_19182_),
    .ZN(_19183_)
  );
  INV_X1 _54918_ (
    .A(_19183_),
    .ZN(_19184_)
  );
  AND2_X1 _54919_ (
    .A1(_19178_),
    .A2(_19183_),
    .ZN(_19185_)
  );
  INV_X1 _54920_ (
    .A(_19185_),
    .ZN(_19186_)
  );
  AND2_X1 _54921_ (
    .A1(_19177_),
    .A2(_19184_),
    .ZN(_19187_)
  );
  INV_X1 _54922_ (
    .A(_19187_),
    .ZN(_19188_)
  );
  AND2_X1 _54923_ (
    .A1(_19186_),
    .A2(_19188_),
    .ZN(_19189_)
  );
  AND2_X1 _54924_ (
    .A1(_11090_),
    .A2(_19189_),
    .ZN(_19190_)
  );
  INV_X1 _54925_ (
    .A(_19190_),
    .ZN(_19191_)
  );
  AND2_X1 _54926_ (
    .A1(_19176_),
    .A2(_19191_),
    .ZN(_19192_)
  );
  INV_X1 _54927_ (
    .A(_19192_),
    .ZN(_19193_)
  );
  AND2_X1 _54928_ (
    .A1(resetn),
    .A2(_19193_),
    .ZN(_00005_[13])
  );
  AND2_X1 _54929_ (
    .A1(reg_pc[14]),
    .A2(decoded_imm[14]),
    .ZN(_19194_)
  );
  INV_X1 _54930_ (
    .A(_19194_),
    .ZN(_19195_)
  );
  AND2_X1 _54931_ (
    .A1(_21090_),
    .A2(_21995_),
    .ZN(_19196_)
  );
  INV_X1 _54932_ (
    .A(_19196_),
    .ZN(_19197_)
  );
  AND2_X1 _54933_ (
    .A1(_19195_),
    .A2(_19197_),
    .ZN(_19198_)
  );
  INV_X1 _54934_ (
    .A(_19198_),
    .ZN(_19199_)
  );
  AND2_X1 _54935_ (
    .A1(_19177_),
    .A2(_19180_),
    .ZN(_19200_)
  );
  INV_X1 _54936_ (
    .A(_19200_),
    .ZN(_19201_)
  );
  AND2_X1 _54937_ (
    .A1(_19178_),
    .A2(_19182_),
    .ZN(_19202_)
  );
  INV_X1 _54938_ (
    .A(_19202_),
    .ZN(_19203_)
  );
  AND2_X1 _54939_ (
    .A1(_19182_),
    .A2(_19201_),
    .ZN(_19204_)
  );
  AND2_X1 _54940_ (
    .A1(_19180_),
    .A2(_19203_),
    .ZN(_19205_)
  );
  AND2_X1 _54941_ (
    .A1(_19198_),
    .A2(_19204_),
    .ZN(_19206_)
  );
  INV_X1 _54942_ (
    .A(_19206_),
    .ZN(_19207_)
  );
  AND2_X1 _54943_ (
    .A1(_19199_),
    .A2(_19205_),
    .ZN(_19208_)
  );
  INV_X1 _54944_ (
    .A(_19208_),
    .ZN(_19209_)
  );
  AND2_X1 _54945_ (
    .A1(_11090_),
    .A2(_19209_),
    .ZN(_19210_)
  );
  AND2_X1 _54946_ (
    .A1(_19207_),
    .A2(_19210_),
    .ZN(_19211_)
  );
  INV_X1 _54947_ (
    .A(_19211_),
    .ZN(_19212_)
  );
  AND2_X1 _54948_ (
    .A1(mem_rdata[14]),
    .A2(_12475_),
    .ZN(_19213_)
  );
  INV_X1 _54949_ (
    .A(_19213_),
    .ZN(_19214_)
  );
  AND2_X1 _54950_ (
    .A1(mem_rdata[30]),
    .A2(_12494_),
    .ZN(_19215_)
  );
  INV_X1 _54951_ (
    .A(_19215_),
    .ZN(_19216_)
  );
  AND2_X1 _54952_ (
    .A1(_19214_),
    .A2(_19216_),
    .ZN(_19217_)
  );
  INV_X1 _54953_ (
    .A(_19217_),
    .ZN(_19218_)
  );
  AND2_X1 _54954_ (
    .A1(_18476_),
    .A2(_19218_),
    .ZN(_19219_)
  );
  INV_X1 _54955_ (
    .A(_19219_),
    .ZN(_19220_)
  );
  AND2_X1 _54956_ (
    .A1(_18899_),
    .A2(_19220_),
    .ZN(_19221_)
  );
  INV_X1 _54957_ (
    .A(_19221_),
    .ZN(_19222_)
  );
  AND2_X1 _54958_ (
    .A1(_18479_),
    .A2(_19222_),
    .ZN(_19223_)
  );
  INV_X1 _54959_ (
    .A(_19223_),
    .ZN(_19224_)
  );
  AND2_X1 _54960_ (
    .A1(reg_op1[14]),
    .A2(_22282_),
    .ZN(_19225_)
  );
  INV_X1 _54961_ (
    .A(_19225_),
    .ZN(_19226_)
  );
  AND2_X1 _54962_ (
    .A1(count_instr[14]),
    .A2(instr_rdinstr),
    .ZN(_19227_)
  );
  INV_X1 _54963_ (
    .A(_19227_),
    .ZN(_19228_)
  );
  AND2_X1 _54964_ (
    .A1(instr_rdcycleh),
    .A2(count_cycle[46]),
    .ZN(_19229_)
  );
  INV_X1 _54965_ (
    .A(_19229_),
    .ZN(_19230_)
  );
  AND2_X1 _54966_ (
    .A1(_19228_),
    .A2(_19230_),
    .ZN(_19231_)
  );
  AND2_X1 _54967_ (
    .A1(count_instr[46]),
    .A2(instr_rdinstrh),
    .ZN(_19232_)
  );
  INV_X1 _54968_ (
    .A(_19232_),
    .ZN(_19233_)
  );
  AND2_X1 _54969_ (
    .A1(instr_rdcycle),
    .A2(count_cycle[14]),
    .ZN(_19234_)
  );
  INV_X1 _54970_ (
    .A(_19234_),
    .ZN(_19235_)
  );
  AND2_X1 _54971_ (
    .A1(_19233_),
    .A2(_19235_),
    .ZN(_19236_)
  );
  AND2_X1 _54972_ (
    .A1(_19231_),
    .A2(_19236_),
    .ZN(_19237_)
  );
  INV_X1 _54973_ (
    .A(_19237_),
    .ZN(_19238_)
  );
  AND2_X1 _54974_ (
    .A1(_22271_),
    .A2(_19238_),
    .ZN(_19239_)
  );
  INV_X1 _54975_ (
    .A(_19239_),
    .ZN(_19240_)
  );
  AND2_X1 _54976_ (
    .A1(_19226_),
    .A2(_19240_),
    .ZN(_19241_)
  );
  AND2_X1 _54977_ (
    .A1(_19224_),
    .A2(_19241_),
    .ZN(_19242_)
  );
  AND2_X1 _54978_ (
    .A1(_19212_),
    .A2(_19242_),
    .ZN(_19243_)
  );
  INV_X1 _54979_ (
    .A(_19243_),
    .ZN(_19244_)
  );
  AND2_X1 _54980_ (
    .A1(resetn),
    .A2(_19244_),
    .ZN(_00005_[14])
  );
  AND2_X1 _54981_ (
    .A1(_19195_),
    .A2(_19207_),
    .ZN(_19245_)
  );
  INV_X1 _54982_ (
    .A(_19245_),
    .ZN(_19246_)
  );
  AND2_X1 _54983_ (
    .A1(reg_pc[15]),
    .A2(decoded_imm[15]),
    .ZN(_19247_)
  );
  INV_X1 _54984_ (
    .A(_19247_),
    .ZN(_19248_)
  );
  AND2_X1 _54985_ (
    .A1(_21089_),
    .A2(_21994_),
    .ZN(_19249_)
  );
  INV_X1 _54986_ (
    .A(_19249_),
    .ZN(_19250_)
  );
  AND2_X1 _54987_ (
    .A1(_19248_),
    .A2(_19250_),
    .ZN(_19251_)
  );
  INV_X1 _54988_ (
    .A(_19251_),
    .ZN(_19252_)
  );
  AND2_X1 _54989_ (
    .A1(_19246_),
    .A2(_19251_),
    .ZN(_19253_)
  );
  INV_X1 _54990_ (
    .A(_19253_),
    .ZN(_19254_)
  );
  AND2_X1 _54991_ (
    .A1(_19245_),
    .A2(_19252_),
    .ZN(_19255_)
  );
  INV_X1 _54992_ (
    .A(_19255_),
    .ZN(_19256_)
  );
  AND2_X1 _54993_ (
    .A1(_11090_),
    .A2(_19256_),
    .ZN(_19257_)
  );
  AND2_X1 _54994_ (
    .A1(_19254_),
    .A2(_19257_),
    .ZN(_19258_)
  );
  INV_X1 _54995_ (
    .A(_19258_),
    .ZN(_19259_)
  );
  AND2_X1 _54996_ (
    .A1(mem_rdata[15]),
    .A2(_12475_),
    .ZN(_19260_)
  );
  INV_X1 _54997_ (
    .A(_19260_),
    .ZN(_19261_)
  );
  AND2_X1 _54998_ (
    .A1(mem_rdata[31]),
    .A2(_12494_),
    .ZN(_19262_)
  );
  INV_X1 _54999_ (
    .A(_19262_),
    .ZN(_19263_)
  );
  AND2_X1 _55000_ (
    .A1(_19261_),
    .A2(_19263_),
    .ZN(_19264_)
  );
  INV_X1 _55001_ (
    .A(_19264_),
    .ZN(_19265_)
  );
  AND2_X1 _55002_ (
    .A1(_18476_),
    .A2(_19265_),
    .ZN(_19266_)
  );
  INV_X1 _55003_ (
    .A(_19266_),
    .ZN(_19267_)
  );
  AND2_X1 _55004_ (
    .A1(_18899_),
    .A2(_19267_),
    .ZN(_19268_)
  );
  INV_X1 _55005_ (
    .A(_19268_),
    .ZN(_19269_)
  );
  AND2_X1 _55006_ (
    .A1(_18479_),
    .A2(_19269_),
    .ZN(_19270_)
  );
  INV_X1 _55007_ (
    .A(_19270_),
    .ZN(_19271_)
  );
  AND2_X1 _55008_ (
    .A1(instr_rdcycleh),
    .A2(count_cycle[47]),
    .ZN(_19272_)
  );
  INV_X1 _55009_ (
    .A(_19272_),
    .ZN(_19273_)
  );
  AND2_X1 _55010_ (
    .A1(count_instr[15]),
    .A2(instr_rdinstr),
    .ZN(_19274_)
  );
  INV_X1 _55011_ (
    .A(_19274_),
    .ZN(_19275_)
  );
  AND2_X1 _55012_ (
    .A1(_19273_),
    .A2(_19275_),
    .ZN(_19276_)
  );
  AND2_X1 _55013_ (
    .A1(instr_rdcycle),
    .A2(count_cycle[15]),
    .ZN(_19277_)
  );
  INV_X1 _55014_ (
    .A(_19277_),
    .ZN(_19278_)
  );
  AND2_X1 _55015_ (
    .A1(count_instr[47]),
    .A2(instr_rdinstrh),
    .ZN(_19279_)
  );
  INV_X1 _55016_ (
    .A(_19279_),
    .ZN(_19280_)
  );
  AND2_X1 _55017_ (
    .A1(_19278_),
    .A2(_19280_),
    .ZN(_19281_)
  );
  AND2_X1 _55018_ (
    .A1(_19276_),
    .A2(_19281_),
    .ZN(_19282_)
  );
  INV_X1 _55019_ (
    .A(_19282_),
    .ZN(_19283_)
  );
  AND2_X1 _55020_ (
    .A1(_22271_),
    .A2(_19283_),
    .ZN(_19284_)
  );
  INV_X1 _55021_ (
    .A(_19284_),
    .ZN(_19285_)
  );
  AND2_X1 _55022_ (
    .A1(reg_op1[15]),
    .A2(_22282_),
    .ZN(_19286_)
  );
  INV_X1 _55023_ (
    .A(_19286_),
    .ZN(_19287_)
  );
  AND2_X1 _55024_ (
    .A1(_19285_),
    .A2(_19287_),
    .ZN(_19288_)
  );
  AND2_X1 _55025_ (
    .A1(_19271_),
    .A2(_19288_),
    .ZN(_19289_)
  );
  AND2_X1 _55026_ (
    .A1(_19259_),
    .A2(_19289_),
    .ZN(_19290_)
  );
  INV_X1 _55027_ (
    .A(_19290_),
    .ZN(_19291_)
  );
  AND2_X1 _55028_ (
    .A1(resetn),
    .A2(_19291_),
    .ZN(_00005_[15])
  );
  AND2_X1 _55029_ (
    .A1(reg_pc[16]),
    .A2(decoded_imm[16]),
    .ZN(_19292_)
  );
  INV_X1 _55030_ (
    .A(_19292_),
    .ZN(_19293_)
  );
  AND2_X1 _55031_ (
    .A1(_21088_),
    .A2(_21993_),
    .ZN(_19294_)
  );
  INV_X1 _55032_ (
    .A(_19294_),
    .ZN(_19295_)
  );
  AND2_X1 _55033_ (
    .A1(_19293_),
    .A2(_19295_),
    .ZN(_19296_)
  );
  INV_X1 _55034_ (
    .A(_19296_),
    .ZN(_19297_)
  );
  AND2_X1 _55035_ (
    .A1(_19245_),
    .A2(_19248_),
    .ZN(_19298_)
  );
  INV_X1 _55036_ (
    .A(_19298_),
    .ZN(_19299_)
  );
  AND2_X1 _55037_ (
    .A1(_19246_),
    .A2(_19250_),
    .ZN(_19300_)
  );
  INV_X1 _55038_ (
    .A(_19300_),
    .ZN(_19301_)
  );
  AND2_X1 _55039_ (
    .A1(_19250_),
    .A2(_19299_),
    .ZN(_19302_)
  );
  AND2_X1 _55040_ (
    .A1(_19248_),
    .A2(_19301_),
    .ZN(_19303_)
  );
  AND2_X1 _55041_ (
    .A1(_19296_),
    .A2(_19302_),
    .ZN(_19304_)
  );
  INV_X1 _55042_ (
    .A(_19304_),
    .ZN(_19305_)
  );
  AND2_X1 _55043_ (
    .A1(_19297_),
    .A2(_19303_),
    .ZN(_19306_)
  );
  INV_X1 _55044_ (
    .A(_19306_),
    .ZN(_19307_)
  );
  AND2_X1 _55045_ (
    .A1(_11090_),
    .A2(_19307_),
    .ZN(_19308_)
  );
  AND2_X1 _55046_ (
    .A1(_19305_),
    .A2(_19308_),
    .ZN(_19309_)
  );
  INV_X1 _55047_ (
    .A(_19309_),
    .ZN(_19310_)
  );
  AND2_X1 _55048_ (
    .A1(latched_is_lh),
    .A2(_19265_),
    .ZN(_19311_)
  );
  INV_X1 _55049_ (
    .A(_19311_),
    .ZN(_19312_)
  );
  AND2_X1 _55050_ (
    .A1(_18899_),
    .A2(_19312_),
    .ZN(_19313_)
  );
  AND2_X1 _55051_ (
    .A1(latched_is_lu),
    .A2(mem_rdata[16]),
    .ZN(_19314_)
  );
  AND2_X1 _55052_ (
    .A1(_12194_),
    .A2(_19314_),
    .ZN(_19315_)
  );
  INV_X1 _55053_ (
    .A(_19315_),
    .ZN(_19316_)
  );
  AND2_X1 _55054_ (
    .A1(_19313_),
    .A2(_19316_),
    .ZN(_19317_)
  );
  INV_X1 _55055_ (
    .A(_19317_),
    .ZN(_19318_)
  );
  AND2_X1 _55056_ (
    .A1(_18479_),
    .A2(_19318_),
    .ZN(_19319_)
  );
  INV_X1 _55057_ (
    .A(_19319_),
    .ZN(_19320_)
  );
  AND2_X1 _55058_ (
    .A1(count_instr[48]),
    .A2(instr_rdinstrh),
    .ZN(_19321_)
  );
  INV_X1 _55059_ (
    .A(_19321_),
    .ZN(_19322_)
  );
  AND2_X1 _55060_ (
    .A1(count_instr[16]),
    .A2(instr_rdinstr),
    .ZN(_19323_)
  );
  INV_X1 _55061_ (
    .A(_19323_),
    .ZN(_19324_)
  );
  AND2_X1 _55062_ (
    .A1(_19322_),
    .A2(_19324_),
    .ZN(_19325_)
  );
  AND2_X1 _55063_ (
    .A1(instr_rdcycle),
    .A2(count_cycle[16]),
    .ZN(_19326_)
  );
  INV_X1 _55064_ (
    .A(_19326_),
    .ZN(_19327_)
  );
  AND2_X1 _55065_ (
    .A1(instr_rdcycleh),
    .A2(count_cycle[48]),
    .ZN(_19328_)
  );
  INV_X1 _55066_ (
    .A(_19328_),
    .ZN(_19329_)
  );
  AND2_X1 _55067_ (
    .A1(_19327_),
    .A2(_19329_),
    .ZN(_19330_)
  );
  AND2_X1 _55068_ (
    .A1(_19325_),
    .A2(_19330_),
    .ZN(_19331_)
  );
  INV_X1 _55069_ (
    .A(_19331_),
    .ZN(_19332_)
  );
  AND2_X1 _55070_ (
    .A1(_22271_),
    .A2(_19332_),
    .ZN(_19333_)
  );
  INV_X1 _55071_ (
    .A(_19333_),
    .ZN(_19334_)
  );
  AND2_X1 _55072_ (
    .A1(reg_op1[16]),
    .A2(_22282_),
    .ZN(_19335_)
  );
  INV_X1 _55073_ (
    .A(_19335_),
    .ZN(_19336_)
  );
  AND2_X1 _55074_ (
    .A1(_19334_),
    .A2(_19336_),
    .ZN(_19337_)
  );
  AND2_X1 _55075_ (
    .A1(_19320_),
    .A2(_19337_),
    .ZN(_19338_)
  );
  AND2_X1 _55076_ (
    .A1(_19310_),
    .A2(_19338_),
    .ZN(_19339_)
  );
  INV_X1 _55077_ (
    .A(_19339_),
    .ZN(_19340_)
  );
  AND2_X1 _55078_ (
    .A1(resetn),
    .A2(_19340_),
    .ZN(_00005_[16])
  );
  AND2_X1 _55079_ (
    .A1(latched_is_lu),
    .A2(mem_rdata[17]),
    .ZN(_19341_)
  );
  AND2_X1 _55080_ (
    .A1(_12194_),
    .A2(_19341_),
    .ZN(_19342_)
  );
  INV_X1 _55081_ (
    .A(_19342_),
    .ZN(_19343_)
  );
  AND2_X1 _55082_ (
    .A1(_19313_),
    .A2(_19343_),
    .ZN(_19344_)
  );
  INV_X1 _55083_ (
    .A(_19344_),
    .ZN(_19345_)
  );
  AND2_X1 _55084_ (
    .A1(_18479_),
    .A2(_19345_),
    .ZN(_19346_)
  );
  INV_X1 _55085_ (
    .A(_19346_),
    .ZN(_19347_)
  );
  AND2_X1 _55086_ (
    .A1(count_instr[17]),
    .A2(instr_rdinstr),
    .ZN(_19348_)
  );
  INV_X1 _55087_ (
    .A(_19348_),
    .ZN(_19349_)
  );
  AND2_X1 _55088_ (
    .A1(instr_rdcycleh),
    .A2(count_cycle[49]),
    .ZN(_19350_)
  );
  INV_X1 _55089_ (
    .A(_19350_),
    .ZN(_19351_)
  );
  AND2_X1 _55090_ (
    .A1(_19349_),
    .A2(_19351_),
    .ZN(_19352_)
  );
  AND2_X1 _55091_ (
    .A1(instr_rdcycle),
    .A2(count_cycle[17]),
    .ZN(_19353_)
  );
  INV_X1 _55092_ (
    .A(_19353_),
    .ZN(_19354_)
  );
  AND2_X1 _55093_ (
    .A1(count_instr[49]),
    .A2(instr_rdinstrh),
    .ZN(_19355_)
  );
  INV_X1 _55094_ (
    .A(_19355_),
    .ZN(_19356_)
  );
  AND2_X1 _55095_ (
    .A1(_19354_),
    .A2(_19356_),
    .ZN(_19357_)
  );
  AND2_X1 _55096_ (
    .A1(_19352_),
    .A2(_19357_),
    .ZN(_19358_)
  );
  INV_X1 _55097_ (
    .A(_19358_),
    .ZN(_19359_)
  );
  AND2_X1 _55098_ (
    .A1(_22271_),
    .A2(_19359_),
    .ZN(_19360_)
  );
  INV_X1 _55099_ (
    .A(_19360_),
    .ZN(_19361_)
  );
  AND2_X1 _55100_ (
    .A1(reg_op1[17]),
    .A2(_22282_),
    .ZN(_19362_)
  );
  INV_X1 _55101_ (
    .A(_19362_),
    .ZN(_19363_)
  );
  AND2_X1 _55102_ (
    .A1(_19361_),
    .A2(_19363_),
    .ZN(_19364_)
  );
  AND2_X1 _55103_ (
    .A1(_19347_),
    .A2(_19364_),
    .ZN(_19365_)
  );
  AND2_X1 _55104_ (
    .A1(_19293_),
    .A2(_19305_),
    .ZN(_19366_)
  );
  INV_X1 _55105_ (
    .A(_19366_),
    .ZN(_19367_)
  );
  AND2_X1 _55106_ (
    .A1(reg_pc[17]),
    .A2(decoded_imm[17]),
    .ZN(_19368_)
  );
  INV_X1 _55107_ (
    .A(_19368_),
    .ZN(_19369_)
  );
  AND2_X1 _55108_ (
    .A1(_21087_),
    .A2(_21992_),
    .ZN(_19370_)
  );
  INV_X1 _55109_ (
    .A(_19370_),
    .ZN(_19371_)
  );
  AND2_X1 _55110_ (
    .A1(_19369_),
    .A2(_19371_),
    .ZN(_19372_)
  );
  INV_X1 _55111_ (
    .A(_19372_),
    .ZN(_19373_)
  );
  AND2_X1 _55112_ (
    .A1(_19367_),
    .A2(_19372_),
    .ZN(_19374_)
  );
  INV_X1 _55113_ (
    .A(_19374_),
    .ZN(_19375_)
  );
  AND2_X1 _55114_ (
    .A1(_19366_),
    .A2(_19373_),
    .ZN(_19376_)
  );
  INV_X1 _55115_ (
    .A(_19376_),
    .ZN(_19377_)
  );
  AND2_X1 _55116_ (
    .A1(_11090_),
    .A2(_19377_),
    .ZN(_19378_)
  );
  AND2_X1 _55117_ (
    .A1(_19375_),
    .A2(_19378_),
    .ZN(_19379_)
  );
  INV_X1 _55118_ (
    .A(_19379_),
    .ZN(_19380_)
  );
  AND2_X1 _55119_ (
    .A1(_19365_),
    .A2(_19380_),
    .ZN(_19381_)
  );
  INV_X1 _55120_ (
    .A(_19381_),
    .ZN(_19382_)
  );
  AND2_X1 _55121_ (
    .A1(resetn),
    .A2(_19382_),
    .ZN(_00005_[17])
  );
  AND2_X1 _55122_ (
    .A1(reg_pc[18]),
    .A2(decoded_imm[18]),
    .ZN(_19383_)
  );
  INV_X1 _55123_ (
    .A(_19383_),
    .ZN(_19384_)
  );
  AND2_X1 _55124_ (
    .A1(_21086_),
    .A2(_21991_),
    .ZN(_19385_)
  );
  INV_X1 _55125_ (
    .A(_19385_),
    .ZN(_19386_)
  );
  AND2_X1 _55126_ (
    .A1(_19384_),
    .A2(_19386_),
    .ZN(_19387_)
  );
  INV_X1 _55127_ (
    .A(_19387_),
    .ZN(_19388_)
  );
  AND2_X1 _55128_ (
    .A1(_19366_),
    .A2(_19369_),
    .ZN(_19389_)
  );
  INV_X1 _55129_ (
    .A(_19389_),
    .ZN(_19390_)
  );
  AND2_X1 _55130_ (
    .A1(_19367_),
    .A2(_19371_),
    .ZN(_19391_)
  );
  INV_X1 _55131_ (
    .A(_19391_),
    .ZN(_19392_)
  );
  AND2_X1 _55132_ (
    .A1(_19371_),
    .A2(_19390_),
    .ZN(_19393_)
  );
  AND2_X1 _55133_ (
    .A1(_19369_),
    .A2(_19392_),
    .ZN(_19394_)
  );
  AND2_X1 _55134_ (
    .A1(_19387_),
    .A2(_19393_),
    .ZN(_19395_)
  );
  INV_X1 _55135_ (
    .A(_19395_),
    .ZN(_19396_)
  );
  AND2_X1 _55136_ (
    .A1(_19388_),
    .A2(_19394_),
    .ZN(_19397_)
  );
  INV_X1 _55137_ (
    .A(_19397_),
    .ZN(_19398_)
  );
  AND2_X1 _55138_ (
    .A1(_19396_),
    .A2(_19398_),
    .ZN(_19399_)
  );
  AND2_X1 _55139_ (
    .A1(_11090_),
    .A2(_19399_),
    .ZN(_19400_)
  );
  INV_X1 _55140_ (
    .A(_19400_),
    .ZN(_19401_)
  );
  AND2_X1 _55141_ (
    .A1(latched_is_lu),
    .A2(mem_rdata[18]),
    .ZN(_19402_)
  );
  AND2_X1 _55142_ (
    .A1(_12194_),
    .A2(_19402_),
    .ZN(_19403_)
  );
  INV_X1 _55143_ (
    .A(_19403_),
    .ZN(_19404_)
  );
  AND2_X1 _55144_ (
    .A1(_19313_),
    .A2(_19404_),
    .ZN(_19405_)
  );
  INV_X1 _55145_ (
    .A(_19405_),
    .ZN(_19406_)
  );
  AND2_X1 _55146_ (
    .A1(_18479_),
    .A2(_19406_),
    .ZN(_19407_)
  );
  INV_X1 _55147_ (
    .A(_19407_),
    .ZN(_19408_)
  );
  AND2_X1 _55148_ (
    .A1(count_instr[18]),
    .A2(instr_rdinstr),
    .ZN(_19409_)
  );
  INV_X1 _55149_ (
    .A(_19409_),
    .ZN(_19410_)
  );
  AND2_X1 _55150_ (
    .A1(instr_rdcycleh),
    .A2(count_cycle[50]),
    .ZN(_19411_)
  );
  INV_X1 _55151_ (
    .A(_19411_),
    .ZN(_19412_)
  );
  AND2_X1 _55152_ (
    .A1(_19410_),
    .A2(_19412_),
    .ZN(_19413_)
  );
  AND2_X1 _55153_ (
    .A1(count_instr[50]),
    .A2(instr_rdinstrh),
    .ZN(_19414_)
  );
  INV_X1 _55154_ (
    .A(_19414_),
    .ZN(_19415_)
  );
  AND2_X1 _55155_ (
    .A1(instr_rdcycle),
    .A2(count_cycle[18]),
    .ZN(_19416_)
  );
  INV_X1 _55156_ (
    .A(_19416_),
    .ZN(_19417_)
  );
  AND2_X1 _55157_ (
    .A1(_19415_),
    .A2(_19417_),
    .ZN(_19418_)
  );
  AND2_X1 _55158_ (
    .A1(_19413_),
    .A2(_19418_),
    .ZN(_19419_)
  );
  INV_X1 _55159_ (
    .A(_19419_),
    .ZN(_19420_)
  );
  AND2_X1 _55160_ (
    .A1(_22271_),
    .A2(_19420_),
    .ZN(_19421_)
  );
  INV_X1 _55161_ (
    .A(_19421_),
    .ZN(_19422_)
  );
  AND2_X1 _55162_ (
    .A1(reg_op1[18]),
    .A2(_22282_),
    .ZN(_19423_)
  );
  INV_X1 _55163_ (
    .A(_19423_),
    .ZN(_19424_)
  );
  AND2_X1 _55164_ (
    .A1(_19422_),
    .A2(_19424_),
    .ZN(_19425_)
  );
  AND2_X1 _55165_ (
    .A1(_19408_),
    .A2(_19425_),
    .ZN(_19426_)
  );
  AND2_X1 _55166_ (
    .A1(_19401_),
    .A2(_19426_),
    .ZN(_19427_)
  );
  INV_X1 _55167_ (
    .A(_19427_),
    .ZN(_19428_)
  );
  AND2_X1 _55168_ (
    .A1(resetn),
    .A2(_19428_),
    .ZN(_00005_[18])
  );
  AND2_X1 _55169_ (
    .A1(_19384_),
    .A2(_19396_),
    .ZN(_19429_)
  );
  INV_X1 _55170_ (
    .A(_19429_),
    .ZN(_19430_)
  );
  AND2_X1 _55171_ (
    .A1(reg_pc[19]),
    .A2(decoded_imm[19]),
    .ZN(_19431_)
  );
  INV_X1 _55172_ (
    .A(_19431_),
    .ZN(_19432_)
  );
  AND2_X1 _55173_ (
    .A1(_21085_),
    .A2(_21990_),
    .ZN(_19433_)
  );
  INV_X1 _55174_ (
    .A(_19433_),
    .ZN(_19434_)
  );
  AND2_X1 _55175_ (
    .A1(_19432_),
    .A2(_19434_),
    .ZN(_19435_)
  );
  INV_X1 _55176_ (
    .A(_19435_),
    .ZN(_19436_)
  );
  AND2_X1 _55177_ (
    .A1(_19430_),
    .A2(_19435_),
    .ZN(_19437_)
  );
  INV_X1 _55178_ (
    .A(_19437_),
    .ZN(_19438_)
  );
  AND2_X1 _55179_ (
    .A1(_19429_),
    .A2(_19436_),
    .ZN(_19439_)
  );
  INV_X1 _55180_ (
    .A(_19439_),
    .ZN(_19440_)
  );
  AND2_X1 _55181_ (
    .A1(_11090_),
    .A2(_19440_),
    .ZN(_19441_)
  );
  AND2_X1 _55182_ (
    .A1(_19438_),
    .A2(_19441_),
    .ZN(_19442_)
  );
  INV_X1 _55183_ (
    .A(_19442_),
    .ZN(_19443_)
  );
  AND2_X1 _55184_ (
    .A1(latched_is_lu),
    .A2(mem_rdata[19]),
    .ZN(_19444_)
  );
  AND2_X1 _55185_ (
    .A1(_12194_),
    .A2(_19444_),
    .ZN(_19445_)
  );
  INV_X1 _55186_ (
    .A(_19445_),
    .ZN(_19446_)
  );
  AND2_X1 _55187_ (
    .A1(_19313_),
    .A2(_19446_),
    .ZN(_19447_)
  );
  INV_X1 _55188_ (
    .A(_19447_),
    .ZN(_19448_)
  );
  AND2_X1 _55189_ (
    .A1(_18479_),
    .A2(_19448_),
    .ZN(_19449_)
  );
  INV_X1 _55190_ (
    .A(_19449_),
    .ZN(_19450_)
  );
  AND2_X1 _55191_ (
    .A1(reg_op1[19]),
    .A2(_22282_),
    .ZN(_19451_)
  );
  INV_X1 _55192_ (
    .A(_19451_),
    .ZN(_19452_)
  );
  AND2_X1 _55193_ (
    .A1(count_instr[19]),
    .A2(instr_rdinstr),
    .ZN(_19453_)
  );
  INV_X1 _55194_ (
    .A(_19453_),
    .ZN(_19454_)
  );
  AND2_X1 _55195_ (
    .A1(instr_rdcycleh),
    .A2(count_cycle[51]),
    .ZN(_19455_)
  );
  INV_X1 _55196_ (
    .A(_19455_),
    .ZN(_19456_)
  );
  AND2_X1 _55197_ (
    .A1(_19454_),
    .A2(_19456_),
    .ZN(_19457_)
  );
  AND2_X1 _55198_ (
    .A1(count_instr[51]),
    .A2(instr_rdinstrh),
    .ZN(_19458_)
  );
  INV_X1 _55199_ (
    .A(_19458_),
    .ZN(_19459_)
  );
  AND2_X1 _55200_ (
    .A1(instr_rdcycle),
    .A2(count_cycle[19]),
    .ZN(_19460_)
  );
  INV_X1 _55201_ (
    .A(_19460_),
    .ZN(_19461_)
  );
  AND2_X1 _55202_ (
    .A1(_19459_),
    .A2(_19461_),
    .ZN(_19462_)
  );
  AND2_X1 _55203_ (
    .A1(_19457_),
    .A2(_19462_),
    .ZN(_19463_)
  );
  INV_X1 _55204_ (
    .A(_19463_),
    .ZN(_19464_)
  );
  AND2_X1 _55205_ (
    .A1(_22271_),
    .A2(_19464_),
    .ZN(_19465_)
  );
  INV_X1 _55206_ (
    .A(_19465_),
    .ZN(_19466_)
  );
  AND2_X1 _55207_ (
    .A1(_19452_),
    .A2(_19466_),
    .ZN(_19467_)
  );
  AND2_X1 _55208_ (
    .A1(_19450_),
    .A2(_19467_),
    .ZN(_19468_)
  );
  AND2_X1 _55209_ (
    .A1(_19443_),
    .A2(_19468_),
    .ZN(_19469_)
  );
  INV_X1 _55210_ (
    .A(_19469_),
    .ZN(_19470_)
  );
  AND2_X1 _55211_ (
    .A1(resetn),
    .A2(_19470_),
    .ZN(_00005_[19])
  );
  AND2_X1 _55212_ (
    .A1(latched_is_lu),
    .A2(mem_rdata[20]),
    .ZN(_19471_)
  );
  AND2_X1 _55213_ (
    .A1(_12194_),
    .A2(_19471_),
    .ZN(_19472_)
  );
  INV_X1 _55214_ (
    .A(_19472_),
    .ZN(_19473_)
  );
  AND2_X1 _55215_ (
    .A1(_19313_),
    .A2(_19473_),
    .ZN(_19474_)
  );
  INV_X1 _55216_ (
    .A(_19474_),
    .ZN(_19475_)
  );
  AND2_X1 _55217_ (
    .A1(_18479_),
    .A2(_19475_),
    .ZN(_19476_)
  );
  INV_X1 _55218_ (
    .A(_19476_),
    .ZN(_19477_)
  );
  AND2_X1 _55219_ (
    .A1(reg_op1[20]),
    .A2(_22282_),
    .ZN(_19478_)
  );
  INV_X1 _55220_ (
    .A(_19478_),
    .ZN(_19479_)
  );
  AND2_X1 _55221_ (
    .A1(count_instr[20]),
    .A2(instr_rdinstr),
    .ZN(_19480_)
  );
  INV_X1 _55222_ (
    .A(_19480_),
    .ZN(_19481_)
  );
  AND2_X1 _55223_ (
    .A1(instr_rdcycleh),
    .A2(count_cycle[52]),
    .ZN(_19482_)
  );
  INV_X1 _55224_ (
    .A(_19482_),
    .ZN(_19483_)
  );
  AND2_X1 _55225_ (
    .A1(_19481_),
    .A2(_19483_),
    .ZN(_19484_)
  );
  AND2_X1 _55226_ (
    .A1(count_instr[52]),
    .A2(instr_rdinstrh),
    .ZN(_19485_)
  );
  INV_X1 _55227_ (
    .A(_19485_),
    .ZN(_19486_)
  );
  AND2_X1 _55228_ (
    .A1(instr_rdcycle),
    .A2(count_cycle[20]),
    .ZN(_19487_)
  );
  INV_X1 _55229_ (
    .A(_19487_),
    .ZN(_19488_)
  );
  AND2_X1 _55230_ (
    .A1(_19486_),
    .A2(_19488_),
    .ZN(_19489_)
  );
  AND2_X1 _55231_ (
    .A1(_19484_),
    .A2(_19489_),
    .ZN(_19490_)
  );
  INV_X1 _55232_ (
    .A(_19490_),
    .ZN(_19491_)
  );
  AND2_X1 _55233_ (
    .A1(_22271_),
    .A2(_19491_),
    .ZN(_19492_)
  );
  INV_X1 _55234_ (
    .A(_19492_),
    .ZN(_19493_)
  );
  AND2_X1 _55235_ (
    .A1(_19479_),
    .A2(_19493_),
    .ZN(_19494_)
  );
  AND2_X1 _55236_ (
    .A1(reg_pc[20]),
    .A2(decoded_imm[20]),
    .ZN(_19495_)
  );
  INV_X1 _55237_ (
    .A(_19495_),
    .ZN(_19496_)
  );
  AND2_X1 _55238_ (
    .A1(_21084_),
    .A2(_21989_),
    .ZN(_19497_)
  );
  INV_X1 _55239_ (
    .A(_19497_),
    .ZN(_19498_)
  );
  AND2_X1 _55240_ (
    .A1(_19496_),
    .A2(_19498_),
    .ZN(_19499_)
  );
  INV_X1 _55241_ (
    .A(_19499_),
    .ZN(_19500_)
  );
  AND2_X1 _55242_ (
    .A1(_19429_),
    .A2(_19432_),
    .ZN(_19501_)
  );
  INV_X1 _55243_ (
    .A(_19501_),
    .ZN(_19502_)
  );
  AND2_X1 _55244_ (
    .A1(_19430_),
    .A2(_19434_),
    .ZN(_19503_)
  );
  INV_X1 _55245_ (
    .A(_19503_),
    .ZN(_19504_)
  );
  AND2_X1 _55246_ (
    .A1(_19434_),
    .A2(_19502_),
    .ZN(_19505_)
  );
  AND2_X1 _55247_ (
    .A1(_19432_),
    .A2(_19504_),
    .ZN(_19506_)
  );
  AND2_X1 _55248_ (
    .A1(_19500_),
    .A2(_19506_),
    .ZN(_19507_)
  );
  INV_X1 _55249_ (
    .A(_19507_),
    .ZN(_19508_)
  );
  AND2_X1 _55250_ (
    .A1(_19499_),
    .A2(_19505_),
    .ZN(_19509_)
  );
  INV_X1 _55251_ (
    .A(_19509_),
    .ZN(_19510_)
  );
  AND2_X1 _55252_ (
    .A1(_11090_),
    .A2(_19510_),
    .ZN(_19511_)
  );
  AND2_X1 _55253_ (
    .A1(_19508_),
    .A2(_19511_),
    .ZN(_19512_)
  );
  INV_X1 _55254_ (
    .A(_19512_),
    .ZN(_19513_)
  );
  AND2_X1 _55255_ (
    .A1(_19494_),
    .A2(_19513_),
    .ZN(_19514_)
  );
  AND2_X1 _55256_ (
    .A1(_19477_),
    .A2(_19514_),
    .ZN(_19515_)
  );
  INV_X1 _55257_ (
    .A(_19515_),
    .ZN(_19516_)
  );
  AND2_X1 _55258_ (
    .A1(resetn),
    .A2(_19516_),
    .ZN(_00005_[20])
  );
  AND2_X1 _55259_ (
    .A1(_19496_),
    .A2(_19510_),
    .ZN(_19517_)
  );
  INV_X1 _55260_ (
    .A(_19517_),
    .ZN(_19518_)
  );
  AND2_X1 _55261_ (
    .A1(reg_pc[21]),
    .A2(decoded_imm[21]),
    .ZN(_19519_)
  );
  INV_X1 _55262_ (
    .A(_19519_),
    .ZN(_19520_)
  );
  AND2_X1 _55263_ (
    .A1(_21083_),
    .A2(_21988_),
    .ZN(_19521_)
  );
  INV_X1 _55264_ (
    .A(_19521_),
    .ZN(_19522_)
  );
  AND2_X1 _55265_ (
    .A1(_19520_),
    .A2(_19522_),
    .ZN(_19523_)
  );
  INV_X1 _55266_ (
    .A(_19523_),
    .ZN(_19524_)
  );
  AND2_X1 _55267_ (
    .A1(_19517_),
    .A2(_19524_),
    .ZN(_19525_)
  );
  INV_X1 _55268_ (
    .A(_19525_),
    .ZN(_19526_)
  );
  AND2_X1 _55269_ (
    .A1(_19518_),
    .A2(_19523_),
    .ZN(_19527_)
  );
  INV_X1 _55270_ (
    .A(_19527_),
    .ZN(_19528_)
  );
  AND2_X1 _55271_ (
    .A1(_19526_),
    .A2(_19528_),
    .ZN(_19529_)
  );
  AND2_X1 _55272_ (
    .A1(_11090_),
    .A2(_19529_),
    .ZN(_19530_)
  );
  INV_X1 _55273_ (
    .A(_19530_),
    .ZN(_19531_)
  );
  AND2_X1 _55274_ (
    .A1(latched_is_lu),
    .A2(mem_rdata[21]),
    .ZN(_19532_)
  );
  AND2_X1 _55275_ (
    .A1(_12194_),
    .A2(_19532_),
    .ZN(_19533_)
  );
  INV_X1 _55276_ (
    .A(_19533_),
    .ZN(_19534_)
  );
  AND2_X1 _55277_ (
    .A1(_19313_),
    .A2(_19534_),
    .ZN(_19535_)
  );
  INV_X1 _55278_ (
    .A(_19535_),
    .ZN(_19536_)
  );
  AND2_X1 _55279_ (
    .A1(_18479_),
    .A2(_19536_),
    .ZN(_19537_)
  );
  INV_X1 _55280_ (
    .A(_19537_),
    .ZN(_19538_)
  );
  AND2_X1 _55281_ (
    .A1(reg_op1[21]),
    .A2(_22282_),
    .ZN(_19539_)
  );
  INV_X1 _55282_ (
    .A(_19539_),
    .ZN(_19540_)
  );
  AND2_X1 _55283_ (
    .A1(count_instr[21]),
    .A2(instr_rdinstr),
    .ZN(_19541_)
  );
  INV_X1 _55284_ (
    .A(_19541_),
    .ZN(_19542_)
  );
  AND2_X1 _55285_ (
    .A1(instr_rdcycleh),
    .A2(count_cycle[53]),
    .ZN(_19543_)
  );
  INV_X1 _55286_ (
    .A(_19543_),
    .ZN(_19544_)
  );
  AND2_X1 _55287_ (
    .A1(_19542_),
    .A2(_19544_),
    .ZN(_19545_)
  );
  AND2_X1 _55288_ (
    .A1(count_instr[53]),
    .A2(instr_rdinstrh),
    .ZN(_19546_)
  );
  INV_X1 _55289_ (
    .A(_19546_),
    .ZN(_19547_)
  );
  AND2_X1 _55290_ (
    .A1(instr_rdcycle),
    .A2(count_cycle[21]),
    .ZN(_19548_)
  );
  INV_X1 _55291_ (
    .A(_19548_),
    .ZN(_19549_)
  );
  AND2_X1 _55292_ (
    .A1(_19547_),
    .A2(_19549_),
    .ZN(_19550_)
  );
  AND2_X1 _55293_ (
    .A1(_19545_),
    .A2(_19550_),
    .ZN(_19551_)
  );
  INV_X1 _55294_ (
    .A(_19551_),
    .ZN(_19552_)
  );
  AND2_X1 _55295_ (
    .A1(_22271_),
    .A2(_19552_),
    .ZN(_19553_)
  );
  INV_X1 _55296_ (
    .A(_19553_),
    .ZN(_19554_)
  );
  AND2_X1 _55297_ (
    .A1(_19540_),
    .A2(_19554_),
    .ZN(_19555_)
  );
  AND2_X1 _55298_ (
    .A1(_19538_),
    .A2(_19555_),
    .ZN(_19556_)
  );
  AND2_X1 _55299_ (
    .A1(_19531_),
    .A2(_19556_),
    .ZN(_19557_)
  );
  INV_X1 _55300_ (
    .A(_19557_),
    .ZN(_19558_)
  );
  AND2_X1 _55301_ (
    .A1(resetn),
    .A2(_19558_),
    .ZN(_00005_[21])
  );
  AND2_X1 _55302_ (
    .A1(reg_pc[22]),
    .A2(decoded_imm[22]),
    .ZN(_19559_)
  );
  INV_X1 _55303_ (
    .A(_19559_),
    .ZN(_19560_)
  );
  AND2_X1 _55304_ (
    .A1(_21082_),
    .A2(_21987_),
    .ZN(_19561_)
  );
  INV_X1 _55305_ (
    .A(_19561_),
    .ZN(_19562_)
  );
  AND2_X1 _55306_ (
    .A1(_19560_),
    .A2(_19562_),
    .ZN(_19563_)
  );
  INV_X1 _55307_ (
    .A(_19563_),
    .ZN(_19564_)
  );
  AND2_X1 _55308_ (
    .A1(_19517_),
    .A2(_19520_),
    .ZN(_19565_)
  );
  INV_X1 _55309_ (
    .A(_19565_),
    .ZN(_19566_)
  );
  AND2_X1 _55310_ (
    .A1(_19518_),
    .A2(_19522_),
    .ZN(_19567_)
  );
  INV_X1 _55311_ (
    .A(_19567_),
    .ZN(_19568_)
  );
  AND2_X1 _55312_ (
    .A1(_19522_),
    .A2(_19566_),
    .ZN(_19569_)
  );
  AND2_X1 _55313_ (
    .A1(_19520_),
    .A2(_19568_),
    .ZN(_19570_)
  );
  AND2_X1 _55314_ (
    .A1(_19563_),
    .A2(_19569_),
    .ZN(_19571_)
  );
  INV_X1 _55315_ (
    .A(_19571_),
    .ZN(_19572_)
  );
  AND2_X1 _55316_ (
    .A1(_19564_),
    .A2(_19570_),
    .ZN(_19573_)
  );
  INV_X1 _55317_ (
    .A(_19573_),
    .ZN(_19574_)
  );
  AND2_X1 _55318_ (
    .A1(_11090_),
    .A2(_19572_),
    .ZN(_19575_)
  );
  AND2_X1 _55319_ (
    .A1(_19574_),
    .A2(_19575_),
    .ZN(_19576_)
  );
  INV_X1 _55320_ (
    .A(_19576_),
    .ZN(_19577_)
  );
  AND2_X1 _55321_ (
    .A1(latched_is_lu),
    .A2(mem_rdata[22]),
    .ZN(_19578_)
  );
  AND2_X1 _55322_ (
    .A1(_12194_),
    .A2(_19578_),
    .ZN(_19579_)
  );
  INV_X1 _55323_ (
    .A(_19579_),
    .ZN(_19580_)
  );
  AND2_X1 _55324_ (
    .A1(_19313_),
    .A2(_19580_),
    .ZN(_19581_)
  );
  INV_X1 _55325_ (
    .A(_19581_),
    .ZN(_19582_)
  );
  AND2_X1 _55326_ (
    .A1(_18479_),
    .A2(_19582_),
    .ZN(_19583_)
  );
  INV_X1 _55327_ (
    .A(_19583_),
    .ZN(_19584_)
  );
  AND2_X1 _55328_ (
    .A1(reg_op1[22]),
    .A2(_22282_),
    .ZN(_19585_)
  );
  INV_X1 _55329_ (
    .A(_19585_),
    .ZN(_19586_)
  );
  AND2_X1 _55330_ (
    .A1(count_instr[54]),
    .A2(instr_rdinstrh),
    .ZN(_19587_)
  );
  INV_X1 _55331_ (
    .A(_19587_),
    .ZN(_19588_)
  );
  AND2_X1 _55332_ (
    .A1(count_instr[22]),
    .A2(instr_rdinstr),
    .ZN(_19589_)
  );
  INV_X1 _55333_ (
    .A(_19589_),
    .ZN(_19590_)
  );
  AND2_X1 _55334_ (
    .A1(_19588_),
    .A2(_19590_),
    .ZN(_19591_)
  );
  AND2_X1 _55335_ (
    .A1(instr_rdcycle),
    .A2(count_cycle[22]),
    .ZN(_19592_)
  );
  INV_X1 _55336_ (
    .A(_19592_),
    .ZN(_19593_)
  );
  AND2_X1 _55337_ (
    .A1(instr_rdcycleh),
    .A2(count_cycle[54]),
    .ZN(_19594_)
  );
  INV_X1 _55338_ (
    .A(_19594_),
    .ZN(_19595_)
  );
  AND2_X1 _55339_ (
    .A1(_19593_),
    .A2(_19595_),
    .ZN(_19596_)
  );
  AND2_X1 _55340_ (
    .A1(_19591_),
    .A2(_19596_),
    .ZN(_19597_)
  );
  INV_X1 _55341_ (
    .A(_19597_),
    .ZN(_19598_)
  );
  AND2_X1 _55342_ (
    .A1(_22271_),
    .A2(_19598_),
    .ZN(_19599_)
  );
  INV_X1 _55343_ (
    .A(_19599_),
    .ZN(_19600_)
  );
  AND2_X1 _55344_ (
    .A1(_19586_),
    .A2(_19600_),
    .ZN(_19601_)
  );
  AND2_X1 _55345_ (
    .A1(_19584_),
    .A2(_19601_),
    .ZN(_19602_)
  );
  AND2_X1 _55346_ (
    .A1(_19577_),
    .A2(_19602_),
    .ZN(_19603_)
  );
  INV_X1 _55347_ (
    .A(_19603_),
    .ZN(_19604_)
  );
  AND2_X1 _55348_ (
    .A1(resetn),
    .A2(_19604_),
    .ZN(_00005_[22])
  );
  AND2_X1 _55349_ (
    .A1(latched_is_lu),
    .A2(mem_rdata[23]),
    .ZN(_19605_)
  );
  AND2_X1 _55350_ (
    .A1(_12194_),
    .A2(_19605_),
    .ZN(_19606_)
  );
  INV_X1 _55351_ (
    .A(_19606_),
    .ZN(_19607_)
  );
  AND2_X1 _55352_ (
    .A1(_19313_),
    .A2(_19607_),
    .ZN(_19608_)
  );
  INV_X1 _55353_ (
    .A(_19608_),
    .ZN(_19609_)
  );
  AND2_X1 _55354_ (
    .A1(_18479_),
    .A2(_19609_),
    .ZN(_19610_)
  );
  INV_X1 _55355_ (
    .A(_19610_),
    .ZN(_19611_)
  );
  AND2_X1 _55356_ (
    .A1(count_instr[55]),
    .A2(instr_rdinstrh),
    .ZN(_19612_)
  );
  INV_X1 _55357_ (
    .A(_19612_),
    .ZN(_19613_)
  );
  AND2_X1 _55358_ (
    .A1(count_instr[23]),
    .A2(instr_rdinstr),
    .ZN(_19614_)
  );
  INV_X1 _55359_ (
    .A(_19614_),
    .ZN(_19615_)
  );
  AND2_X1 _55360_ (
    .A1(_19613_),
    .A2(_19615_),
    .ZN(_19616_)
  );
  AND2_X1 _55361_ (
    .A1(instr_rdcycle),
    .A2(count_cycle[23]),
    .ZN(_19617_)
  );
  INV_X1 _55362_ (
    .A(_19617_),
    .ZN(_19618_)
  );
  AND2_X1 _55363_ (
    .A1(instr_rdcycleh),
    .A2(count_cycle[55]),
    .ZN(_19619_)
  );
  INV_X1 _55364_ (
    .A(_19619_),
    .ZN(_19620_)
  );
  AND2_X1 _55365_ (
    .A1(_19618_),
    .A2(_19620_),
    .ZN(_19621_)
  );
  AND2_X1 _55366_ (
    .A1(_19616_),
    .A2(_19621_),
    .ZN(_19622_)
  );
  INV_X1 _55367_ (
    .A(_19622_),
    .ZN(_19623_)
  );
  AND2_X1 _55368_ (
    .A1(_22271_),
    .A2(_19623_),
    .ZN(_19624_)
  );
  INV_X1 _55369_ (
    .A(_19624_),
    .ZN(_19625_)
  );
  AND2_X1 _55370_ (
    .A1(reg_op1[23]),
    .A2(_22282_),
    .ZN(_19626_)
  );
  INV_X1 _55371_ (
    .A(_19626_),
    .ZN(_19627_)
  );
  AND2_X1 _55372_ (
    .A1(_19625_),
    .A2(_19627_),
    .ZN(_19628_)
  );
  AND2_X1 _55373_ (
    .A1(_19611_),
    .A2(_19628_),
    .ZN(_19629_)
  );
  AND2_X1 _55374_ (
    .A1(_19560_),
    .A2(_19572_),
    .ZN(_19630_)
  );
  INV_X1 _55375_ (
    .A(_19630_),
    .ZN(_19631_)
  );
  AND2_X1 _55376_ (
    .A1(reg_pc[23]),
    .A2(decoded_imm[23]),
    .ZN(_19632_)
  );
  INV_X1 _55377_ (
    .A(_19632_),
    .ZN(_19633_)
  );
  AND2_X1 _55378_ (
    .A1(_21081_),
    .A2(_21986_),
    .ZN(_19634_)
  );
  INV_X1 _55379_ (
    .A(_19634_),
    .ZN(_19635_)
  );
  AND2_X1 _55380_ (
    .A1(_19633_),
    .A2(_19635_),
    .ZN(_19636_)
  );
  INV_X1 _55381_ (
    .A(_19636_),
    .ZN(_19637_)
  );
  AND2_X1 _55382_ (
    .A1(_19630_),
    .A2(_19636_),
    .ZN(_19638_)
  );
  INV_X1 _55383_ (
    .A(_19638_),
    .ZN(_19639_)
  );
  AND2_X1 _55384_ (
    .A1(_19631_),
    .A2(_19637_),
    .ZN(_19640_)
  );
  INV_X1 _55385_ (
    .A(_19640_),
    .ZN(_19641_)
  );
  AND2_X1 _55386_ (
    .A1(_19639_),
    .A2(_19641_),
    .ZN(_19642_)
  );
  INV_X1 _55387_ (
    .A(_19642_),
    .ZN(_19643_)
  );
  AND2_X1 _55388_ (
    .A1(_11090_),
    .A2(_19643_),
    .ZN(_19644_)
  );
  INV_X1 _55389_ (
    .A(_19644_),
    .ZN(_19645_)
  );
  AND2_X1 _55390_ (
    .A1(_19629_),
    .A2(_19645_),
    .ZN(_19646_)
  );
  INV_X1 _55391_ (
    .A(_19646_),
    .ZN(_19647_)
  );
  AND2_X1 _55392_ (
    .A1(resetn),
    .A2(_19647_),
    .ZN(_00005_[23])
  );
  AND2_X1 _55393_ (
    .A1(reg_pc[24]),
    .A2(decoded_imm[24]),
    .ZN(_19648_)
  );
  INV_X1 _55394_ (
    .A(_19648_),
    .ZN(_19649_)
  );
  AND2_X1 _55395_ (
    .A1(_21080_),
    .A2(_21985_),
    .ZN(_19650_)
  );
  INV_X1 _55396_ (
    .A(_19650_),
    .ZN(_19651_)
  );
  AND2_X1 _55397_ (
    .A1(_19649_),
    .A2(_19651_),
    .ZN(_19652_)
  );
  INV_X1 _55398_ (
    .A(_19652_),
    .ZN(_19653_)
  );
  AND2_X1 _55399_ (
    .A1(_19630_),
    .A2(_19633_),
    .ZN(_19654_)
  );
  INV_X1 _55400_ (
    .A(_19654_),
    .ZN(_19655_)
  );
  AND2_X1 _55401_ (
    .A1(_19631_),
    .A2(_19635_),
    .ZN(_19656_)
  );
  INV_X1 _55402_ (
    .A(_19656_),
    .ZN(_19657_)
  );
  AND2_X1 _55403_ (
    .A1(_19635_),
    .A2(_19655_),
    .ZN(_19658_)
  );
  AND2_X1 _55404_ (
    .A1(_19633_),
    .A2(_19657_),
    .ZN(_19659_)
  );
  AND2_X1 _55405_ (
    .A1(_19652_),
    .A2(_19658_),
    .ZN(_19660_)
  );
  INV_X1 _55406_ (
    .A(_19660_),
    .ZN(_19661_)
  );
  AND2_X1 _55407_ (
    .A1(_19653_),
    .A2(_19659_),
    .ZN(_19662_)
  );
  INV_X1 _55408_ (
    .A(_19662_),
    .ZN(_19663_)
  );
  AND2_X1 _55409_ (
    .A1(_11090_),
    .A2(_19661_),
    .ZN(_19664_)
  );
  AND2_X1 _55410_ (
    .A1(_19663_),
    .A2(_19664_),
    .ZN(_19665_)
  );
  INV_X1 _55411_ (
    .A(_19665_),
    .ZN(_19666_)
  );
  AND2_X1 _55412_ (
    .A1(latched_is_lu),
    .A2(mem_rdata[24]),
    .ZN(_19667_)
  );
  AND2_X1 _55413_ (
    .A1(_12194_),
    .A2(_19667_),
    .ZN(_19668_)
  );
  INV_X1 _55414_ (
    .A(_19668_),
    .ZN(_19669_)
  );
  AND2_X1 _55415_ (
    .A1(_19313_),
    .A2(_19669_),
    .ZN(_19670_)
  );
  INV_X1 _55416_ (
    .A(_19670_),
    .ZN(_19671_)
  );
  AND2_X1 _55417_ (
    .A1(_18479_),
    .A2(_19671_),
    .ZN(_19672_)
  );
  INV_X1 _55418_ (
    .A(_19672_),
    .ZN(_19673_)
  );
  AND2_X1 _55419_ (
    .A1(count_instr[24]),
    .A2(instr_rdinstr),
    .ZN(_19674_)
  );
  INV_X1 _55420_ (
    .A(_19674_),
    .ZN(_19675_)
  );
  AND2_X1 _55421_ (
    .A1(instr_rdcycleh),
    .A2(count_cycle[56]),
    .ZN(_19676_)
  );
  INV_X1 _55422_ (
    .A(_19676_),
    .ZN(_19677_)
  );
  AND2_X1 _55423_ (
    .A1(_19675_),
    .A2(_19677_),
    .ZN(_19678_)
  );
  AND2_X1 _55424_ (
    .A1(count_instr[56]),
    .A2(instr_rdinstrh),
    .ZN(_19679_)
  );
  INV_X1 _55425_ (
    .A(_19679_),
    .ZN(_19680_)
  );
  AND2_X1 _55426_ (
    .A1(instr_rdcycle),
    .A2(count_cycle[24]),
    .ZN(_19681_)
  );
  INV_X1 _55427_ (
    .A(_19681_),
    .ZN(_19682_)
  );
  AND2_X1 _55428_ (
    .A1(_19680_),
    .A2(_19682_),
    .ZN(_19683_)
  );
  AND2_X1 _55429_ (
    .A1(_19678_),
    .A2(_19683_),
    .ZN(_19684_)
  );
  INV_X1 _55430_ (
    .A(_19684_),
    .ZN(_19685_)
  );
  AND2_X1 _55431_ (
    .A1(_22271_),
    .A2(_19685_),
    .ZN(_19686_)
  );
  INV_X1 _55432_ (
    .A(_19686_),
    .ZN(_19687_)
  );
  AND2_X1 _55433_ (
    .A1(reg_op1[24]),
    .A2(_22282_),
    .ZN(_19688_)
  );
  INV_X1 _55434_ (
    .A(_19688_),
    .ZN(_19689_)
  );
  AND2_X1 _55435_ (
    .A1(_19687_),
    .A2(_19689_),
    .ZN(_19690_)
  );
  AND2_X1 _55436_ (
    .A1(_19673_),
    .A2(_19690_),
    .ZN(_19691_)
  );
  AND2_X1 _55437_ (
    .A1(_19666_),
    .A2(_19691_),
    .ZN(_19692_)
  );
  INV_X1 _55438_ (
    .A(_19692_),
    .ZN(_19693_)
  );
  AND2_X1 _55439_ (
    .A1(resetn),
    .A2(_19693_),
    .ZN(_00005_[24])
  );
  AND2_X1 _55440_ (
    .A1(latched_is_lu),
    .A2(mem_rdata[25]),
    .ZN(_19694_)
  );
  AND2_X1 _55441_ (
    .A1(_12194_),
    .A2(_19694_),
    .ZN(_19695_)
  );
  INV_X1 _55442_ (
    .A(_19695_),
    .ZN(_19696_)
  );
  AND2_X1 _55443_ (
    .A1(_19313_),
    .A2(_19696_),
    .ZN(_19697_)
  );
  INV_X1 _55444_ (
    .A(_19697_),
    .ZN(_19698_)
  );
  AND2_X1 _55445_ (
    .A1(_18479_),
    .A2(_19698_),
    .ZN(_19699_)
  );
  INV_X1 _55446_ (
    .A(_19699_),
    .ZN(_19700_)
  );
  AND2_X1 _55447_ (
    .A1(reg_op1[25]),
    .A2(_22282_),
    .ZN(_19701_)
  );
  INV_X1 _55448_ (
    .A(_19701_),
    .ZN(_19702_)
  );
  AND2_X1 _55449_ (
    .A1(count_instr[25]),
    .A2(instr_rdinstr),
    .ZN(_19703_)
  );
  INV_X1 _55450_ (
    .A(_19703_),
    .ZN(_19704_)
  );
  AND2_X1 _55451_ (
    .A1(instr_rdcycleh),
    .A2(count_cycle[57]),
    .ZN(_19705_)
  );
  INV_X1 _55452_ (
    .A(_19705_),
    .ZN(_19706_)
  );
  AND2_X1 _55453_ (
    .A1(_19704_),
    .A2(_19706_),
    .ZN(_19707_)
  );
  AND2_X1 _55454_ (
    .A1(instr_rdcycle),
    .A2(count_cycle[25]),
    .ZN(_19708_)
  );
  INV_X1 _55455_ (
    .A(_19708_),
    .ZN(_19709_)
  );
  AND2_X1 _55456_ (
    .A1(count_instr[57]),
    .A2(instr_rdinstrh),
    .ZN(_19710_)
  );
  INV_X1 _55457_ (
    .A(_19710_),
    .ZN(_19711_)
  );
  AND2_X1 _55458_ (
    .A1(_19709_),
    .A2(_19711_),
    .ZN(_19712_)
  );
  AND2_X1 _55459_ (
    .A1(_19707_),
    .A2(_19712_),
    .ZN(_19713_)
  );
  INV_X1 _55460_ (
    .A(_19713_),
    .ZN(_19714_)
  );
  AND2_X1 _55461_ (
    .A1(_22271_),
    .A2(_19714_),
    .ZN(_19715_)
  );
  INV_X1 _55462_ (
    .A(_19715_),
    .ZN(_19716_)
  );
  AND2_X1 _55463_ (
    .A1(_19702_),
    .A2(_19716_),
    .ZN(_19717_)
  );
  AND2_X1 _55464_ (
    .A1(_19700_),
    .A2(_19717_),
    .ZN(_19718_)
  );
  INV_X1 _55465_ (
    .A(_19718_),
    .ZN(_19719_)
  );
  AND2_X1 _55466_ (
    .A1(resetn),
    .A2(_19719_),
    .ZN(_19720_)
  );
  INV_X1 _55467_ (
    .A(_19720_),
    .ZN(_19721_)
  );
  AND2_X1 _55468_ (
    .A1(_19649_),
    .A2(_19661_),
    .ZN(_19722_)
  );
  INV_X1 _55469_ (
    .A(_19722_),
    .ZN(_19723_)
  );
  AND2_X1 _55470_ (
    .A1(reg_pc[25]),
    .A2(decoded_imm[25]),
    .ZN(_19724_)
  );
  INV_X1 _55471_ (
    .A(_19724_),
    .ZN(_19725_)
  );
  AND2_X1 _55472_ (
    .A1(_21079_),
    .A2(_21984_),
    .ZN(_19726_)
  );
  INV_X1 _55473_ (
    .A(_19726_),
    .ZN(_19727_)
  );
  AND2_X1 _55474_ (
    .A1(_19725_),
    .A2(_19727_),
    .ZN(_19728_)
  );
  INV_X1 _55475_ (
    .A(_19728_),
    .ZN(_19729_)
  );
  AND2_X1 _55476_ (
    .A1(_19723_),
    .A2(_19728_),
    .ZN(_19730_)
  );
  INV_X1 _55477_ (
    .A(_19730_),
    .ZN(_19731_)
  );
  AND2_X1 _55478_ (
    .A1(_19722_),
    .A2(_19729_),
    .ZN(_19732_)
  );
  INV_X1 _55479_ (
    .A(_19732_),
    .ZN(_19733_)
  );
  AND2_X1 _55480_ (
    .A1(_11098_),
    .A2(_19733_),
    .ZN(_19734_)
  );
  AND2_X1 _55481_ (
    .A1(_19731_),
    .A2(_19734_),
    .ZN(_19735_)
  );
  INV_X1 _55482_ (
    .A(_19735_),
    .ZN(_19736_)
  );
  AND2_X1 _55483_ (
    .A1(_19721_),
    .A2(_19736_),
    .ZN(_19737_)
  );
  INV_X1 _55484_ (
    .A(_19737_),
    .ZN(_00005_[25])
  );
  AND2_X1 _55485_ (
    .A1(latched_is_lu),
    .A2(mem_rdata[26]),
    .ZN(_19738_)
  );
  AND2_X1 _55486_ (
    .A1(_12194_),
    .A2(_19738_),
    .ZN(_19739_)
  );
  INV_X1 _55487_ (
    .A(_19739_),
    .ZN(_19740_)
  );
  AND2_X1 _55488_ (
    .A1(_19313_),
    .A2(_19740_),
    .ZN(_19741_)
  );
  INV_X1 _55489_ (
    .A(_19741_),
    .ZN(_19742_)
  );
  AND2_X1 _55490_ (
    .A1(_18479_),
    .A2(_19742_),
    .ZN(_19743_)
  );
  INV_X1 _55491_ (
    .A(_19743_),
    .ZN(_19744_)
  );
  AND2_X1 _55492_ (
    .A1(reg_op1[26]),
    .A2(_22282_),
    .ZN(_19745_)
  );
  INV_X1 _55493_ (
    .A(_19745_),
    .ZN(_19746_)
  );
  AND2_X1 _55494_ (
    .A1(count_instr[26]),
    .A2(instr_rdinstr),
    .ZN(_19747_)
  );
  INV_X1 _55495_ (
    .A(_19747_),
    .ZN(_19748_)
  );
  AND2_X1 _55496_ (
    .A1(instr_rdcycleh),
    .A2(count_cycle[58]),
    .ZN(_19749_)
  );
  INV_X1 _55497_ (
    .A(_19749_),
    .ZN(_19750_)
  );
  AND2_X1 _55498_ (
    .A1(_19748_),
    .A2(_19750_),
    .ZN(_19751_)
  );
  AND2_X1 _55499_ (
    .A1(count_instr[58]),
    .A2(instr_rdinstrh),
    .ZN(_19752_)
  );
  INV_X1 _55500_ (
    .A(_19752_),
    .ZN(_19753_)
  );
  AND2_X1 _55501_ (
    .A1(instr_rdcycle),
    .A2(count_cycle[26]),
    .ZN(_19754_)
  );
  INV_X1 _55502_ (
    .A(_19754_),
    .ZN(_19755_)
  );
  AND2_X1 _55503_ (
    .A1(_19753_),
    .A2(_19755_),
    .ZN(_19756_)
  );
  AND2_X1 _55504_ (
    .A1(_19751_),
    .A2(_19756_),
    .ZN(_19757_)
  );
  INV_X1 _55505_ (
    .A(_19757_),
    .ZN(_19758_)
  );
  AND2_X1 _55506_ (
    .A1(_22271_),
    .A2(_19758_),
    .ZN(_19759_)
  );
  INV_X1 _55507_ (
    .A(_19759_),
    .ZN(_19760_)
  );
  AND2_X1 _55508_ (
    .A1(_19746_),
    .A2(_19760_),
    .ZN(_19761_)
  );
  AND2_X1 _55509_ (
    .A1(_19744_),
    .A2(_19761_),
    .ZN(_19762_)
  );
  AND2_X1 _55510_ (
    .A1(reg_pc[26]),
    .A2(decoded_imm[26]),
    .ZN(_19763_)
  );
  INV_X1 _55511_ (
    .A(_19763_),
    .ZN(_19764_)
  );
  AND2_X1 _55512_ (
    .A1(_21078_),
    .A2(_21983_),
    .ZN(_19765_)
  );
  INV_X1 _55513_ (
    .A(_19765_),
    .ZN(_19766_)
  );
  AND2_X1 _55514_ (
    .A1(_19764_),
    .A2(_19766_),
    .ZN(_19767_)
  );
  INV_X1 _55515_ (
    .A(_19767_),
    .ZN(_19768_)
  );
  AND2_X1 _55516_ (
    .A1(_19723_),
    .A2(_19727_),
    .ZN(_19769_)
  );
  INV_X1 _55517_ (
    .A(_19769_),
    .ZN(_19770_)
  );
  AND2_X1 _55518_ (
    .A1(_19722_),
    .A2(_19725_),
    .ZN(_19771_)
  );
  INV_X1 _55519_ (
    .A(_19771_),
    .ZN(_19772_)
  );
  AND2_X1 _55520_ (
    .A1(_19725_),
    .A2(_19770_),
    .ZN(_19773_)
  );
  AND2_X1 _55521_ (
    .A1(_19727_),
    .A2(_19772_),
    .ZN(_19774_)
  );
  AND2_X1 _55522_ (
    .A1(_19767_),
    .A2(_19774_),
    .ZN(_19775_)
  );
  INV_X1 _55523_ (
    .A(_19775_),
    .ZN(_19776_)
  );
  AND2_X1 _55524_ (
    .A1(_19768_),
    .A2(_19773_),
    .ZN(_19777_)
  );
  INV_X1 _55525_ (
    .A(_19777_),
    .ZN(_19778_)
  );
  AND2_X1 _55526_ (
    .A1(_11090_),
    .A2(_19778_),
    .ZN(_19779_)
  );
  AND2_X1 _55527_ (
    .A1(_19776_),
    .A2(_19779_),
    .ZN(_19780_)
  );
  INV_X1 _55528_ (
    .A(_19780_),
    .ZN(_19781_)
  );
  AND2_X1 _55529_ (
    .A1(_19762_),
    .A2(_19781_),
    .ZN(_19782_)
  );
  INV_X1 _55530_ (
    .A(_19782_),
    .ZN(_19783_)
  );
  AND2_X1 _55531_ (
    .A1(resetn),
    .A2(_19783_),
    .ZN(_00005_[26])
  );
  AND2_X1 _55532_ (
    .A1(latched_is_lu),
    .A2(mem_rdata[27]),
    .ZN(_19784_)
  );
  AND2_X1 _55533_ (
    .A1(_12194_),
    .A2(_19784_),
    .ZN(_19785_)
  );
  INV_X1 _55534_ (
    .A(_19785_),
    .ZN(_19786_)
  );
  AND2_X1 _55535_ (
    .A1(_19313_),
    .A2(_19786_),
    .ZN(_19787_)
  );
  INV_X1 _55536_ (
    .A(_19787_),
    .ZN(_19788_)
  );
  AND2_X1 _55537_ (
    .A1(_18479_),
    .A2(_19788_),
    .ZN(_19789_)
  );
  INV_X1 _55538_ (
    .A(_19789_),
    .ZN(_19790_)
  );
  AND2_X1 _55539_ (
    .A1(count_instr[27]),
    .A2(instr_rdinstr),
    .ZN(_19791_)
  );
  INV_X1 _55540_ (
    .A(_19791_),
    .ZN(_19792_)
  );
  AND2_X1 _55541_ (
    .A1(instr_rdcycleh),
    .A2(count_cycle[59]),
    .ZN(_19793_)
  );
  INV_X1 _55542_ (
    .A(_19793_),
    .ZN(_19794_)
  );
  AND2_X1 _55543_ (
    .A1(_19792_),
    .A2(_19794_),
    .ZN(_19795_)
  );
  AND2_X1 _55544_ (
    .A1(instr_rdcycle),
    .A2(count_cycle[27]),
    .ZN(_19796_)
  );
  INV_X1 _55545_ (
    .A(_19796_),
    .ZN(_19797_)
  );
  AND2_X1 _55546_ (
    .A1(count_instr[59]),
    .A2(instr_rdinstrh),
    .ZN(_19798_)
  );
  INV_X1 _55547_ (
    .A(_19798_),
    .ZN(_19799_)
  );
  AND2_X1 _55548_ (
    .A1(_19797_),
    .A2(_19799_),
    .ZN(_19800_)
  );
  AND2_X1 _55549_ (
    .A1(_19795_),
    .A2(_19800_),
    .ZN(_19801_)
  );
  INV_X1 _55550_ (
    .A(_19801_),
    .ZN(_19802_)
  );
  AND2_X1 _55551_ (
    .A1(_22271_),
    .A2(_19802_),
    .ZN(_19803_)
  );
  INV_X1 _55552_ (
    .A(_19803_),
    .ZN(_19804_)
  );
  AND2_X1 _55553_ (
    .A1(reg_op1[27]),
    .A2(_22282_),
    .ZN(_19805_)
  );
  INV_X1 _55554_ (
    .A(_19805_),
    .ZN(_19806_)
  );
  AND2_X1 _55555_ (
    .A1(_19804_),
    .A2(_19806_),
    .ZN(_19807_)
  );
  AND2_X1 _55556_ (
    .A1(_19790_),
    .A2(_19807_),
    .ZN(_19808_)
  );
  AND2_X1 _55557_ (
    .A1(_19764_),
    .A2(_19776_),
    .ZN(_19809_)
  );
  INV_X1 _55558_ (
    .A(_19809_),
    .ZN(_19810_)
  );
  AND2_X1 _55559_ (
    .A1(reg_pc[27]),
    .A2(decoded_imm[27]),
    .ZN(_19811_)
  );
  INV_X1 _55560_ (
    .A(_19811_),
    .ZN(_19812_)
  );
  AND2_X1 _55561_ (
    .A1(_21077_),
    .A2(_21982_),
    .ZN(_19813_)
  );
  INV_X1 _55562_ (
    .A(_19813_),
    .ZN(_19814_)
  );
  AND2_X1 _55563_ (
    .A1(_19812_),
    .A2(_19814_),
    .ZN(_19815_)
  );
  INV_X1 _55564_ (
    .A(_19815_),
    .ZN(_19816_)
  );
  AND2_X1 _55565_ (
    .A1(_19810_),
    .A2(_19815_),
    .ZN(_19817_)
  );
  INV_X1 _55566_ (
    .A(_19817_),
    .ZN(_19818_)
  );
  AND2_X1 _55567_ (
    .A1(_19809_),
    .A2(_19816_),
    .ZN(_19819_)
  );
  INV_X1 _55568_ (
    .A(_19819_),
    .ZN(_19820_)
  );
  AND2_X1 _55569_ (
    .A1(_19818_),
    .A2(_19820_),
    .ZN(_19821_)
  );
  AND2_X1 _55570_ (
    .A1(_11090_),
    .A2(_19821_),
    .ZN(_19822_)
  );
  INV_X1 _55571_ (
    .A(_19822_),
    .ZN(_19823_)
  );
  AND2_X1 _55572_ (
    .A1(_19808_),
    .A2(_19823_),
    .ZN(_19824_)
  );
  INV_X1 _55573_ (
    .A(_19824_),
    .ZN(_19825_)
  );
  AND2_X1 _55574_ (
    .A1(resetn),
    .A2(_19825_),
    .ZN(_00005_[27])
  );
  AND2_X1 _55575_ (
    .A1(reg_pc[28]),
    .A2(decoded_imm[28]),
    .ZN(_19826_)
  );
  INV_X1 _55576_ (
    .A(_19826_),
    .ZN(_19827_)
  );
  AND2_X1 _55577_ (
    .A1(_21076_),
    .A2(_21981_),
    .ZN(_19828_)
  );
  INV_X1 _55578_ (
    .A(_19828_),
    .ZN(_19829_)
  );
  AND2_X1 _55579_ (
    .A1(_19827_),
    .A2(_19829_),
    .ZN(_19830_)
  );
  INV_X1 _55580_ (
    .A(_19830_),
    .ZN(_19831_)
  );
  AND2_X1 _55581_ (
    .A1(_19810_),
    .A2(_19814_),
    .ZN(_19832_)
  );
  INV_X1 _55582_ (
    .A(_19832_),
    .ZN(_19833_)
  );
  AND2_X1 _55583_ (
    .A1(_19809_),
    .A2(_19812_),
    .ZN(_19834_)
  );
  INV_X1 _55584_ (
    .A(_19834_),
    .ZN(_19835_)
  );
  AND2_X1 _55585_ (
    .A1(_19812_),
    .A2(_19833_),
    .ZN(_19836_)
  );
  AND2_X1 _55586_ (
    .A1(_19814_),
    .A2(_19835_),
    .ZN(_19837_)
  );
  AND2_X1 _55587_ (
    .A1(_19830_),
    .A2(_19837_),
    .ZN(_19838_)
  );
  INV_X1 _55588_ (
    .A(_19838_),
    .ZN(_19839_)
  );
  AND2_X1 _55589_ (
    .A1(_19831_),
    .A2(_19836_),
    .ZN(_19840_)
  );
  INV_X1 _55590_ (
    .A(_19840_),
    .ZN(_19841_)
  );
  AND2_X1 _55591_ (
    .A1(latched_is_lu),
    .A2(mem_rdata[28]),
    .ZN(_19842_)
  );
  AND2_X1 _55592_ (
    .A1(_12194_),
    .A2(_19842_),
    .ZN(_19843_)
  );
  INV_X1 _55593_ (
    .A(_19843_),
    .ZN(_19844_)
  );
  AND2_X1 _55594_ (
    .A1(_19313_),
    .A2(_19844_),
    .ZN(_19845_)
  );
  INV_X1 _55595_ (
    .A(_19845_),
    .ZN(_19846_)
  );
  AND2_X1 _55596_ (
    .A1(_18479_),
    .A2(_19846_),
    .ZN(_19847_)
  );
  INV_X1 _55597_ (
    .A(_19847_),
    .ZN(_19848_)
  );
  AND2_X1 _55598_ (
    .A1(count_instr[28]),
    .A2(instr_rdinstr),
    .ZN(_19849_)
  );
  INV_X1 _55599_ (
    .A(_19849_),
    .ZN(_19850_)
  );
  AND2_X1 _55600_ (
    .A1(instr_rdcycleh),
    .A2(count_cycle[60]),
    .ZN(_19851_)
  );
  INV_X1 _55601_ (
    .A(_19851_),
    .ZN(_19852_)
  );
  AND2_X1 _55602_ (
    .A1(_19850_),
    .A2(_19852_),
    .ZN(_19853_)
  );
  AND2_X1 _55603_ (
    .A1(count_instr[60]),
    .A2(instr_rdinstrh),
    .ZN(_19854_)
  );
  INV_X1 _55604_ (
    .A(_19854_),
    .ZN(_19855_)
  );
  AND2_X1 _55605_ (
    .A1(instr_rdcycle),
    .A2(count_cycle[28]),
    .ZN(_19856_)
  );
  INV_X1 _55606_ (
    .A(_19856_),
    .ZN(_19857_)
  );
  AND2_X1 _55607_ (
    .A1(_19855_),
    .A2(_19857_),
    .ZN(_19858_)
  );
  AND2_X1 _55608_ (
    .A1(_19853_),
    .A2(_19858_),
    .ZN(_19859_)
  );
  INV_X1 _55609_ (
    .A(_19859_),
    .ZN(_19860_)
  );
  AND2_X1 _55610_ (
    .A1(_22271_),
    .A2(_19860_),
    .ZN(_19861_)
  );
  INV_X1 _55611_ (
    .A(_19861_),
    .ZN(_19862_)
  );
  AND2_X1 _55612_ (
    .A1(reg_op1[28]),
    .A2(_22282_),
    .ZN(_19863_)
  );
  INV_X1 _55613_ (
    .A(_19863_),
    .ZN(_19864_)
  );
  AND2_X1 _55614_ (
    .A1(_19862_),
    .A2(_19864_),
    .ZN(_19865_)
  );
  AND2_X1 _55615_ (
    .A1(_11090_),
    .A2(_19839_),
    .ZN(_19866_)
  );
  AND2_X1 _55616_ (
    .A1(_19841_),
    .A2(_19866_),
    .ZN(_19867_)
  );
  INV_X1 _55617_ (
    .A(_19867_),
    .ZN(_19868_)
  );
  AND2_X1 _55618_ (
    .A1(_19865_),
    .A2(_19868_),
    .ZN(_19869_)
  );
  AND2_X1 _55619_ (
    .A1(_19848_),
    .A2(_19869_),
    .ZN(_19870_)
  );
  INV_X1 _55620_ (
    .A(_19870_),
    .ZN(_19871_)
  );
  AND2_X1 _55621_ (
    .A1(resetn),
    .A2(_19871_),
    .ZN(_00005_[28])
  );
  AND2_X1 _55622_ (
    .A1(_19827_),
    .A2(_19839_),
    .ZN(_19872_)
  );
  INV_X1 _55623_ (
    .A(_19872_),
    .ZN(_19873_)
  );
  AND2_X1 _55624_ (
    .A1(reg_pc[29]),
    .A2(decoded_imm[29]),
    .ZN(_19874_)
  );
  INV_X1 _55625_ (
    .A(_19874_),
    .ZN(_19875_)
  );
  AND2_X1 _55626_ (
    .A1(_21075_),
    .A2(_21980_),
    .ZN(_19876_)
  );
  INV_X1 _55627_ (
    .A(_19876_),
    .ZN(_19877_)
  );
  AND2_X1 _55628_ (
    .A1(_19875_),
    .A2(_19877_),
    .ZN(_19878_)
  );
  INV_X1 _55629_ (
    .A(_19878_),
    .ZN(_19879_)
  );
  AND2_X1 _55630_ (
    .A1(_19873_),
    .A2(_19878_),
    .ZN(_19880_)
  );
  INV_X1 _55631_ (
    .A(_19880_),
    .ZN(_19881_)
  );
  AND2_X1 _55632_ (
    .A1(_19872_),
    .A2(_19879_),
    .ZN(_19882_)
  );
  INV_X1 _55633_ (
    .A(_19882_),
    .ZN(_19883_)
  );
  AND2_X1 _55634_ (
    .A1(_11090_),
    .A2(_19883_),
    .ZN(_19884_)
  );
  AND2_X1 _55635_ (
    .A1(_19881_),
    .A2(_19884_),
    .ZN(_19885_)
  );
  INV_X1 _55636_ (
    .A(_19885_),
    .ZN(_19886_)
  );
  AND2_X1 _55637_ (
    .A1(latched_is_lu),
    .A2(mem_rdata[29]),
    .ZN(_19887_)
  );
  AND2_X1 _55638_ (
    .A1(_12194_),
    .A2(_19887_),
    .ZN(_19888_)
  );
  INV_X1 _55639_ (
    .A(_19888_),
    .ZN(_19889_)
  );
  AND2_X1 _55640_ (
    .A1(_19313_),
    .A2(_19889_),
    .ZN(_19890_)
  );
  INV_X1 _55641_ (
    .A(_19890_),
    .ZN(_19891_)
  );
  AND2_X1 _55642_ (
    .A1(_18479_),
    .A2(_19891_),
    .ZN(_19892_)
  );
  INV_X1 _55643_ (
    .A(_19892_),
    .ZN(_19893_)
  );
  AND2_X1 _55644_ (
    .A1(count_instr[29]),
    .A2(instr_rdinstr),
    .ZN(_19894_)
  );
  INV_X1 _55645_ (
    .A(_19894_),
    .ZN(_19895_)
  );
  AND2_X1 _55646_ (
    .A1(instr_rdcycleh),
    .A2(count_cycle[61]),
    .ZN(_19896_)
  );
  INV_X1 _55647_ (
    .A(_19896_),
    .ZN(_19897_)
  );
  AND2_X1 _55648_ (
    .A1(_19895_),
    .A2(_19897_),
    .ZN(_19898_)
  );
  AND2_X1 _55649_ (
    .A1(count_instr[61]),
    .A2(instr_rdinstrh),
    .ZN(_19899_)
  );
  INV_X1 _55650_ (
    .A(_19899_),
    .ZN(_19900_)
  );
  AND2_X1 _55651_ (
    .A1(instr_rdcycle),
    .A2(count_cycle[29]),
    .ZN(_19901_)
  );
  INV_X1 _55652_ (
    .A(_19901_),
    .ZN(_19902_)
  );
  AND2_X1 _55653_ (
    .A1(_19900_),
    .A2(_19902_),
    .ZN(_19903_)
  );
  AND2_X1 _55654_ (
    .A1(_19898_),
    .A2(_19903_),
    .ZN(_19904_)
  );
  INV_X1 _55655_ (
    .A(_19904_),
    .ZN(_19905_)
  );
  AND2_X1 _55656_ (
    .A1(_22271_),
    .A2(_19905_),
    .ZN(_19906_)
  );
  INV_X1 _55657_ (
    .A(_19906_),
    .ZN(_19907_)
  );
  AND2_X1 _55658_ (
    .A1(reg_op1[29]),
    .A2(_22282_),
    .ZN(_19908_)
  );
  INV_X1 _55659_ (
    .A(_19908_),
    .ZN(_19909_)
  );
  AND2_X1 _55660_ (
    .A1(_19907_),
    .A2(_19909_),
    .ZN(_19910_)
  );
  AND2_X1 _55661_ (
    .A1(_19893_),
    .A2(_19910_),
    .ZN(_19911_)
  );
  AND2_X1 _55662_ (
    .A1(_19886_),
    .A2(_19911_),
    .ZN(_19912_)
  );
  INV_X1 _55663_ (
    .A(_19912_),
    .ZN(_19913_)
  );
  AND2_X1 _55664_ (
    .A1(resetn),
    .A2(_19913_),
    .ZN(_00005_[29])
  );
  AND2_X1 _55665_ (
    .A1(latched_is_lu),
    .A2(mem_rdata[30]),
    .ZN(_19914_)
  );
  AND2_X1 _55666_ (
    .A1(_12194_),
    .A2(_19914_),
    .ZN(_19915_)
  );
  INV_X1 _55667_ (
    .A(_19915_),
    .ZN(_19916_)
  );
  AND2_X1 _55668_ (
    .A1(_19313_),
    .A2(_19916_),
    .ZN(_19917_)
  );
  INV_X1 _55669_ (
    .A(_19917_),
    .ZN(_19918_)
  );
  AND2_X1 _55670_ (
    .A1(_18479_),
    .A2(_19918_),
    .ZN(_19919_)
  );
  INV_X1 _55671_ (
    .A(_19919_),
    .ZN(_19920_)
  );
  AND2_X1 _55672_ (
    .A1(reg_op1[30]),
    .A2(_22282_),
    .ZN(_19921_)
  );
  INV_X1 _55673_ (
    .A(_19921_),
    .ZN(_19922_)
  );
  AND2_X1 _55674_ (
    .A1(count_instr[62]),
    .A2(instr_rdinstrh),
    .ZN(_19923_)
  );
  INV_X1 _55675_ (
    .A(_19923_),
    .ZN(_19924_)
  );
  AND2_X1 _55676_ (
    .A1(count_instr[30]),
    .A2(instr_rdinstr),
    .ZN(_19925_)
  );
  INV_X1 _55677_ (
    .A(_19925_),
    .ZN(_19926_)
  );
  AND2_X1 _55678_ (
    .A1(_19924_),
    .A2(_19926_),
    .ZN(_19927_)
  );
  AND2_X1 _55679_ (
    .A1(instr_rdcycle),
    .A2(count_cycle[30]),
    .ZN(_19928_)
  );
  INV_X1 _55680_ (
    .A(_19928_),
    .ZN(_19929_)
  );
  AND2_X1 _55681_ (
    .A1(instr_rdcycleh),
    .A2(count_cycle[62]),
    .ZN(_19930_)
  );
  INV_X1 _55682_ (
    .A(_19930_),
    .ZN(_19931_)
  );
  AND2_X1 _55683_ (
    .A1(_19929_),
    .A2(_19931_),
    .ZN(_19932_)
  );
  AND2_X1 _55684_ (
    .A1(_19927_),
    .A2(_19932_),
    .ZN(_19933_)
  );
  INV_X1 _55685_ (
    .A(_19933_),
    .ZN(_19934_)
  );
  AND2_X1 _55686_ (
    .A1(_22271_),
    .A2(_19934_),
    .ZN(_19935_)
  );
  INV_X1 _55687_ (
    .A(_19935_),
    .ZN(_19936_)
  );
  AND2_X1 _55688_ (
    .A1(_19922_),
    .A2(_19936_),
    .ZN(_19937_)
  );
  AND2_X1 _55689_ (
    .A1(_19875_),
    .A2(_19881_),
    .ZN(_19938_)
  );
  INV_X1 _55690_ (
    .A(_19938_),
    .ZN(_19939_)
  );
  AND2_X1 _55691_ (
    .A1(reg_pc[30]),
    .A2(decoded_imm[30]),
    .ZN(_19940_)
  );
  INV_X1 _55692_ (
    .A(_19940_),
    .ZN(_19941_)
  );
  AND2_X1 _55693_ (
    .A1(_21074_),
    .A2(_21979_),
    .ZN(_19942_)
  );
  INV_X1 _55694_ (
    .A(_19942_),
    .ZN(_19943_)
  );
  AND2_X1 _55695_ (
    .A1(_19941_),
    .A2(_19943_),
    .ZN(_19944_)
  );
  INV_X1 _55696_ (
    .A(_19944_),
    .ZN(_19945_)
  );
  AND2_X1 _55697_ (
    .A1(_19938_),
    .A2(_19945_),
    .ZN(_19946_)
  );
  INV_X1 _55698_ (
    .A(_19946_),
    .ZN(_19947_)
  );
  AND2_X1 _55699_ (
    .A1(_19939_),
    .A2(_19944_),
    .ZN(_19948_)
  );
  INV_X1 _55700_ (
    .A(_19948_),
    .ZN(_19949_)
  );
  AND2_X1 _55701_ (
    .A1(_11090_),
    .A2(_19949_),
    .ZN(_19950_)
  );
  AND2_X1 _55702_ (
    .A1(_19947_),
    .A2(_19950_),
    .ZN(_19951_)
  );
  INV_X1 _55703_ (
    .A(_19951_),
    .ZN(_19952_)
  );
  AND2_X1 _55704_ (
    .A1(_19937_),
    .A2(_19952_),
    .ZN(_19953_)
  );
  AND2_X1 _55705_ (
    .A1(_19920_),
    .A2(_19953_),
    .ZN(_19954_)
  );
  INV_X1 _55706_ (
    .A(_19954_),
    .ZN(_19955_)
  );
  AND2_X1 _55707_ (
    .A1(resetn),
    .A2(_19955_),
    .ZN(_00005_[30])
  );
  AND2_X1 _55708_ (
    .A1(latched_is_lu),
    .A2(mem_rdata[31]),
    .ZN(_19956_)
  );
  AND2_X1 _55709_ (
    .A1(_12194_),
    .A2(_19956_),
    .ZN(_19957_)
  );
  INV_X1 _55710_ (
    .A(_19957_),
    .ZN(_19958_)
  );
  AND2_X1 _55711_ (
    .A1(_19313_),
    .A2(_19958_),
    .ZN(_19959_)
  );
  INV_X1 _55712_ (
    .A(_19959_),
    .ZN(_19960_)
  );
  AND2_X1 _55713_ (
    .A1(_18479_),
    .A2(_19960_),
    .ZN(_19961_)
  );
  INV_X1 _55714_ (
    .A(_19961_),
    .ZN(_19962_)
  );
  AND2_X1 _55715_ (
    .A1(count_instr[31]),
    .A2(instr_rdinstr),
    .ZN(_19963_)
  );
  INV_X1 _55716_ (
    .A(_19963_),
    .ZN(_19964_)
  );
  AND2_X1 _55717_ (
    .A1(instr_rdcycleh),
    .A2(count_cycle[63]),
    .ZN(_19965_)
  );
  INV_X1 _55718_ (
    .A(_19965_),
    .ZN(_19966_)
  );
  AND2_X1 _55719_ (
    .A1(_19964_),
    .A2(_19966_),
    .ZN(_19967_)
  );
  AND2_X1 _55720_ (
    .A1(count_instr[63]),
    .A2(instr_rdinstrh),
    .ZN(_19968_)
  );
  INV_X1 _55721_ (
    .A(_19968_),
    .ZN(_19969_)
  );
  AND2_X1 _55722_ (
    .A1(instr_rdcycle),
    .A2(count_cycle[31]),
    .ZN(_19970_)
  );
  INV_X1 _55723_ (
    .A(_19970_),
    .ZN(_19971_)
  );
  AND2_X1 _55724_ (
    .A1(_19969_),
    .A2(_19971_),
    .ZN(_19972_)
  );
  AND2_X1 _55725_ (
    .A1(_19967_),
    .A2(_19972_),
    .ZN(_19973_)
  );
  INV_X1 _55726_ (
    .A(_19973_),
    .ZN(_19974_)
  );
  AND2_X1 _55727_ (
    .A1(_22271_),
    .A2(_19974_),
    .ZN(_19975_)
  );
  INV_X1 _55728_ (
    .A(_19975_),
    .ZN(_19976_)
  );
  AND2_X1 _55729_ (
    .A1(reg_op1[31]),
    .A2(_22282_),
    .ZN(_19977_)
  );
  INV_X1 _55730_ (
    .A(_19977_),
    .ZN(_19978_)
  );
  AND2_X1 _55731_ (
    .A1(_19976_),
    .A2(_19978_),
    .ZN(_19979_)
  );
  AND2_X1 _55732_ (
    .A1(_19962_),
    .A2(_19979_),
    .ZN(_19980_)
  );
  INV_X1 _55733_ (
    .A(_19980_),
    .ZN(_19981_)
  );
  AND2_X1 _55734_ (
    .A1(resetn),
    .A2(_19981_),
    .ZN(_19982_)
  );
  INV_X1 _55735_ (
    .A(_19982_),
    .ZN(_19983_)
  );
  AND2_X1 _55736_ (
    .A1(_19941_),
    .A2(_19949_),
    .ZN(_19984_)
  );
  INV_X1 _55737_ (
    .A(_19984_),
    .ZN(_19985_)
  );
  AND2_X1 _55738_ (
    .A1(reg_pc[31]),
    .A2(_21978_),
    .ZN(_19986_)
  );
  INV_X1 _55739_ (
    .A(_19986_),
    .ZN(_19987_)
  );
  AND2_X1 _55740_ (
    .A1(_21073_),
    .A2(decoded_imm[31]),
    .ZN(_19988_)
  );
  INV_X1 _55741_ (
    .A(_19988_),
    .ZN(_19989_)
  );
  AND2_X1 _55742_ (
    .A1(_21073_),
    .A2(_21978_),
    .ZN(_19990_)
  );
  INV_X1 _55743_ (
    .A(_19990_),
    .ZN(_19991_)
  );
  AND2_X1 _55744_ (
    .A1(reg_pc[31]),
    .A2(decoded_imm[31]),
    .ZN(_19992_)
  );
  INV_X1 _55745_ (
    .A(_19992_),
    .ZN(_19993_)
  );
  AND2_X1 _55746_ (
    .A1(_19987_),
    .A2(_19989_),
    .ZN(_19994_)
  );
  AND2_X1 _55747_ (
    .A1(_19991_),
    .A2(_19993_),
    .ZN(_19995_)
  );
  AND2_X1 _55748_ (
    .A1(_19984_),
    .A2(_19994_),
    .ZN(_19996_)
  );
  INV_X1 _55749_ (
    .A(_19996_),
    .ZN(_19997_)
  );
  AND2_X1 _55750_ (
    .A1(_19985_),
    .A2(_19995_),
    .ZN(_19998_)
  );
  INV_X1 _55751_ (
    .A(_19998_),
    .ZN(_19999_)
  );
  AND2_X1 _55752_ (
    .A1(_19997_),
    .A2(_19999_),
    .ZN(_20000_)
  );
  AND2_X1 _55753_ (
    .A1(_11098_),
    .A2(_20000_),
    .ZN(_20001_)
  );
  INV_X1 _55754_ (
    .A(_20001_),
    .ZN(_20002_)
  );
  AND2_X1 _55755_ (
    .A1(_19983_),
    .A2(_20002_),
    .ZN(_20003_)
  );
  INV_X1 _55756_ (
    .A(_20003_),
    .ZN(_00005_[31])
  );
  AND2_X1 _55757_ (
    .A1(decoded_rs2[0]),
    .A2(_18235_),
    .ZN(_20004_)
  );
  INV_X1 _55758_ (
    .A(_20004_),
    .ZN(_20005_)
  );
  AND2_X1 _55759_ (
    .A1(_29149_[0]),
    .A2(_22572_),
    .ZN(_20006_)
  );
  INV_X1 _55760_ (
    .A(_20006_),
    .ZN(_20007_)
  );
  AND2_X1 _55761_ (
    .A1(reg_sh[0]),
    .A2(_22573_),
    .ZN(_20008_)
  );
  INV_X1 _55762_ (
    .A(_20008_),
    .ZN(_20009_)
  );
  AND2_X1 _55763_ (
    .A1(_20007_),
    .A2(_20009_),
    .ZN(_20010_)
  );
  INV_X1 _55764_ (
    .A(_20010_),
    .ZN(_20011_)
  );
  AND2_X1 _55765_ (
    .A1(_22295_),
    .A2(_20011_),
    .ZN(_20012_)
  );
  INV_X1 _55766_ (
    .A(_20012_),
    .ZN(_20013_)
  );
  AND2_X1 _55767_ (
    .A1(_20005_),
    .A2(_20013_),
    .ZN(_20014_)
  );
  AND2_X1 _55768_ (
    .A1(_05141_),
    .A2(_20014_),
    .ZN(_20015_)
  );
  INV_X1 _55769_ (
    .A(_20015_),
    .ZN(_20016_)
  );
  AND2_X1 _55770_ (
    .A1(resetn),
    .A2(_20016_),
    .ZN(_00006_[0])
  );
  AND2_X1 _55771_ (
    .A1(decoded_rs2[1]),
    .A2(_18235_),
    .ZN(_20017_)
  );
  INV_X1 _55772_ (
    .A(_20017_),
    .ZN(_20018_)
  );
  AND2_X1 _55773_ (
    .A1(reg_sh[0]),
    .A2(_29149_[1]),
    .ZN(_20019_)
  );
  INV_X1 _55774_ (
    .A(_20019_),
    .ZN(_20020_)
  );
  AND2_X1 _55775_ (
    .A1(_22036_),
    .A2(_22068_),
    .ZN(_20021_)
  );
  INV_X1 _55776_ (
    .A(_20021_),
    .ZN(_20022_)
  );
  AND2_X1 _55777_ (
    .A1(_20020_),
    .A2(_20022_),
    .ZN(_20023_)
  );
  AND2_X1 _55778_ (
    .A1(_22572_),
    .A2(_20023_),
    .ZN(_20024_)
  );
  INV_X1 _55779_ (
    .A(_20024_),
    .ZN(_20025_)
  );
  AND2_X1 _55780_ (
    .A1(reg_sh[1]),
    .A2(_22573_),
    .ZN(_20026_)
  );
  INV_X1 _55781_ (
    .A(_20026_),
    .ZN(_20027_)
  );
  AND2_X1 _55782_ (
    .A1(_20025_),
    .A2(_20027_),
    .ZN(_20028_)
  );
  INV_X1 _55783_ (
    .A(_20028_),
    .ZN(_20029_)
  );
  AND2_X1 _55784_ (
    .A1(_22295_),
    .A2(_20029_),
    .ZN(_20030_)
  );
  INV_X1 _55785_ (
    .A(_20030_),
    .ZN(_20031_)
  );
  AND2_X1 _55786_ (
    .A1(_20018_),
    .A2(_20031_),
    .ZN(_20032_)
  );
  AND2_X1 _55787_ (
    .A1(_05312_),
    .A2(_20032_),
    .ZN(_20033_)
  );
  INV_X1 _55788_ (
    .A(_20033_),
    .ZN(_20034_)
  );
  AND2_X1 _55789_ (
    .A1(resetn),
    .A2(_20034_),
    .ZN(_00006_[1])
  );
  AND2_X1 _55790_ (
    .A1(decoded_rs2[2]),
    .A2(_18235_),
    .ZN(_20035_)
  );
  INV_X1 _55791_ (
    .A(_20035_),
    .ZN(_20036_)
  );
  AND2_X1 _55792_ (
    .A1(_22030_),
    .A2(_20020_),
    .ZN(_20037_)
  );
  INV_X1 _55793_ (
    .A(_20037_),
    .ZN(_20038_)
  );
  AND2_X1 _55794_ (
    .A1(_22572_),
    .A2(_20038_),
    .ZN(_20039_)
  );
  INV_X1 _55795_ (
    .A(_20039_),
    .ZN(_20040_)
  );
  AND2_X1 _55796_ (
    .A1(_29150_[2]),
    .A2(_20039_),
    .ZN(_20041_)
  );
  INV_X1 _55797_ (
    .A(_20041_),
    .ZN(_20042_)
  );
  AND2_X1 _55798_ (
    .A1(_22145_),
    .A2(_20040_),
    .ZN(_20043_)
  );
  INV_X1 _55799_ (
    .A(_20043_),
    .ZN(_20044_)
  );
  AND2_X1 _55800_ (
    .A1(_22295_),
    .A2(_20044_),
    .ZN(_20045_)
  );
  AND2_X1 _55801_ (
    .A1(_20042_),
    .A2(_20045_),
    .ZN(_20046_)
  );
  INV_X1 _55802_ (
    .A(_20046_),
    .ZN(_20047_)
  );
  AND2_X1 _55803_ (
    .A1(_20036_),
    .A2(_20047_),
    .ZN(_20048_)
  );
  AND2_X1 _55804_ (
    .A1(_05483_),
    .A2(_20048_),
    .ZN(_20049_)
  );
  INV_X1 _55805_ (
    .A(_20049_),
    .ZN(_20050_)
  );
  AND2_X1 _55806_ (
    .A1(resetn),
    .A2(_20050_),
    .ZN(_00006_[2])
  );
  AND2_X1 _55807_ (
    .A1(decoded_rs2[3]),
    .A2(_18235_),
    .ZN(_20051_)
  );
  INV_X1 _55808_ (
    .A(_20051_),
    .ZN(_20052_)
  );
  AND2_X1 _55809_ (
    .A1(_22037_),
    .A2(_20042_),
    .ZN(_20053_)
  );
  INV_X1 _55810_ (
    .A(_20053_),
    .ZN(_20054_)
  );
  AND2_X1 _55811_ (
    .A1(_22217_),
    .A2(_20053_),
    .ZN(_20055_)
  );
  INV_X1 _55812_ (
    .A(_20055_),
    .ZN(_20056_)
  );
  AND2_X1 _55813_ (
    .A1(_29149_[3]),
    .A2(_20054_),
    .ZN(_20057_)
  );
  INV_X1 _55814_ (
    .A(_20057_),
    .ZN(_20058_)
  );
  AND2_X1 _55815_ (
    .A1(_22295_),
    .A2(_20058_),
    .ZN(_20059_)
  );
  AND2_X1 _55816_ (
    .A1(_20056_),
    .A2(_20059_),
    .ZN(_20060_)
  );
  INV_X1 _55817_ (
    .A(_20060_),
    .ZN(_20061_)
  );
  AND2_X1 _55818_ (
    .A1(_20052_),
    .A2(_20061_),
    .ZN(_20062_)
  );
  AND2_X1 _55819_ (
    .A1(_05659_),
    .A2(_20062_),
    .ZN(_20063_)
  );
  INV_X1 _55820_ (
    .A(_20063_),
    .ZN(_20064_)
  );
  AND2_X1 _55821_ (
    .A1(resetn),
    .A2(_20064_),
    .ZN(_00006_[3])
  );
  AND2_X1 _55822_ (
    .A1(_22029_),
    .A2(_20058_),
    .ZN(_20065_)
  );
  INV_X1 _55823_ (
    .A(_20065_),
    .ZN(_20066_)
  );
  AND2_X1 _55824_ (
    .A1(_22069_),
    .A2(_20066_),
    .ZN(_20067_)
  );
  INV_X1 _55825_ (
    .A(_20067_),
    .ZN(_20068_)
  );
  AND2_X1 _55826_ (
    .A1(_29149_[4]),
    .A2(_20065_),
    .ZN(_20069_)
  );
  INV_X1 _55827_ (
    .A(_20069_),
    .ZN(_20070_)
  );
  AND2_X1 _55828_ (
    .A1(_20068_),
    .A2(_20070_),
    .ZN(_20071_)
  );
  INV_X1 _55829_ (
    .A(_20071_),
    .ZN(_20072_)
  );
  AND2_X1 _55830_ (
    .A1(_22295_),
    .A2(_20072_),
    .ZN(_20073_)
  );
  INV_X1 _55831_ (
    .A(_20073_),
    .ZN(_20074_)
  );
  AND2_X1 _55832_ (
    .A1(decoded_imm_j[4]),
    .A2(_18235_),
    .ZN(_20075_)
  );
  INV_X1 _55833_ (
    .A(_20075_),
    .ZN(_20076_)
  );
  AND2_X1 _55834_ (
    .A1(_20074_),
    .A2(_20076_),
    .ZN(_20077_)
  );
  AND2_X1 _55835_ (
    .A1(_05832_),
    .A2(_20077_),
    .ZN(_20078_)
  );
  INV_X1 _55836_ (
    .A(_20078_),
    .ZN(_20079_)
  );
  AND2_X1 _55837_ (
    .A1(resetn),
    .A2(_20079_),
    .ZN(_00006_[4])
  );
  AND2_X1 _55838_ (
    .A1(is_compare),
    .A2(_11087_),
    .ZN(_20080_)
  );
  INV_X1 _55839_ (
    .A(_20080_),
    .ZN(_20081_)
  );
  AND2_X1 _55840_ (
    .A1(_21049_),
    .A2(is_lui_auipc_jal_jalr_addi_add_sub),
    .ZN(_20082_)
  );
  INV_X1 _55841_ (
    .A(_20082_),
    .ZN(_20083_)
  );
  AND2_X1 _55842_ (
    .A1(_22527_),
    .A2(_20083_),
    .ZN(_20084_)
  );
  INV_X1 _55843_ (
    .A(_20084_),
    .ZN(_20085_)
  );
  AND2_X1 _55844_ (
    .A1(_10975_),
    .A2(_20085_),
    .ZN(_20086_)
  );
  INV_X1 _55845_ (
    .A(_20086_),
    .ZN(_20087_)
  );
  AND2_X1 _55846_ (
    .A1(reg_op1[0]),
    .A2(_29151_[0]),
    .ZN(_20088_)
  );
  INV_X1 _55847_ (
    .A(_20088_),
    .ZN(_20089_)
  );
  AND2_X1 _55848_ (
    .A1(_10674_),
    .A2(_20089_),
    .ZN(_20090_)
  );
  INV_X1 _55849_ (
    .A(_20090_),
    .ZN(_20091_)
  );
  AND2_X1 _55850_ (
    .A1(instr_sub),
    .A2(is_lui_auipc_jal_jalr_addi_add_sub),
    .ZN(_20092_)
  );
  INV_X1 _55851_ (
    .A(_20092_),
    .ZN(_20093_)
  );
  AND2_X1 _55852_ (
    .A1(_20091_),
    .A2(_20092_),
    .ZN(_20094_)
  );
  INV_X1 _55853_ (
    .A(_20094_),
    .ZN(_20095_)
  );
  AND2_X1 _55854_ (
    .A1(_21041_),
    .A2(_21051_),
    .ZN(_20096_)
  );
  INV_X1 _55855_ (
    .A(_20096_),
    .ZN(_20097_)
  );
  AND2_X1 _55856_ (
    .A1(_10971_),
    .A2(_20097_),
    .ZN(_20098_)
  );
  INV_X1 _55857_ (
    .A(_20098_),
    .ZN(_20099_)
  );
  AND2_X1 _55858_ (
    .A1(_22532_),
    .A2(_10974_),
    .ZN(_20100_)
  );
  INV_X1 _55859_ (
    .A(_20100_),
    .ZN(_20101_)
  );
  AND2_X1 _55860_ (
    .A1(_20099_),
    .A2(_20101_),
    .ZN(_20102_)
  );
  AND2_X1 _55861_ (
    .A1(_20095_),
    .A2(_20102_),
    .ZN(_20103_)
  );
  AND2_X1 _55862_ (
    .A1(_20087_),
    .A2(_20103_),
    .ZN(_20104_)
  );
  AND2_X1 _55863_ (
    .A1(_20081_),
    .A2(_20104_),
    .ZN(_20105_)
  );
  INV_X1 _55864_ (
    .A(_20105_),
    .ZN(alu_out[0])
  );
  AND2_X1 _55865_ (
    .A1(_10673_),
    .A2(_10678_),
    .ZN(_20106_)
  );
  INV_X1 _55866_ (
    .A(_20106_),
    .ZN(_20107_)
  );
  AND2_X1 _55867_ (
    .A1(instr_sub),
    .A2(_10680_),
    .ZN(_20108_)
  );
  AND2_X1 _55868_ (
    .A1(_20107_),
    .A2(_20108_),
    .ZN(_20109_)
  );
  INV_X1 _55869_ (
    .A(_20109_),
    .ZN(_20110_)
  );
  AND2_X1 _55870_ (
    .A1(_10855_),
    .A2(_10971_),
    .ZN(_20111_)
  );
  INV_X1 _55871_ (
    .A(_20111_),
    .ZN(_20112_)
  );
  AND2_X1 _55872_ (
    .A1(_10856_),
    .A2(_10972_),
    .ZN(_20113_)
  );
  INV_X1 _55873_ (
    .A(_20113_),
    .ZN(_20114_)
  );
  AND2_X1 _55874_ (
    .A1(_21049_),
    .A2(_20112_),
    .ZN(_20115_)
  );
  AND2_X1 _55875_ (
    .A1(_20114_),
    .A2(_20115_),
    .ZN(_20116_)
  );
  INV_X1 _55876_ (
    .A(_20116_),
    .ZN(_20117_)
  );
  AND2_X1 _55877_ (
    .A1(_20110_),
    .A2(_20117_),
    .ZN(_20118_)
  );
  INV_X1 _55878_ (
    .A(_20118_),
    .ZN(_20119_)
  );
  AND2_X1 _55879_ (
    .A1(is_lui_auipc_jal_jalr_addi_add_sub),
    .A2(_20119_),
    .ZN(_20120_)
  );
  INV_X1 _55880_ (
    .A(_20120_),
    .ZN(_20121_)
  );
  AND2_X1 _55881_ (
    .A1(_22528_),
    .A2(_10855_),
    .ZN(_20122_)
  );
  INV_X1 _55882_ (
    .A(_20122_),
    .ZN(_20123_)
  );
  AND2_X1 _55883_ (
    .A1(_10851_),
    .A2(_20097_),
    .ZN(_20124_)
  );
  INV_X1 _55884_ (
    .A(_20124_),
    .ZN(_20125_)
  );
  AND2_X1 _55885_ (
    .A1(_22532_),
    .A2(_10854_),
    .ZN(_20126_)
  );
  INV_X1 _55886_ (
    .A(_20126_),
    .ZN(_20127_)
  );
  AND2_X1 _55887_ (
    .A1(_20125_),
    .A2(_20127_),
    .ZN(_20128_)
  );
  AND2_X1 _55888_ (
    .A1(_20123_),
    .A2(_20128_),
    .ZN(_20129_)
  );
  AND2_X1 _55889_ (
    .A1(_20121_),
    .A2(_20129_),
    .ZN(_20130_)
  );
  INV_X1 _55890_ (
    .A(_20130_),
    .ZN(alu_out[1])
  );
  AND2_X1 _55891_ (
    .A1(_10681_),
    .A2(_10686_),
    .ZN(_20131_)
  );
  INV_X1 _55892_ (
    .A(_20131_),
    .ZN(_20132_)
  );
  AND2_X1 _55893_ (
    .A1(instr_sub),
    .A2(_10688_),
    .ZN(_20133_)
  );
  AND2_X1 _55894_ (
    .A1(_20132_),
    .A2(_20133_),
    .ZN(_20134_)
  );
  INV_X1 _55895_ (
    .A(_20134_),
    .ZN(_20135_)
  );
  AND2_X1 _55896_ (
    .A1(_10852_),
    .A2(_20112_),
    .ZN(_20136_)
  );
  INV_X1 _55897_ (
    .A(_20136_),
    .ZN(_20137_)
  );
  AND2_X1 _55898_ (
    .A1(_11035_),
    .A2(_20137_),
    .ZN(_20138_)
  );
  INV_X1 _55899_ (
    .A(_20138_),
    .ZN(_20139_)
  );
  AND2_X1 _55900_ (
    .A1(_11036_),
    .A2(_20136_),
    .ZN(_20140_)
  );
  INV_X1 _55901_ (
    .A(_20140_),
    .ZN(_20141_)
  );
  AND2_X1 _55902_ (
    .A1(_21049_),
    .A2(_20141_),
    .ZN(_20142_)
  );
  AND2_X1 _55903_ (
    .A1(_20139_),
    .A2(_20142_),
    .ZN(_20143_)
  );
  INV_X1 _55904_ (
    .A(_20143_),
    .ZN(_20144_)
  );
  AND2_X1 _55905_ (
    .A1(_20135_),
    .A2(_20144_),
    .ZN(_20145_)
  );
  INV_X1 _55906_ (
    .A(_20145_),
    .ZN(_20146_)
  );
  AND2_X1 _55907_ (
    .A1(is_lui_auipc_jal_jalr_addi_add_sub),
    .A2(_20146_),
    .ZN(_20147_)
  );
  INV_X1 _55908_ (
    .A(_20147_),
    .ZN(_20148_)
  );
  AND2_X1 _55909_ (
    .A1(_22528_),
    .A2(_11035_),
    .ZN(_20149_)
  );
  INV_X1 _55910_ (
    .A(_20149_),
    .ZN(_20150_)
  );
  AND2_X1 _55911_ (
    .A1(_11031_),
    .A2(_20097_),
    .ZN(_20151_)
  );
  INV_X1 _55912_ (
    .A(_20151_),
    .ZN(_20152_)
  );
  AND2_X1 _55913_ (
    .A1(_22532_),
    .A2(_11034_),
    .ZN(_20153_)
  );
  INV_X1 _55914_ (
    .A(_20153_),
    .ZN(_20154_)
  );
  AND2_X1 _55915_ (
    .A1(_20152_),
    .A2(_20154_),
    .ZN(_20155_)
  );
  AND2_X1 _55916_ (
    .A1(_20150_),
    .A2(_20155_),
    .ZN(_20156_)
  );
  AND2_X1 _55917_ (
    .A1(_20148_),
    .A2(_20156_),
    .ZN(_20157_)
  );
  INV_X1 _55918_ (
    .A(_20157_),
    .ZN(alu_out[2])
  );
  AND2_X1 _55919_ (
    .A1(_11032_),
    .A2(_20139_),
    .ZN(_20158_)
  );
  INV_X1 _55920_ (
    .A(_20158_),
    .ZN(_20159_)
  );
  AND2_X1 _55921_ (
    .A1(_10927_),
    .A2(_20159_),
    .ZN(_20160_)
  );
  INV_X1 _55922_ (
    .A(_20160_),
    .ZN(_20161_)
  );
  AND2_X1 _55923_ (
    .A1(_10928_),
    .A2(_20158_),
    .ZN(_20162_)
  );
  INV_X1 _55924_ (
    .A(_20162_),
    .ZN(_20163_)
  );
  AND2_X1 _55925_ (
    .A1(_21049_),
    .A2(_20163_),
    .ZN(_20164_)
  );
  AND2_X1 _55926_ (
    .A1(_20161_),
    .A2(_20164_),
    .ZN(_20165_)
  );
  INV_X1 _55927_ (
    .A(_20165_),
    .ZN(_20166_)
  );
  AND2_X1 _55928_ (
    .A1(_10666_),
    .A2(_10668_),
    .ZN(_20167_)
  );
  INV_X1 _55929_ (
    .A(_20167_),
    .ZN(_20168_)
  );
  AND2_X1 _55930_ (
    .A1(_10689_),
    .A2(_20168_),
    .ZN(_20169_)
  );
  INV_X1 _55931_ (
    .A(_20169_),
    .ZN(_20170_)
  );
  AND2_X1 _55932_ (
    .A1(_10690_),
    .A2(_20167_),
    .ZN(_20171_)
  );
  INV_X1 _55933_ (
    .A(_20171_),
    .ZN(_20172_)
  );
  AND2_X1 _55934_ (
    .A1(_20170_),
    .A2(_20172_),
    .ZN(_20173_)
  );
  AND2_X1 _55935_ (
    .A1(instr_sub),
    .A2(_20173_),
    .ZN(_20174_)
  );
  INV_X1 _55936_ (
    .A(_20174_),
    .ZN(_20175_)
  );
  AND2_X1 _55937_ (
    .A1(_20166_),
    .A2(_20175_),
    .ZN(_20176_)
  );
  INV_X1 _55938_ (
    .A(_20176_),
    .ZN(_20177_)
  );
  AND2_X1 _55939_ (
    .A1(is_lui_auipc_jal_jalr_addi_add_sub),
    .A2(_20177_),
    .ZN(_20178_)
  );
  INV_X1 _55940_ (
    .A(_20178_),
    .ZN(_20179_)
  );
  AND2_X1 _55941_ (
    .A1(_22528_),
    .A2(_10927_),
    .ZN(_20180_)
  );
  INV_X1 _55942_ (
    .A(_20180_),
    .ZN(_20181_)
  );
  AND2_X1 _55943_ (
    .A1(_10923_),
    .A2(_20097_),
    .ZN(_20182_)
  );
  INV_X1 _55944_ (
    .A(_20182_),
    .ZN(_20183_)
  );
  AND2_X1 _55945_ (
    .A1(_22532_),
    .A2(_10926_),
    .ZN(_20184_)
  );
  INV_X1 _55946_ (
    .A(_20184_),
    .ZN(_20185_)
  );
  AND2_X1 _55947_ (
    .A1(_20183_),
    .A2(_20185_),
    .ZN(_20186_)
  );
  AND2_X1 _55948_ (
    .A1(_20181_),
    .A2(_20186_),
    .ZN(_20187_)
  );
  AND2_X1 _55949_ (
    .A1(_20179_),
    .A2(_20187_),
    .ZN(_20188_)
  );
  INV_X1 _55950_ (
    .A(_20188_),
    .ZN(alu_out[3])
  );
  AND2_X1 _55951_ (
    .A1(_10664_),
    .A2(_10695_),
    .ZN(_20189_)
  );
  INV_X1 _55952_ (
    .A(_20189_),
    .ZN(_20190_)
  );
  AND2_X1 _55953_ (
    .A1(_10698_),
    .A2(_20092_),
    .ZN(_20191_)
  );
  AND2_X1 _55954_ (
    .A1(_20190_),
    .A2(_20191_),
    .ZN(_20192_)
  );
  INV_X1 _55955_ (
    .A(_20192_),
    .ZN(_20193_)
  );
  AND2_X1 _55956_ (
    .A1(_10924_),
    .A2(_20161_),
    .ZN(_20194_)
  );
  INV_X1 _55957_ (
    .A(_20194_),
    .ZN(_20195_)
  );
  AND2_X1 _55958_ (
    .A1(_11005_),
    .A2(_20195_),
    .ZN(_20196_)
  );
  INV_X1 _55959_ (
    .A(_20196_),
    .ZN(_20197_)
  );
  AND2_X1 _55960_ (
    .A1(_11006_),
    .A2(_20194_),
    .ZN(_20198_)
  );
  INV_X1 _55961_ (
    .A(_20198_),
    .ZN(_20199_)
  );
  AND2_X1 _55962_ (
    .A1(_20082_),
    .A2(_20199_),
    .ZN(_20200_)
  );
  AND2_X1 _55963_ (
    .A1(_20197_),
    .A2(_20200_),
    .ZN(_20201_)
  );
  INV_X1 _55964_ (
    .A(_20201_),
    .ZN(_20202_)
  );
  AND2_X1 _55965_ (
    .A1(_22528_),
    .A2(_11005_),
    .ZN(_20203_)
  );
  INV_X1 _55966_ (
    .A(_20203_),
    .ZN(_20204_)
  );
  AND2_X1 _55967_ (
    .A1(_11001_),
    .A2(_20097_),
    .ZN(_20205_)
  );
  INV_X1 _55968_ (
    .A(_20205_),
    .ZN(_20206_)
  );
  AND2_X1 _55969_ (
    .A1(_22532_),
    .A2(_11004_),
    .ZN(_20207_)
  );
  INV_X1 _55970_ (
    .A(_20207_),
    .ZN(_20208_)
  );
  AND2_X1 _55971_ (
    .A1(_20206_),
    .A2(_20208_),
    .ZN(_20209_)
  );
  AND2_X1 _55972_ (
    .A1(_20204_),
    .A2(_20209_),
    .ZN(_20210_)
  );
  AND2_X1 _55973_ (
    .A1(_20193_),
    .A2(_20210_),
    .ZN(_20211_)
  );
  AND2_X1 _55974_ (
    .A1(_20202_),
    .A2(_20211_),
    .ZN(_20212_)
  );
  INV_X1 _55975_ (
    .A(_20212_),
    .ZN(alu_out[4])
  );
  AND2_X1 _55976_ (
    .A1(_11002_),
    .A2(_20197_),
    .ZN(_20213_)
  );
  INV_X1 _55977_ (
    .A(_20213_),
    .ZN(_20214_)
  );
  AND2_X1 _55978_ (
    .A1(_10994_),
    .A2(_20213_),
    .ZN(_20215_)
  );
  INV_X1 _55979_ (
    .A(_20215_),
    .ZN(_20216_)
  );
  AND2_X1 _55980_ (
    .A1(_10993_),
    .A2(_20214_),
    .ZN(_20217_)
  );
  INV_X1 _55981_ (
    .A(_20217_),
    .ZN(_20218_)
  );
  AND2_X1 _55982_ (
    .A1(_20216_),
    .A2(_20218_),
    .ZN(_20219_)
  );
  AND2_X1 _55983_ (
    .A1(_20082_),
    .A2(_20219_),
    .ZN(_20220_)
  );
  INV_X1 _55984_ (
    .A(_20220_),
    .ZN(_20221_)
  );
  AND2_X1 _55985_ (
    .A1(_10656_),
    .A2(_10658_),
    .ZN(_20222_)
  );
  INV_X1 _55986_ (
    .A(_20222_),
    .ZN(_20223_)
  );
  AND2_X1 _55987_ (
    .A1(_10700_),
    .A2(_20222_),
    .ZN(_20224_)
  );
  INV_X1 _55988_ (
    .A(_20224_),
    .ZN(_20225_)
  );
  AND2_X1 _55989_ (
    .A1(_10699_),
    .A2(_20223_),
    .ZN(_20226_)
  );
  INV_X1 _55990_ (
    .A(_20226_),
    .ZN(_20227_)
  );
  AND2_X1 _55991_ (
    .A1(_20092_),
    .A2(_20227_),
    .ZN(_20228_)
  );
  AND2_X1 _55992_ (
    .A1(_20225_),
    .A2(_20228_),
    .ZN(_20229_)
  );
  INV_X1 _55993_ (
    .A(_20229_),
    .ZN(_20230_)
  );
  AND2_X1 _55994_ (
    .A1(_22528_),
    .A2(_10993_),
    .ZN(_20231_)
  );
  INV_X1 _55995_ (
    .A(_20231_),
    .ZN(_20232_)
  );
  AND2_X1 _55996_ (
    .A1(_10989_),
    .A2(_20097_),
    .ZN(_20233_)
  );
  INV_X1 _55997_ (
    .A(_20233_),
    .ZN(_20234_)
  );
  AND2_X1 _55998_ (
    .A1(_22532_),
    .A2(_10992_),
    .ZN(_20235_)
  );
  INV_X1 _55999_ (
    .A(_20235_),
    .ZN(_20236_)
  );
  AND2_X1 _56000_ (
    .A1(_20234_),
    .A2(_20236_),
    .ZN(_20237_)
  );
  AND2_X1 _56001_ (
    .A1(_20232_),
    .A2(_20237_),
    .ZN(_20238_)
  );
  AND2_X1 _56002_ (
    .A1(_20230_),
    .A2(_20238_),
    .ZN(_20239_)
  );
  AND2_X1 _56003_ (
    .A1(_20221_),
    .A2(_20239_),
    .ZN(_20240_)
  );
  INV_X1 _56004_ (
    .A(_20240_),
    .ZN(alu_out[5])
  );
  AND2_X1 _56005_ (
    .A1(_10990_),
    .A2(_20218_),
    .ZN(_20241_)
  );
  INV_X1 _56006_ (
    .A(_20241_),
    .ZN(_20242_)
  );
  AND2_X1 _56007_ (
    .A1(_10934_),
    .A2(_20241_),
    .ZN(_20243_)
  );
  INV_X1 _56008_ (
    .A(_20243_),
    .ZN(_20244_)
  );
  AND2_X1 _56009_ (
    .A1(_10933_),
    .A2(_20242_),
    .ZN(_20245_)
  );
  INV_X1 _56010_ (
    .A(_20245_),
    .ZN(_20246_)
  );
  AND2_X1 _56011_ (
    .A1(_20244_),
    .A2(_20246_),
    .ZN(_20247_)
  );
  AND2_X1 _56012_ (
    .A1(_20082_),
    .A2(_20247_),
    .ZN(_20248_)
  );
  INV_X1 _56013_ (
    .A(_20248_),
    .ZN(_20249_)
  );
  AND2_X1 _56014_ (
    .A1(_10654_),
    .A2(_10705_),
    .ZN(_20250_)
  );
  INV_X1 _56015_ (
    .A(_20250_),
    .ZN(_20251_)
  );
  AND2_X1 _56016_ (
    .A1(_10708_),
    .A2(_20092_),
    .ZN(_20252_)
  );
  AND2_X1 _56017_ (
    .A1(_20251_),
    .A2(_20252_),
    .ZN(_20253_)
  );
  INV_X1 _56018_ (
    .A(_20253_),
    .ZN(_20254_)
  );
  AND2_X1 _56019_ (
    .A1(_22528_),
    .A2(_10933_),
    .ZN(_20255_)
  );
  INV_X1 _56020_ (
    .A(_20255_),
    .ZN(_20256_)
  );
  AND2_X1 _56021_ (
    .A1(_10929_),
    .A2(_20097_),
    .ZN(_20257_)
  );
  INV_X1 _56022_ (
    .A(_20257_),
    .ZN(_20258_)
  );
  AND2_X1 _56023_ (
    .A1(_22532_),
    .A2(_10932_),
    .ZN(_20259_)
  );
  INV_X1 _56024_ (
    .A(_20259_),
    .ZN(_20260_)
  );
  AND2_X1 _56025_ (
    .A1(_20258_),
    .A2(_20260_),
    .ZN(_20261_)
  );
  AND2_X1 _56026_ (
    .A1(_20256_),
    .A2(_20261_),
    .ZN(_20262_)
  );
  AND2_X1 _56027_ (
    .A1(_20254_),
    .A2(_20262_),
    .ZN(_20263_)
  );
  AND2_X1 _56028_ (
    .A1(_20249_),
    .A2(_20263_),
    .ZN(_20264_)
  );
  INV_X1 _56029_ (
    .A(_20264_),
    .ZN(alu_out[6])
  );
  AND2_X1 _56030_ (
    .A1(_10930_),
    .A2(_20246_),
    .ZN(_20265_)
  );
  INV_X1 _56031_ (
    .A(_20265_),
    .ZN(_20266_)
  );
  AND2_X1 _56032_ (
    .A1(_10963_),
    .A2(_20265_),
    .ZN(_20267_)
  );
  INV_X1 _56033_ (
    .A(_20267_),
    .ZN(_20268_)
  );
  AND2_X1 _56034_ (
    .A1(_10964_),
    .A2(_20266_),
    .ZN(_20269_)
  );
  INV_X1 _56035_ (
    .A(_20269_),
    .ZN(_20270_)
  );
  AND2_X1 _56036_ (
    .A1(_20268_),
    .A2(_20270_),
    .ZN(_20271_)
  );
  AND2_X1 _56037_ (
    .A1(_21049_),
    .A2(_20271_),
    .ZN(_20272_)
  );
  INV_X1 _56038_ (
    .A(_20272_),
    .ZN(_20273_)
  );
  AND2_X1 _56039_ (
    .A1(_10646_),
    .A2(_10648_),
    .ZN(_20274_)
  );
  INV_X1 _56040_ (
    .A(_20274_),
    .ZN(_20275_)
  );
  AND2_X1 _56041_ (
    .A1(_10709_),
    .A2(_20274_),
    .ZN(_20276_)
  );
  INV_X1 _56042_ (
    .A(_20276_),
    .ZN(_20277_)
  );
  AND2_X1 _56043_ (
    .A1(_10710_),
    .A2(_20275_),
    .ZN(_20278_)
  );
  INV_X1 _56044_ (
    .A(_20278_),
    .ZN(_20279_)
  );
  AND2_X1 _56045_ (
    .A1(instr_sub),
    .A2(_20277_),
    .ZN(_20280_)
  );
  AND2_X1 _56046_ (
    .A1(_20279_),
    .A2(_20280_),
    .ZN(_20281_)
  );
  INV_X1 _56047_ (
    .A(_20281_),
    .ZN(_20282_)
  );
  AND2_X1 _56048_ (
    .A1(is_lui_auipc_jal_jalr_addi_add_sub),
    .A2(_20282_),
    .ZN(_20283_)
  );
  AND2_X1 _56049_ (
    .A1(_20273_),
    .A2(_20283_),
    .ZN(_20284_)
  );
  INV_X1 _56050_ (
    .A(_20284_),
    .ZN(_20285_)
  );
  AND2_X1 _56051_ (
    .A1(_22528_),
    .A2(_10963_),
    .ZN(_20286_)
  );
  INV_X1 _56052_ (
    .A(_20286_),
    .ZN(_20287_)
  );
  AND2_X1 _56053_ (
    .A1(_10959_),
    .A2(_20097_),
    .ZN(_20288_)
  );
  INV_X1 _56054_ (
    .A(_20288_),
    .ZN(_20289_)
  );
  AND2_X1 _56055_ (
    .A1(_22532_),
    .A2(_10962_),
    .ZN(_20290_)
  );
  INV_X1 _56056_ (
    .A(_20290_),
    .ZN(_20291_)
  );
  AND2_X1 _56057_ (
    .A1(_20289_),
    .A2(_20291_),
    .ZN(_20292_)
  );
  AND2_X1 _56058_ (
    .A1(_20287_),
    .A2(_20292_),
    .ZN(_20293_)
  );
  AND2_X1 _56059_ (
    .A1(_20285_),
    .A2(_20293_),
    .ZN(_20294_)
  );
  INV_X1 _56060_ (
    .A(_20294_),
    .ZN(alu_out[7])
  );
  AND2_X1 _56061_ (
    .A1(_10962_),
    .A2(_20266_),
    .ZN(_20295_)
  );
  INV_X1 _56062_ (
    .A(_20295_),
    .ZN(_20296_)
  );
  AND2_X1 _56063_ (
    .A1(_10960_),
    .A2(_20265_),
    .ZN(_20297_)
  );
  INV_X1 _56064_ (
    .A(_20297_),
    .ZN(_20298_)
  );
  AND2_X1 _56065_ (
    .A1(_10960_),
    .A2(_20296_),
    .ZN(_20299_)
  );
  AND2_X1 _56066_ (
    .A1(_10962_),
    .A2(_20298_),
    .ZN(_20300_)
  );
  AND2_X1 _56067_ (
    .A1(_10873_),
    .A2(_20300_),
    .ZN(_20301_)
  );
  INV_X1 _56068_ (
    .A(_20301_),
    .ZN(_20302_)
  );
  AND2_X1 _56069_ (
    .A1(_10874_),
    .A2(_20299_),
    .ZN(_20303_)
  );
  INV_X1 _56070_ (
    .A(_20303_),
    .ZN(_20304_)
  );
  AND2_X1 _56071_ (
    .A1(_20302_),
    .A2(_20304_),
    .ZN(_20305_)
  );
  AND2_X1 _56072_ (
    .A1(_20082_),
    .A2(_20305_),
    .ZN(_20306_)
  );
  INV_X1 _56073_ (
    .A(_20306_),
    .ZN(_20307_)
  );
  AND2_X1 _56074_ (
    .A1(_10644_),
    .A2(_10715_),
    .ZN(_20308_)
  );
  INV_X1 _56075_ (
    .A(_20308_),
    .ZN(_20309_)
  );
  AND2_X1 _56076_ (
    .A1(_10718_),
    .A2(_20092_),
    .ZN(_20310_)
  );
  AND2_X1 _56077_ (
    .A1(_20309_),
    .A2(_20310_),
    .ZN(_20311_)
  );
  INV_X1 _56078_ (
    .A(_20311_),
    .ZN(_20312_)
  );
  AND2_X1 _56079_ (
    .A1(_22528_),
    .A2(_10873_),
    .ZN(_20313_)
  );
  INV_X1 _56080_ (
    .A(_20313_),
    .ZN(_20314_)
  );
  AND2_X1 _56081_ (
    .A1(_10869_),
    .A2(_20097_),
    .ZN(_20315_)
  );
  INV_X1 _56082_ (
    .A(_20315_),
    .ZN(_20316_)
  );
  AND2_X1 _56083_ (
    .A1(_22532_),
    .A2(_10872_),
    .ZN(_20317_)
  );
  INV_X1 _56084_ (
    .A(_20317_),
    .ZN(_20318_)
  );
  AND2_X1 _56085_ (
    .A1(_20316_),
    .A2(_20318_),
    .ZN(_20319_)
  );
  AND2_X1 _56086_ (
    .A1(_20314_),
    .A2(_20319_),
    .ZN(_20320_)
  );
  AND2_X1 _56087_ (
    .A1(_20312_),
    .A2(_20320_),
    .ZN(_20321_)
  );
  AND2_X1 _56088_ (
    .A1(_20307_),
    .A2(_20321_),
    .ZN(_20322_)
  );
  INV_X1 _56089_ (
    .A(_20322_),
    .ZN(alu_out[8])
  );
  AND2_X1 _56090_ (
    .A1(_10870_),
    .A2(_20302_),
    .ZN(_20323_)
  );
  INV_X1 _56091_ (
    .A(_20323_),
    .ZN(_20324_)
  );
  AND2_X1 _56092_ (
    .A1(_10861_),
    .A2(_20324_),
    .ZN(_20325_)
  );
  INV_X1 _56093_ (
    .A(_20325_),
    .ZN(_20326_)
  );
  AND2_X1 _56094_ (
    .A1(_10862_),
    .A2(_20323_),
    .ZN(_20327_)
  );
  INV_X1 _56095_ (
    .A(_20327_),
    .ZN(_20328_)
  );
  AND2_X1 _56096_ (
    .A1(_20326_),
    .A2(_20328_),
    .ZN(_20329_)
  );
  AND2_X1 _56097_ (
    .A1(_10636_),
    .A2(_10638_),
    .ZN(_20330_)
  );
  INV_X1 _56098_ (
    .A(_20330_),
    .ZN(_20331_)
  );
  AND2_X1 _56099_ (
    .A1(_10719_),
    .A2(_20331_),
    .ZN(_20332_)
  );
  INV_X1 _56100_ (
    .A(_20332_),
    .ZN(_20333_)
  );
  AND2_X1 _56101_ (
    .A1(_10720_),
    .A2(_20330_),
    .ZN(_20334_)
  );
  INV_X1 _56102_ (
    .A(_20334_),
    .ZN(_20335_)
  );
  AND2_X1 _56103_ (
    .A1(_20333_),
    .A2(_20335_),
    .ZN(_20336_)
  );
  AND2_X1 _56104_ (
    .A1(instr_sub),
    .A2(_20336_),
    .ZN(_20337_)
  );
  INV_X1 _56105_ (
    .A(_20337_),
    .ZN(_20338_)
  );
  AND2_X1 _56106_ (
    .A1(_21049_),
    .A2(_20329_),
    .ZN(_20339_)
  );
  INV_X1 _56107_ (
    .A(_20339_),
    .ZN(_20340_)
  );
  AND2_X1 _56108_ (
    .A1(_20338_),
    .A2(_20340_),
    .ZN(_20341_)
  );
  INV_X1 _56109_ (
    .A(_20341_),
    .ZN(_20342_)
  );
  AND2_X1 _56110_ (
    .A1(is_lui_auipc_jal_jalr_addi_add_sub),
    .A2(_20342_),
    .ZN(_20343_)
  );
  INV_X1 _56111_ (
    .A(_20343_),
    .ZN(_20344_)
  );
  AND2_X1 _56112_ (
    .A1(_22528_),
    .A2(_10861_),
    .ZN(_20345_)
  );
  INV_X1 _56113_ (
    .A(_20345_),
    .ZN(_20346_)
  );
  AND2_X1 _56114_ (
    .A1(_10857_),
    .A2(_20097_),
    .ZN(_20347_)
  );
  INV_X1 _56115_ (
    .A(_20347_),
    .ZN(_20348_)
  );
  AND2_X1 _56116_ (
    .A1(_22532_),
    .A2(_10860_),
    .ZN(_20349_)
  );
  INV_X1 _56117_ (
    .A(_20349_),
    .ZN(_20350_)
  );
  AND2_X1 _56118_ (
    .A1(_20348_),
    .A2(_20350_),
    .ZN(_20351_)
  );
  AND2_X1 _56119_ (
    .A1(_20346_),
    .A2(_20351_),
    .ZN(_20352_)
  );
  AND2_X1 _56120_ (
    .A1(_20344_),
    .A2(_20352_),
    .ZN(_20353_)
  );
  INV_X1 _56121_ (
    .A(_20353_),
    .ZN(alu_out[9])
  );
  AND2_X1 _56122_ (
    .A1(_10634_),
    .A2(_10725_),
    .ZN(_20354_)
  );
  INV_X1 _56123_ (
    .A(_20354_),
    .ZN(_20355_)
  );
  AND2_X1 _56124_ (
    .A1(instr_sub),
    .A2(_10728_),
    .ZN(_20356_)
  );
  AND2_X1 _56125_ (
    .A1(_20355_),
    .A2(_20356_),
    .ZN(_20357_)
  );
  INV_X1 _56126_ (
    .A(_20357_),
    .ZN(_20358_)
  );
  AND2_X1 _56127_ (
    .A1(_10860_),
    .A2(_20324_),
    .ZN(_20359_)
  );
  INV_X1 _56128_ (
    .A(_20359_),
    .ZN(_20360_)
  );
  AND2_X1 _56129_ (
    .A1(_10858_),
    .A2(_20323_),
    .ZN(_20361_)
  );
  INV_X1 _56130_ (
    .A(_20361_),
    .ZN(_20362_)
  );
  AND2_X1 _56131_ (
    .A1(_10858_),
    .A2(_20360_),
    .ZN(_20363_)
  );
  AND2_X1 _56132_ (
    .A1(_10860_),
    .A2(_20362_),
    .ZN(_20364_)
  );
  AND2_X1 _56133_ (
    .A1(_10897_),
    .A2(_20364_),
    .ZN(_20365_)
  );
  INV_X1 _56134_ (
    .A(_20365_),
    .ZN(_20366_)
  );
  AND2_X1 _56135_ (
    .A1(_10898_),
    .A2(_20363_),
    .ZN(_20367_)
  );
  INV_X1 _56136_ (
    .A(_20367_),
    .ZN(_20368_)
  );
  AND2_X1 _56137_ (
    .A1(_21049_),
    .A2(_20366_),
    .ZN(_20369_)
  );
  AND2_X1 _56138_ (
    .A1(_20368_),
    .A2(_20369_),
    .ZN(_20370_)
  );
  INV_X1 _56139_ (
    .A(_20370_),
    .ZN(_20371_)
  );
  AND2_X1 _56140_ (
    .A1(_20358_),
    .A2(_20371_),
    .ZN(_20372_)
  );
  INV_X1 _56141_ (
    .A(_20372_),
    .ZN(_20373_)
  );
  AND2_X1 _56142_ (
    .A1(is_lui_auipc_jal_jalr_addi_add_sub),
    .A2(_20373_),
    .ZN(_20374_)
  );
  INV_X1 _56143_ (
    .A(_20374_),
    .ZN(_20375_)
  );
  AND2_X1 _56144_ (
    .A1(_22528_),
    .A2(_10897_),
    .ZN(_20376_)
  );
  INV_X1 _56145_ (
    .A(_20376_),
    .ZN(_20377_)
  );
  AND2_X1 _56146_ (
    .A1(_22532_),
    .A2(_10896_),
    .ZN(_20378_)
  );
  INV_X1 _56147_ (
    .A(_20378_),
    .ZN(_20379_)
  );
  AND2_X1 _56148_ (
    .A1(_10893_),
    .A2(_20097_),
    .ZN(_20380_)
  );
  INV_X1 _56149_ (
    .A(_20380_),
    .ZN(_20381_)
  );
  AND2_X1 _56150_ (
    .A1(_20379_),
    .A2(_20381_),
    .ZN(_20382_)
  );
  AND2_X1 _56151_ (
    .A1(_20377_),
    .A2(_20382_),
    .ZN(_20383_)
  );
  AND2_X1 _56152_ (
    .A1(_20375_),
    .A2(_20383_),
    .ZN(_20384_)
  );
  INV_X1 _56153_ (
    .A(_20384_),
    .ZN(alu_out[10])
  );
  AND2_X1 _56154_ (
    .A1(_10894_),
    .A2(_20366_),
    .ZN(_20385_)
  );
  INV_X1 _56155_ (
    .A(_20385_),
    .ZN(_20386_)
  );
  AND2_X1 _56156_ (
    .A1(_10909_),
    .A2(_20386_),
    .ZN(_20387_)
  );
  INV_X1 _56157_ (
    .A(_20387_),
    .ZN(_20388_)
  );
  AND2_X1 _56158_ (
    .A1(_10910_),
    .A2(_20385_),
    .ZN(_20389_)
  );
  INV_X1 _56159_ (
    .A(_20389_),
    .ZN(_20390_)
  );
  AND2_X1 _56160_ (
    .A1(_20388_),
    .A2(_20390_),
    .ZN(_20391_)
  );
  AND2_X1 _56161_ (
    .A1(_10626_),
    .A2(_10628_),
    .ZN(_20392_)
  );
  INV_X1 _56162_ (
    .A(_20392_),
    .ZN(_20393_)
  );
  AND2_X1 _56163_ (
    .A1(_10729_),
    .A2(_20393_),
    .ZN(_20394_)
  );
  INV_X1 _56164_ (
    .A(_20394_),
    .ZN(_20395_)
  );
  AND2_X1 _56165_ (
    .A1(_10730_),
    .A2(_20392_),
    .ZN(_20396_)
  );
  INV_X1 _56166_ (
    .A(_20396_),
    .ZN(_20397_)
  );
  AND2_X1 _56167_ (
    .A1(_20395_),
    .A2(_20397_),
    .ZN(_20398_)
  );
  AND2_X1 _56168_ (
    .A1(instr_sub),
    .A2(_20398_),
    .ZN(_20399_)
  );
  INV_X1 _56169_ (
    .A(_20399_),
    .ZN(_20400_)
  );
  AND2_X1 _56170_ (
    .A1(_21049_),
    .A2(_20391_),
    .ZN(_20401_)
  );
  INV_X1 _56171_ (
    .A(_20401_),
    .ZN(_20402_)
  );
  AND2_X1 _56172_ (
    .A1(_20400_),
    .A2(_20402_),
    .ZN(_20403_)
  );
  INV_X1 _56173_ (
    .A(_20403_),
    .ZN(_20404_)
  );
  AND2_X1 _56174_ (
    .A1(is_lui_auipc_jal_jalr_addi_add_sub),
    .A2(_20404_),
    .ZN(_20405_)
  );
  INV_X1 _56175_ (
    .A(_20405_),
    .ZN(_20406_)
  );
  AND2_X1 _56176_ (
    .A1(_22528_),
    .A2(_10909_),
    .ZN(_20407_)
  );
  INV_X1 _56177_ (
    .A(_20407_),
    .ZN(_20408_)
  );
  AND2_X1 _56178_ (
    .A1(_22532_),
    .A2(_10908_),
    .ZN(_20409_)
  );
  INV_X1 _56179_ (
    .A(_20409_),
    .ZN(_20410_)
  );
  AND2_X1 _56180_ (
    .A1(_10905_),
    .A2(_20097_),
    .ZN(_20411_)
  );
  INV_X1 _56181_ (
    .A(_20411_),
    .ZN(_20412_)
  );
  AND2_X1 _56182_ (
    .A1(_20410_),
    .A2(_20412_),
    .ZN(_20413_)
  );
  AND2_X1 _56183_ (
    .A1(_20408_),
    .A2(_20413_),
    .ZN(_20414_)
  );
  AND2_X1 _56184_ (
    .A1(_20406_),
    .A2(_20414_),
    .ZN(_20415_)
  );
  INV_X1 _56185_ (
    .A(_20415_),
    .ZN(alu_out[11])
  );
  AND2_X1 _56186_ (
    .A1(_10908_),
    .A2(_20386_),
    .ZN(_20416_)
  );
  INV_X1 _56187_ (
    .A(_20416_),
    .ZN(_20417_)
  );
  AND2_X1 _56188_ (
    .A1(_10906_),
    .A2(_20385_),
    .ZN(_20418_)
  );
  INV_X1 _56189_ (
    .A(_20418_),
    .ZN(_20419_)
  );
  AND2_X1 _56190_ (
    .A1(_10906_),
    .A2(_20417_),
    .ZN(_20420_)
  );
  AND2_X1 _56191_ (
    .A1(_10908_),
    .A2(_20419_),
    .ZN(_20421_)
  );
  AND2_X1 _56192_ (
    .A1(_11012_),
    .A2(_20420_),
    .ZN(_20422_)
  );
  INV_X1 _56193_ (
    .A(_20422_),
    .ZN(_20423_)
  );
  AND2_X1 _56194_ (
    .A1(_11011_),
    .A2(_20421_),
    .ZN(_20424_)
  );
  INV_X1 _56195_ (
    .A(_20424_),
    .ZN(_20425_)
  );
  AND2_X1 _56196_ (
    .A1(_10624_),
    .A2(_10735_),
    .ZN(_20426_)
  );
  INV_X1 _56197_ (
    .A(_20426_),
    .ZN(_20427_)
  );
  AND2_X1 _56198_ (
    .A1(_21049_),
    .A2(_20425_),
    .ZN(_20428_)
  );
  AND2_X1 _56199_ (
    .A1(_20423_),
    .A2(_20428_),
    .ZN(_20429_)
  );
  INV_X1 _56200_ (
    .A(_20429_),
    .ZN(_20430_)
  );
  AND2_X1 _56201_ (
    .A1(instr_sub),
    .A2(_10738_),
    .ZN(_20431_)
  );
  AND2_X1 _56202_ (
    .A1(_20427_),
    .A2(_20431_),
    .ZN(_20432_)
  );
  INV_X1 _56203_ (
    .A(_20432_),
    .ZN(_20433_)
  );
  AND2_X1 _56204_ (
    .A1(_20430_),
    .A2(_20433_),
    .ZN(_20434_)
  );
  INV_X1 _56205_ (
    .A(_20434_),
    .ZN(_20435_)
  );
  AND2_X1 _56206_ (
    .A1(is_lui_auipc_jal_jalr_addi_add_sub),
    .A2(_20435_),
    .ZN(_20436_)
  );
  INV_X1 _56207_ (
    .A(_20436_),
    .ZN(_20437_)
  );
  AND2_X1 _56208_ (
    .A1(_22528_),
    .A2(_11011_),
    .ZN(_20438_)
  );
  INV_X1 _56209_ (
    .A(_20438_),
    .ZN(_20439_)
  );
  AND2_X1 _56210_ (
    .A1(_11007_),
    .A2(_20097_),
    .ZN(_20440_)
  );
  INV_X1 _56211_ (
    .A(_20440_),
    .ZN(_20441_)
  );
  AND2_X1 _56212_ (
    .A1(_22532_),
    .A2(_11010_),
    .ZN(_20442_)
  );
  INV_X1 _56213_ (
    .A(_20442_),
    .ZN(_20443_)
  );
  AND2_X1 _56214_ (
    .A1(_20441_),
    .A2(_20443_),
    .ZN(_20444_)
  );
  AND2_X1 _56215_ (
    .A1(_20439_),
    .A2(_20444_),
    .ZN(_20445_)
  );
  AND2_X1 _56216_ (
    .A1(_20437_),
    .A2(_20445_),
    .ZN(_20446_)
  );
  INV_X1 _56217_ (
    .A(_20446_),
    .ZN(alu_out[12])
  );
  AND2_X1 _56218_ (
    .A1(_11008_),
    .A2(_20425_),
    .ZN(_20447_)
  );
  INV_X1 _56219_ (
    .A(_20447_),
    .ZN(_20448_)
  );
  AND2_X1 _56220_ (
    .A1(_10969_),
    .A2(_20448_),
    .ZN(_20449_)
  );
  INV_X1 _56221_ (
    .A(_20449_),
    .ZN(_20450_)
  );
  AND2_X1 _56222_ (
    .A1(_10970_),
    .A2(_20447_),
    .ZN(_20451_)
  );
  INV_X1 _56223_ (
    .A(_20451_),
    .ZN(_20452_)
  );
  AND2_X1 _56224_ (
    .A1(_21049_),
    .A2(_20452_),
    .ZN(_20453_)
  );
  AND2_X1 _56225_ (
    .A1(_20450_),
    .A2(_20453_),
    .ZN(_20454_)
  );
  INV_X1 _56226_ (
    .A(_20454_),
    .ZN(_20455_)
  );
  AND2_X1 _56227_ (
    .A1(_10616_),
    .A2(_10618_),
    .ZN(_20456_)
  );
  INV_X1 _56228_ (
    .A(_20456_),
    .ZN(_20457_)
  );
  AND2_X1 _56229_ (
    .A1(_10739_),
    .A2(_20457_),
    .ZN(_20458_)
  );
  INV_X1 _56230_ (
    .A(_20458_),
    .ZN(_20459_)
  );
  AND2_X1 _56231_ (
    .A1(_10740_),
    .A2(_20456_),
    .ZN(_20460_)
  );
  INV_X1 _56232_ (
    .A(_20460_),
    .ZN(_20461_)
  );
  AND2_X1 _56233_ (
    .A1(instr_sub),
    .A2(_20461_),
    .ZN(_20462_)
  );
  AND2_X1 _56234_ (
    .A1(_20459_),
    .A2(_20462_),
    .ZN(_20463_)
  );
  INV_X1 _56235_ (
    .A(_20463_),
    .ZN(_20464_)
  );
  AND2_X1 _56236_ (
    .A1(_20455_),
    .A2(_20464_),
    .ZN(_20465_)
  );
  INV_X1 _56237_ (
    .A(_20465_),
    .ZN(_20466_)
  );
  AND2_X1 _56238_ (
    .A1(is_lui_auipc_jal_jalr_addi_add_sub),
    .A2(_20466_),
    .ZN(_20467_)
  );
  INV_X1 _56239_ (
    .A(_20467_),
    .ZN(_20468_)
  );
  AND2_X1 _56240_ (
    .A1(_22528_),
    .A2(_10969_),
    .ZN(_20469_)
  );
  INV_X1 _56241_ (
    .A(_20469_),
    .ZN(_20470_)
  );
  AND2_X1 _56242_ (
    .A1(_10965_),
    .A2(_20097_),
    .ZN(_20471_)
  );
  INV_X1 _56243_ (
    .A(_20471_),
    .ZN(_20472_)
  );
  AND2_X1 _56244_ (
    .A1(_22532_),
    .A2(_10968_),
    .ZN(_20473_)
  );
  INV_X1 _56245_ (
    .A(_20473_),
    .ZN(_20474_)
  );
  AND2_X1 _56246_ (
    .A1(_20472_),
    .A2(_20474_),
    .ZN(_20475_)
  );
  AND2_X1 _56247_ (
    .A1(_20470_),
    .A2(_20475_),
    .ZN(_20476_)
  );
  AND2_X1 _56248_ (
    .A1(_20468_),
    .A2(_20476_),
    .ZN(_20477_)
  );
  INV_X1 _56249_ (
    .A(_20477_),
    .ZN(alu_out[13])
  );
  AND2_X1 _56250_ (
    .A1(_10614_),
    .A2(_10745_),
    .ZN(_20478_)
  );
  INV_X1 _56251_ (
    .A(_20478_),
    .ZN(_20479_)
  );
  AND2_X1 _56252_ (
    .A1(instr_sub),
    .A2(_10748_),
    .ZN(_20480_)
  );
  AND2_X1 _56253_ (
    .A1(_20479_),
    .A2(_20480_),
    .ZN(_20481_)
  );
  INV_X1 _56254_ (
    .A(_20481_),
    .ZN(_20482_)
  );
  AND2_X1 _56255_ (
    .A1(_10966_),
    .A2(_11008_),
    .ZN(_20483_)
  );
  INV_X1 _56256_ (
    .A(_20483_),
    .ZN(_20484_)
  );
  AND2_X1 _56257_ (
    .A1(_20425_),
    .A2(_20483_),
    .ZN(_20485_)
  );
  INV_X1 _56258_ (
    .A(_20485_),
    .ZN(_20486_)
  );
  AND2_X1 _56259_ (
    .A1(_10968_),
    .A2(_20486_),
    .ZN(_20487_)
  );
  INV_X1 _56260_ (
    .A(_20487_),
    .ZN(_20488_)
  );
  AND2_X1 _56261_ (
    .A1(_10891_),
    .A2(_20487_),
    .ZN(_20489_)
  );
  INV_X1 _56262_ (
    .A(_20489_),
    .ZN(_20490_)
  );
  AND2_X1 _56263_ (
    .A1(_10892_),
    .A2(_20488_),
    .ZN(_20491_)
  );
  INV_X1 _56264_ (
    .A(_20491_),
    .ZN(_20492_)
  );
  AND2_X1 _56265_ (
    .A1(_21049_),
    .A2(_20490_),
    .ZN(_20493_)
  );
  AND2_X1 _56266_ (
    .A1(_20492_),
    .A2(_20493_),
    .ZN(_20494_)
  );
  INV_X1 _56267_ (
    .A(_20494_),
    .ZN(_20495_)
  );
  AND2_X1 _56268_ (
    .A1(_20482_),
    .A2(_20495_),
    .ZN(_20496_)
  );
  INV_X1 _56269_ (
    .A(_20496_),
    .ZN(_20497_)
  );
  AND2_X1 _56270_ (
    .A1(is_lui_auipc_jal_jalr_addi_add_sub),
    .A2(_20497_),
    .ZN(_20498_)
  );
  INV_X1 _56271_ (
    .A(_20498_),
    .ZN(_20499_)
  );
  AND2_X1 _56272_ (
    .A1(_22528_),
    .A2(_10891_),
    .ZN(_20500_)
  );
  INV_X1 _56273_ (
    .A(_20500_),
    .ZN(_20501_)
  );
  AND2_X1 _56274_ (
    .A1(_22532_),
    .A2(_10890_),
    .ZN(_20502_)
  );
  INV_X1 _56275_ (
    .A(_20502_),
    .ZN(_20503_)
  );
  AND2_X1 _56276_ (
    .A1(_10887_),
    .A2(_20097_),
    .ZN(_20504_)
  );
  INV_X1 _56277_ (
    .A(_20504_),
    .ZN(_20505_)
  );
  AND2_X1 _56278_ (
    .A1(_20503_),
    .A2(_20505_),
    .ZN(_20506_)
  );
  AND2_X1 _56279_ (
    .A1(_20501_),
    .A2(_20506_),
    .ZN(_20507_)
  );
  AND2_X1 _56280_ (
    .A1(_20499_),
    .A2(_20507_),
    .ZN(_20508_)
  );
  INV_X1 _56281_ (
    .A(_20508_),
    .ZN(alu_out[14])
  );
  AND2_X1 _56282_ (
    .A1(_10606_),
    .A2(_10608_),
    .ZN(_20509_)
  );
  INV_X1 _56283_ (
    .A(_20509_),
    .ZN(_20510_)
  );
  AND2_X1 _56284_ (
    .A1(_10749_),
    .A2(_20509_),
    .ZN(_20511_)
  );
  INV_X1 _56285_ (
    .A(_20511_),
    .ZN(_20512_)
  );
  AND2_X1 _56286_ (
    .A1(_10750_),
    .A2(_20510_),
    .ZN(_20513_)
  );
  INV_X1 _56287_ (
    .A(_20513_),
    .ZN(_20514_)
  );
  AND2_X1 _56288_ (
    .A1(instr_sub),
    .A2(_20512_),
    .ZN(_20515_)
  );
  AND2_X1 _56289_ (
    .A1(_20514_),
    .A2(_20515_),
    .ZN(_20516_)
  );
  INV_X1 _56290_ (
    .A(_20516_),
    .ZN(_20517_)
  );
  AND2_X1 _56291_ (
    .A1(_10888_),
    .A2(_20490_),
    .ZN(_20518_)
  );
  INV_X1 _56292_ (
    .A(_20518_),
    .ZN(_20519_)
  );
  AND2_X1 _56293_ (
    .A1(_10867_),
    .A2(_20519_),
    .ZN(_20520_)
  );
  INV_X1 _56294_ (
    .A(_20520_),
    .ZN(_20521_)
  );
  AND2_X1 _56295_ (
    .A1(_10868_),
    .A2(_20518_),
    .ZN(_20522_)
  );
  INV_X1 _56296_ (
    .A(_20522_),
    .ZN(_20523_)
  );
  AND2_X1 _56297_ (
    .A1(is_lui_auipc_jal_jalr_addi_add_sub),
    .A2(_20523_),
    .ZN(_20524_)
  );
  AND2_X1 _56298_ (
    .A1(_20521_),
    .A2(_20524_),
    .ZN(_20525_)
  );
  INV_X1 _56299_ (
    .A(_20525_),
    .ZN(_20526_)
  );
  AND2_X1 _56300_ (
    .A1(_20093_),
    .A2(_20526_),
    .ZN(_20527_)
  );
  INV_X1 _56301_ (
    .A(_20527_),
    .ZN(_20528_)
  );
  AND2_X1 _56302_ (
    .A1(_20517_),
    .A2(_20528_),
    .ZN(_20529_)
  );
  INV_X1 _56303_ (
    .A(_20529_),
    .ZN(_20530_)
  );
  AND2_X1 _56304_ (
    .A1(_22528_),
    .A2(_10867_),
    .ZN(_20531_)
  );
  INV_X1 _56305_ (
    .A(_20531_),
    .ZN(_20532_)
  );
  AND2_X1 _56306_ (
    .A1(_22532_),
    .A2(_10866_),
    .ZN(_20533_)
  );
  INV_X1 _56307_ (
    .A(_20533_),
    .ZN(_20534_)
  );
  AND2_X1 _56308_ (
    .A1(_10863_),
    .A2(_20097_),
    .ZN(_20535_)
  );
  INV_X1 _56309_ (
    .A(_20535_),
    .ZN(_20536_)
  );
  AND2_X1 _56310_ (
    .A1(_20534_),
    .A2(_20536_),
    .ZN(_20537_)
  );
  AND2_X1 _56311_ (
    .A1(_20532_),
    .A2(_20537_),
    .ZN(_20538_)
  );
  AND2_X1 _56312_ (
    .A1(_20530_),
    .A2(_20538_),
    .ZN(_20539_)
  );
  INV_X1 _56313_ (
    .A(_20539_),
    .ZN(alu_out[15])
  );
  AND2_X1 _56314_ (
    .A1(_10604_),
    .A2(_10755_),
    .ZN(_20540_)
  );
  INV_X1 _56315_ (
    .A(_20540_),
    .ZN(_20541_)
  );
  AND2_X1 _56316_ (
    .A1(instr_sub),
    .A2(_10758_),
    .ZN(_20542_)
  );
  AND2_X1 _56317_ (
    .A1(_20541_),
    .A2(_20542_),
    .ZN(_20543_)
  );
  INV_X1 _56318_ (
    .A(_20543_),
    .ZN(_20544_)
  );
  AND2_X1 _56319_ (
    .A1(_10867_),
    .A2(_10891_),
    .ZN(_20545_)
  );
  AND2_X1 _56320_ (
    .A1(_10969_),
    .A2(_20545_),
    .ZN(_20546_)
  );
  AND2_X1 _56321_ (
    .A1(_20424_),
    .A2(_20546_),
    .ZN(_20547_)
  );
  INV_X1 _56322_ (
    .A(_20547_),
    .ZN(_20548_)
  );
  AND2_X1 _56323_ (
    .A1(_10864_),
    .A2(_10888_),
    .ZN(_20549_)
  );
  INV_X1 _56324_ (
    .A(_20549_),
    .ZN(_20550_)
  );
  AND2_X1 _56325_ (
    .A1(_10866_),
    .A2(_20550_),
    .ZN(_20551_)
  );
  INV_X1 _56326_ (
    .A(_20551_),
    .ZN(_20552_)
  );
  AND2_X1 _56327_ (
    .A1(_10968_),
    .A2(_20484_),
    .ZN(_20553_)
  );
  AND2_X1 _56328_ (
    .A1(_20545_),
    .A2(_20553_),
    .ZN(_20554_)
  );
  INV_X1 _56329_ (
    .A(_20554_),
    .ZN(_20555_)
  );
  AND2_X1 _56330_ (
    .A1(_20552_),
    .A2(_20555_),
    .ZN(_20556_)
  );
  AND2_X1 _56331_ (
    .A1(_20548_),
    .A2(_20556_),
    .ZN(_20557_)
  );
  INV_X1 _56332_ (
    .A(_20557_),
    .ZN(_20558_)
  );
  AND2_X1 _56333_ (
    .A1(_10946_),
    .A2(_20557_),
    .ZN(_20559_)
  );
  INV_X1 _56334_ (
    .A(_20559_),
    .ZN(_20560_)
  );
  AND2_X1 _56335_ (
    .A1(_10945_),
    .A2(_20558_),
    .ZN(_20561_)
  );
  INV_X1 _56336_ (
    .A(_20561_),
    .ZN(_20562_)
  );
  AND2_X1 _56337_ (
    .A1(_20560_),
    .A2(_20562_),
    .ZN(_20563_)
  );
  AND2_X1 _56338_ (
    .A1(_21049_),
    .A2(_20563_),
    .ZN(_20564_)
  );
  INV_X1 _56339_ (
    .A(_20564_),
    .ZN(_20565_)
  );
  AND2_X1 _56340_ (
    .A1(_20544_),
    .A2(_20565_),
    .ZN(_20566_)
  );
  INV_X1 _56341_ (
    .A(_20566_),
    .ZN(_20567_)
  );
  AND2_X1 _56342_ (
    .A1(is_lui_auipc_jal_jalr_addi_add_sub),
    .A2(_20567_),
    .ZN(_20568_)
  );
  INV_X1 _56343_ (
    .A(_20568_),
    .ZN(_20569_)
  );
  AND2_X1 _56344_ (
    .A1(_22528_),
    .A2(_10945_),
    .ZN(_20570_)
  );
  INV_X1 _56345_ (
    .A(_20570_),
    .ZN(_20571_)
  );
  AND2_X1 _56346_ (
    .A1(_10941_),
    .A2(_20097_),
    .ZN(_20572_)
  );
  INV_X1 _56347_ (
    .A(_20572_),
    .ZN(_20573_)
  );
  AND2_X1 _56348_ (
    .A1(_22532_),
    .A2(_10944_),
    .ZN(_20574_)
  );
  INV_X1 _56349_ (
    .A(_20574_),
    .ZN(_20575_)
  );
  AND2_X1 _56350_ (
    .A1(_20573_),
    .A2(_20575_),
    .ZN(_20576_)
  );
  AND2_X1 _56351_ (
    .A1(_20571_),
    .A2(_20576_),
    .ZN(_20577_)
  );
  AND2_X1 _56352_ (
    .A1(_20569_),
    .A2(_20577_),
    .ZN(_20578_)
  );
  INV_X1 _56353_ (
    .A(_20578_),
    .ZN(alu_out[16])
  );
  AND2_X1 _56354_ (
    .A1(_10596_),
    .A2(_10598_),
    .ZN(_20579_)
  );
  INV_X1 _56355_ (
    .A(_20579_),
    .ZN(_20580_)
  );
  AND2_X1 _56356_ (
    .A1(_10760_),
    .A2(_20579_),
    .ZN(_20581_)
  );
  INV_X1 _56357_ (
    .A(_20581_),
    .ZN(_20582_)
  );
  AND2_X1 _56358_ (
    .A1(_10759_),
    .A2(_20580_),
    .ZN(_20583_)
  );
  INV_X1 _56359_ (
    .A(_20583_),
    .ZN(_20584_)
  );
  AND2_X1 _56360_ (
    .A1(instr_sub),
    .A2(_20584_),
    .ZN(_20585_)
  );
  AND2_X1 _56361_ (
    .A1(_20582_),
    .A2(_20585_),
    .ZN(_20586_)
  );
  INV_X1 _56362_ (
    .A(_20586_),
    .ZN(_20587_)
  );
  AND2_X1 _56363_ (
    .A1(_10942_),
    .A2(_20562_),
    .ZN(_20588_)
  );
  INV_X1 _56364_ (
    .A(_20588_),
    .ZN(_20589_)
  );
  AND2_X1 _56365_ (
    .A1(_10958_),
    .A2(_20588_),
    .ZN(_20590_)
  );
  INV_X1 _56366_ (
    .A(_20590_),
    .ZN(_20591_)
  );
  AND2_X1 _56367_ (
    .A1(_10957_),
    .A2(_20589_),
    .ZN(_20592_)
  );
  INV_X1 _56368_ (
    .A(_20592_),
    .ZN(_20593_)
  );
  AND2_X1 _56369_ (
    .A1(_20591_),
    .A2(_20593_),
    .ZN(_20594_)
  );
  AND2_X1 _56370_ (
    .A1(_21049_),
    .A2(_20594_),
    .ZN(_20595_)
  );
  INV_X1 _56371_ (
    .A(_20595_),
    .ZN(_20596_)
  );
  AND2_X1 _56372_ (
    .A1(_20587_),
    .A2(_20596_),
    .ZN(_20597_)
  );
  INV_X1 _56373_ (
    .A(_20597_),
    .ZN(_20598_)
  );
  AND2_X1 _56374_ (
    .A1(is_lui_auipc_jal_jalr_addi_add_sub),
    .A2(_20598_),
    .ZN(_20599_)
  );
  INV_X1 _56375_ (
    .A(_20599_),
    .ZN(_20600_)
  );
  AND2_X1 _56376_ (
    .A1(_22528_),
    .A2(_10957_),
    .ZN(_20601_)
  );
  INV_X1 _56377_ (
    .A(_20601_),
    .ZN(_20602_)
  );
  AND2_X1 _56378_ (
    .A1(_10953_),
    .A2(_20097_),
    .ZN(_20603_)
  );
  INV_X1 _56379_ (
    .A(_20603_),
    .ZN(_20604_)
  );
  AND2_X1 _56380_ (
    .A1(_22532_),
    .A2(_10956_),
    .ZN(_20605_)
  );
  INV_X1 _56381_ (
    .A(_20605_),
    .ZN(_20606_)
  );
  AND2_X1 _56382_ (
    .A1(_20604_),
    .A2(_20606_),
    .ZN(_20607_)
  );
  AND2_X1 _56383_ (
    .A1(_20602_),
    .A2(_20607_),
    .ZN(_20608_)
  );
  AND2_X1 _56384_ (
    .A1(_20600_),
    .A2(_20608_),
    .ZN(_20609_)
  );
  INV_X1 _56385_ (
    .A(_20609_),
    .ZN(alu_out[17])
  );
  AND2_X1 _56386_ (
    .A1(_10594_),
    .A2(_10765_),
    .ZN(_20610_)
  );
  INV_X1 _56387_ (
    .A(_20610_),
    .ZN(_20611_)
  );
  AND2_X1 _56388_ (
    .A1(_10954_),
    .A2(_20588_),
    .ZN(_20612_)
  );
  INV_X1 _56389_ (
    .A(_20612_),
    .ZN(_20613_)
  );
  AND2_X1 _56390_ (
    .A1(_10956_),
    .A2(_20589_),
    .ZN(_20614_)
  );
  INV_X1 _56391_ (
    .A(_20614_),
    .ZN(_20615_)
  );
  AND2_X1 _56392_ (
    .A1(_10956_),
    .A2(_20613_),
    .ZN(_20616_)
  );
  AND2_X1 _56393_ (
    .A1(_10954_),
    .A2(_20615_),
    .ZN(_20617_)
  );
  AND2_X1 _56394_ (
    .A1(_10916_),
    .A2(_20617_),
    .ZN(_20618_)
  );
  INV_X1 _56395_ (
    .A(_20618_),
    .ZN(_20619_)
  );
  AND2_X1 _56396_ (
    .A1(_10915_),
    .A2(_20616_),
    .ZN(_20620_)
  );
  INV_X1 _56397_ (
    .A(_20620_),
    .ZN(_20621_)
  );
  AND2_X1 _56398_ (
    .A1(_21049_),
    .A2(_20621_),
    .ZN(_20622_)
  );
  AND2_X1 _56399_ (
    .A1(_20619_),
    .A2(_20622_),
    .ZN(_20623_)
  );
  INV_X1 _56400_ (
    .A(_20623_),
    .ZN(_20624_)
  );
  AND2_X1 _56401_ (
    .A1(instr_sub),
    .A2(_10768_),
    .ZN(_20625_)
  );
  AND2_X1 _56402_ (
    .A1(_20611_),
    .A2(_20625_),
    .ZN(_20626_)
  );
  INV_X1 _56403_ (
    .A(_20626_),
    .ZN(_20627_)
  );
  AND2_X1 _56404_ (
    .A1(_20624_),
    .A2(_20627_),
    .ZN(_20628_)
  );
  INV_X1 _56405_ (
    .A(_20628_),
    .ZN(_20629_)
  );
  AND2_X1 _56406_ (
    .A1(is_lui_auipc_jal_jalr_addi_add_sub),
    .A2(_20629_),
    .ZN(_20630_)
  );
  INV_X1 _56407_ (
    .A(_20630_),
    .ZN(_20631_)
  );
  AND2_X1 _56408_ (
    .A1(_22528_),
    .A2(_10915_),
    .ZN(_20632_)
  );
  INV_X1 _56409_ (
    .A(_20632_),
    .ZN(_20633_)
  );
  AND2_X1 _56410_ (
    .A1(_22532_),
    .A2(_10914_),
    .ZN(_20634_)
  );
  INV_X1 _56411_ (
    .A(_20634_),
    .ZN(_20635_)
  );
  AND2_X1 _56412_ (
    .A1(_10911_),
    .A2(_20097_),
    .ZN(_20636_)
  );
  INV_X1 _56413_ (
    .A(_20636_),
    .ZN(_20637_)
  );
  AND2_X1 _56414_ (
    .A1(_20635_),
    .A2(_20637_),
    .ZN(_20638_)
  );
  AND2_X1 _56415_ (
    .A1(_20633_),
    .A2(_20638_),
    .ZN(_20639_)
  );
  AND2_X1 _56416_ (
    .A1(_20631_),
    .A2(_20639_),
    .ZN(_20640_)
  );
  INV_X1 _56417_ (
    .A(_20640_),
    .ZN(alu_out[18])
  );
  AND2_X1 _56418_ (
    .A1(_10586_),
    .A2(_10588_),
    .ZN(_20641_)
  );
  INV_X1 _56419_ (
    .A(_20641_),
    .ZN(_20642_)
  );
  AND2_X1 _56420_ (
    .A1(_10769_),
    .A2(_20642_),
    .ZN(_20643_)
  );
  INV_X1 _56421_ (
    .A(_20643_),
    .ZN(_20644_)
  );
  AND2_X1 _56422_ (
    .A1(_10770_),
    .A2(_20641_),
    .ZN(_20645_)
  );
  INV_X1 _56423_ (
    .A(_20645_),
    .ZN(_20646_)
  );
  AND2_X1 _56424_ (
    .A1(_20644_),
    .A2(_20646_),
    .ZN(_20647_)
  );
  AND2_X1 _56425_ (
    .A1(instr_sub),
    .A2(_20647_),
    .ZN(_20648_)
  );
  INV_X1 _56426_ (
    .A(_20648_),
    .ZN(_20649_)
  );
  AND2_X1 _56427_ (
    .A1(_10912_),
    .A2(_20621_),
    .ZN(_20650_)
  );
  INV_X1 _56428_ (
    .A(_20650_),
    .ZN(_20651_)
  );
  AND2_X1 _56429_ (
    .A1(_10885_),
    .A2(_20651_),
    .ZN(_20652_)
  );
  INV_X1 _56430_ (
    .A(_20652_),
    .ZN(_20653_)
  );
  AND2_X1 _56431_ (
    .A1(_10886_),
    .A2(_20650_),
    .ZN(_20654_)
  );
  INV_X1 _56432_ (
    .A(_20654_),
    .ZN(_20655_)
  );
  AND2_X1 _56433_ (
    .A1(_21049_),
    .A2(_20655_),
    .ZN(_20656_)
  );
  AND2_X1 _56434_ (
    .A1(_20653_),
    .A2(_20656_),
    .ZN(_20657_)
  );
  INV_X1 _56435_ (
    .A(_20657_),
    .ZN(_20658_)
  );
  AND2_X1 _56436_ (
    .A1(_20649_),
    .A2(_20658_),
    .ZN(_20659_)
  );
  INV_X1 _56437_ (
    .A(_20659_),
    .ZN(_20660_)
  );
  AND2_X1 _56438_ (
    .A1(is_lui_auipc_jal_jalr_addi_add_sub),
    .A2(_20660_),
    .ZN(_20661_)
  );
  INV_X1 _56439_ (
    .A(_20661_),
    .ZN(_20662_)
  );
  AND2_X1 _56440_ (
    .A1(_22528_),
    .A2(_10885_),
    .ZN(_20663_)
  );
  INV_X1 _56441_ (
    .A(_20663_),
    .ZN(_20664_)
  );
  AND2_X1 _56442_ (
    .A1(_10881_),
    .A2(_20097_),
    .ZN(_20665_)
  );
  INV_X1 _56443_ (
    .A(_20665_),
    .ZN(_20666_)
  );
  AND2_X1 _56444_ (
    .A1(_22532_),
    .A2(_10884_),
    .ZN(_20667_)
  );
  INV_X1 _56445_ (
    .A(_20667_),
    .ZN(_20668_)
  );
  AND2_X1 _56446_ (
    .A1(_20666_),
    .A2(_20668_),
    .ZN(_20669_)
  );
  AND2_X1 _56447_ (
    .A1(_20664_),
    .A2(_20669_),
    .ZN(_20670_)
  );
  AND2_X1 _56448_ (
    .A1(_20662_),
    .A2(_20670_),
    .ZN(_20671_)
  );
  INV_X1 _56449_ (
    .A(_20671_),
    .ZN(alu_out[19])
  );
  AND2_X1 _56450_ (
    .A1(_10584_),
    .A2(_10775_),
    .ZN(_20672_)
  );
  INV_X1 _56451_ (
    .A(_20672_),
    .ZN(_20673_)
  );
  AND2_X1 _56452_ (
    .A1(_10884_),
    .A2(_20651_),
    .ZN(_20674_)
  );
  INV_X1 _56453_ (
    .A(_20674_),
    .ZN(_20675_)
  );
  AND2_X1 _56454_ (
    .A1(_10882_),
    .A2(_20650_),
    .ZN(_20676_)
  );
  INV_X1 _56455_ (
    .A(_20676_),
    .ZN(_20677_)
  );
  AND2_X1 _56456_ (
    .A1(_10882_),
    .A2(_20675_),
    .ZN(_20678_)
  );
  AND2_X1 _56457_ (
    .A1(_10884_),
    .A2(_20677_),
    .ZN(_20679_)
  );
  AND2_X1 _56458_ (
    .A1(_11042_),
    .A2(_20678_),
    .ZN(_20680_)
  );
  INV_X1 _56459_ (
    .A(_20680_),
    .ZN(_20681_)
  );
  AND2_X1 _56460_ (
    .A1(_11041_),
    .A2(_20679_),
    .ZN(_20682_)
  );
  INV_X1 _56461_ (
    .A(_20682_),
    .ZN(_20683_)
  );
  AND2_X1 _56462_ (
    .A1(_21049_),
    .A2(_20683_),
    .ZN(_20684_)
  );
  AND2_X1 _56463_ (
    .A1(_20681_),
    .A2(_20684_),
    .ZN(_20685_)
  );
  INV_X1 _56464_ (
    .A(_20685_),
    .ZN(_20686_)
  );
  AND2_X1 _56465_ (
    .A1(instr_sub),
    .A2(_10778_),
    .ZN(_20687_)
  );
  AND2_X1 _56466_ (
    .A1(_20673_),
    .A2(_20687_),
    .ZN(_20688_)
  );
  INV_X1 _56467_ (
    .A(_20688_),
    .ZN(_20689_)
  );
  AND2_X1 _56468_ (
    .A1(_20686_),
    .A2(_20689_),
    .ZN(_20690_)
  );
  INV_X1 _56469_ (
    .A(_20690_),
    .ZN(_20691_)
  );
  AND2_X1 _56470_ (
    .A1(is_lui_auipc_jal_jalr_addi_add_sub),
    .A2(_20691_),
    .ZN(_20692_)
  );
  INV_X1 _56471_ (
    .A(_20692_),
    .ZN(_20693_)
  );
  AND2_X1 _56472_ (
    .A1(_22528_),
    .A2(_11041_),
    .ZN(_20694_)
  );
  INV_X1 _56473_ (
    .A(_20694_),
    .ZN(_20695_)
  );
  AND2_X1 _56474_ (
    .A1(_11037_),
    .A2(_20097_),
    .ZN(_20696_)
  );
  INV_X1 _56475_ (
    .A(_20696_),
    .ZN(_20697_)
  );
  AND2_X1 _56476_ (
    .A1(_22532_),
    .A2(_11040_),
    .ZN(_20698_)
  );
  INV_X1 _56477_ (
    .A(_20698_),
    .ZN(_20699_)
  );
  AND2_X1 _56478_ (
    .A1(_20697_),
    .A2(_20699_),
    .ZN(_20700_)
  );
  AND2_X1 _56479_ (
    .A1(_20695_),
    .A2(_20700_),
    .ZN(_20701_)
  );
  AND2_X1 _56480_ (
    .A1(_20693_),
    .A2(_20701_),
    .ZN(_20702_)
  );
  INV_X1 _56481_ (
    .A(_20702_),
    .ZN(alu_out[20])
  );
  AND2_X1 _56482_ (
    .A1(_10576_),
    .A2(_10578_),
    .ZN(_20703_)
  );
  INV_X1 _56483_ (
    .A(_20703_),
    .ZN(_20704_)
  );
  AND2_X1 _56484_ (
    .A1(_10779_),
    .A2(_20703_),
    .ZN(_20705_)
  );
  INV_X1 _56485_ (
    .A(_20705_),
    .ZN(_20706_)
  );
  AND2_X1 _56486_ (
    .A1(_10780_),
    .A2(_20704_),
    .ZN(_20707_)
  );
  INV_X1 _56487_ (
    .A(_20707_),
    .ZN(_20708_)
  );
  AND2_X1 _56488_ (
    .A1(instr_sub),
    .A2(_20708_),
    .ZN(_20709_)
  );
  AND2_X1 _56489_ (
    .A1(_20706_),
    .A2(_20709_),
    .ZN(_20710_)
  );
  INV_X1 _56490_ (
    .A(_20710_),
    .ZN(_20711_)
  );
  AND2_X1 _56491_ (
    .A1(_11038_),
    .A2(_20683_),
    .ZN(_20712_)
  );
  INV_X1 _56492_ (
    .A(_20712_),
    .ZN(_20713_)
  );
  AND2_X1 _56493_ (
    .A1(_11030_),
    .A2(_20713_),
    .ZN(_20714_)
  );
  INV_X1 _56494_ (
    .A(_20714_),
    .ZN(_20715_)
  );
  AND2_X1 _56495_ (
    .A1(_11029_),
    .A2(_20712_),
    .ZN(_20716_)
  );
  INV_X1 _56496_ (
    .A(_20716_),
    .ZN(_20717_)
  );
  AND2_X1 _56497_ (
    .A1(_20715_),
    .A2(_20717_),
    .ZN(_20718_)
  );
  AND2_X1 _56498_ (
    .A1(_21049_),
    .A2(_20718_),
    .ZN(_20719_)
  );
  INV_X1 _56499_ (
    .A(_20719_),
    .ZN(_20720_)
  );
  AND2_X1 _56500_ (
    .A1(is_lui_auipc_jal_jalr_addi_add_sub),
    .A2(_20711_),
    .ZN(_20721_)
  );
  AND2_X1 _56501_ (
    .A1(_20720_),
    .A2(_20721_),
    .ZN(_20722_)
  );
  INV_X1 _56502_ (
    .A(_20722_),
    .ZN(_20723_)
  );
  AND2_X1 _56503_ (
    .A1(_22528_),
    .A2(_11029_),
    .ZN(_20724_)
  );
  INV_X1 _56504_ (
    .A(_20724_),
    .ZN(_20725_)
  );
  AND2_X1 _56505_ (
    .A1(_11025_),
    .A2(_20097_),
    .ZN(_20726_)
  );
  INV_X1 _56506_ (
    .A(_20726_),
    .ZN(_20727_)
  );
  AND2_X1 _56507_ (
    .A1(_22532_),
    .A2(_11028_),
    .ZN(_20728_)
  );
  INV_X1 _56508_ (
    .A(_20728_),
    .ZN(_20729_)
  );
  AND2_X1 _56509_ (
    .A1(_20727_),
    .A2(_20729_),
    .ZN(_20730_)
  );
  AND2_X1 _56510_ (
    .A1(_20725_),
    .A2(_20730_),
    .ZN(_20731_)
  );
  AND2_X1 _56511_ (
    .A1(_20723_),
    .A2(_20731_),
    .ZN(_20732_)
  );
  INV_X1 _56512_ (
    .A(_20732_),
    .ZN(alu_out[21])
  );
  AND2_X1 _56513_ (
    .A1(_10574_),
    .A2(_10785_),
    .ZN(_20733_)
  );
  INV_X1 _56514_ (
    .A(_20733_),
    .ZN(_20734_)
  );
  AND2_X1 _56515_ (
    .A1(instr_sub),
    .A2(_10788_),
    .ZN(_20735_)
  );
  AND2_X1 _56516_ (
    .A1(_20734_),
    .A2(_20735_),
    .ZN(_20736_)
  );
  INV_X1 _56517_ (
    .A(_20736_),
    .ZN(_20737_)
  );
  AND2_X1 _56518_ (
    .A1(_11026_),
    .A2(_20712_),
    .ZN(_20738_)
  );
  INV_X1 _56519_ (
    .A(_20738_),
    .ZN(_20739_)
  );
  AND2_X1 _56520_ (
    .A1(_11028_),
    .A2(_20713_),
    .ZN(_20740_)
  );
  INV_X1 _56521_ (
    .A(_20740_),
    .ZN(_20741_)
  );
  AND2_X1 _56522_ (
    .A1(_11028_),
    .A2(_20739_),
    .ZN(_20742_)
  );
  AND2_X1 _56523_ (
    .A1(_11026_),
    .A2(_20741_),
    .ZN(_20743_)
  );
  AND2_X1 _56524_ (
    .A1(_10981_),
    .A2(_20742_),
    .ZN(_20744_)
  );
  INV_X1 _56525_ (
    .A(_20744_),
    .ZN(_20745_)
  );
  AND2_X1 _56526_ (
    .A1(_10982_),
    .A2(_20743_),
    .ZN(_20746_)
  );
  INV_X1 _56527_ (
    .A(_20746_),
    .ZN(_20747_)
  );
  AND2_X1 _56528_ (
    .A1(_21049_),
    .A2(_20745_),
    .ZN(_20748_)
  );
  AND2_X1 _56529_ (
    .A1(_20747_),
    .A2(_20748_),
    .ZN(_20749_)
  );
  INV_X1 _56530_ (
    .A(_20749_),
    .ZN(_20750_)
  );
  AND2_X1 _56531_ (
    .A1(_20737_),
    .A2(_20750_),
    .ZN(_20751_)
  );
  INV_X1 _56532_ (
    .A(_20751_),
    .ZN(_20752_)
  );
  AND2_X1 _56533_ (
    .A1(is_lui_auipc_jal_jalr_addi_add_sub),
    .A2(_20752_),
    .ZN(_20753_)
  );
  INV_X1 _56534_ (
    .A(_20753_),
    .ZN(_20754_)
  );
  AND2_X1 _56535_ (
    .A1(_22528_),
    .A2(_10981_),
    .ZN(_20755_)
  );
  INV_X1 _56536_ (
    .A(_20755_),
    .ZN(_20756_)
  );
  AND2_X1 _56537_ (
    .A1(_10977_),
    .A2(_20097_),
    .ZN(_20757_)
  );
  INV_X1 _56538_ (
    .A(_20757_),
    .ZN(_20758_)
  );
  AND2_X1 _56539_ (
    .A1(_22532_),
    .A2(_10980_),
    .ZN(_20759_)
  );
  INV_X1 _56540_ (
    .A(_20759_),
    .ZN(_20760_)
  );
  AND2_X1 _56541_ (
    .A1(_20758_),
    .A2(_20760_),
    .ZN(_20761_)
  );
  AND2_X1 _56542_ (
    .A1(_20756_),
    .A2(_20761_),
    .ZN(_20762_)
  );
  AND2_X1 _56543_ (
    .A1(_20754_),
    .A2(_20762_),
    .ZN(_20763_)
  );
  INV_X1 _56544_ (
    .A(_20763_),
    .ZN(alu_out[22])
  );
  AND2_X1 _56545_ (
    .A1(_10566_),
    .A2(_10568_),
    .ZN(_20764_)
  );
  INV_X1 _56546_ (
    .A(_20764_),
    .ZN(_20765_)
  );
  AND2_X1 _56547_ (
    .A1(_10789_),
    .A2(_20764_),
    .ZN(_20766_)
  );
  INV_X1 _56548_ (
    .A(_20766_),
    .ZN(_20767_)
  );
  AND2_X1 _56549_ (
    .A1(_10790_),
    .A2(_20765_),
    .ZN(_20768_)
  );
  INV_X1 _56550_ (
    .A(_20768_),
    .ZN(_20769_)
  );
  AND2_X1 _56551_ (
    .A1(instr_sub),
    .A2(_20769_),
    .ZN(_20770_)
  );
  AND2_X1 _56552_ (
    .A1(_20767_),
    .A2(_20770_),
    .ZN(_20771_)
  );
  INV_X1 _56553_ (
    .A(_20771_),
    .ZN(_20772_)
  );
  AND2_X1 _56554_ (
    .A1(_10978_),
    .A2(_20745_),
    .ZN(_20773_)
  );
  INV_X1 _56555_ (
    .A(_20773_),
    .ZN(_20774_)
  );
  AND2_X1 _56556_ (
    .A1(_10904_),
    .A2(_20774_),
    .ZN(_20775_)
  );
  INV_X1 _56557_ (
    .A(_20775_),
    .ZN(_20776_)
  );
  AND2_X1 _56558_ (
    .A1(_10903_),
    .A2(_20773_),
    .ZN(_20777_)
  );
  INV_X1 _56559_ (
    .A(_20777_),
    .ZN(_20778_)
  );
  AND2_X1 _56560_ (
    .A1(_20776_),
    .A2(_20778_),
    .ZN(_20779_)
  );
  AND2_X1 _56561_ (
    .A1(_21049_),
    .A2(_20779_),
    .ZN(_20780_)
  );
  INV_X1 _56562_ (
    .A(_20780_),
    .ZN(_20781_)
  );
  AND2_X1 _56563_ (
    .A1(is_lui_auipc_jal_jalr_addi_add_sub),
    .A2(_20772_),
    .ZN(_20782_)
  );
  AND2_X1 _56564_ (
    .A1(_20781_),
    .A2(_20782_),
    .ZN(_20783_)
  );
  INV_X1 _56565_ (
    .A(_20783_),
    .ZN(_20784_)
  );
  AND2_X1 _56566_ (
    .A1(_22528_),
    .A2(_10903_),
    .ZN(_20785_)
  );
  INV_X1 _56567_ (
    .A(_20785_),
    .ZN(_20786_)
  );
  AND2_X1 _56568_ (
    .A1(_10899_),
    .A2(_20097_),
    .ZN(_20787_)
  );
  INV_X1 _56569_ (
    .A(_20787_),
    .ZN(_20788_)
  );
  AND2_X1 _56570_ (
    .A1(_22532_),
    .A2(_10902_),
    .ZN(_20789_)
  );
  INV_X1 _56571_ (
    .A(_20789_),
    .ZN(_20790_)
  );
  AND2_X1 _56572_ (
    .A1(_20788_),
    .A2(_20790_),
    .ZN(_20791_)
  );
  AND2_X1 _56573_ (
    .A1(_20786_),
    .A2(_20791_),
    .ZN(_20792_)
  );
  AND2_X1 _56574_ (
    .A1(_20784_),
    .A2(_20792_),
    .ZN(_20793_)
  );
  INV_X1 _56575_ (
    .A(_20793_),
    .ZN(alu_out[23])
  );
  AND2_X1 _56576_ (
    .A1(_10564_),
    .A2(_10795_),
    .ZN(_20794_)
  );
  INV_X1 _56577_ (
    .A(_20794_),
    .ZN(_20795_)
  );
  AND2_X1 _56578_ (
    .A1(instr_sub),
    .A2(_10798_),
    .ZN(_20796_)
  );
  AND2_X1 _56579_ (
    .A1(_20795_),
    .A2(_20796_),
    .ZN(_20797_)
  );
  INV_X1 _56580_ (
    .A(_20797_),
    .ZN(_20798_)
  );
  AND2_X1 _56581_ (
    .A1(_10900_),
    .A2(_20773_),
    .ZN(_20799_)
  );
  INV_X1 _56582_ (
    .A(_20799_),
    .ZN(_20800_)
  );
  AND2_X1 _56583_ (
    .A1(_10902_),
    .A2(_20774_),
    .ZN(_20801_)
  );
  INV_X1 _56584_ (
    .A(_20801_),
    .ZN(_20802_)
  );
  AND2_X1 _56585_ (
    .A1(_10902_),
    .A2(_20800_),
    .ZN(_20803_)
  );
  AND2_X1 _56586_ (
    .A1(_10900_),
    .A2(_20802_),
    .ZN(_20804_)
  );
  AND2_X1 _56587_ (
    .A1(_10951_),
    .A2(_20803_),
    .ZN(_20805_)
  );
  INV_X1 _56588_ (
    .A(_20805_),
    .ZN(_20806_)
  );
  AND2_X1 _56589_ (
    .A1(_10952_),
    .A2(_20804_),
    .ZN(_20807_)
  );
  INV_X1 _56590_ (
    .A(_20807_),
    .ZN(_20808_)
  );
  AND2_X1 _56591_ (
    .A1(_21049_),
    .A2(_20806_),
    .ZN(_20809_)
  );
  AND2_X1 _56592_ (
    .A1(_20808_),
    .A2(_20809_),
    .ZN(_20810_)
  );
  INV_X1 _56593_ (
    .A(_20810_),
    .ZN(_20811_)
  );
  AND2_X1 _56594_ (
    .A1(_20798_),
    .A2(_20811_),
    .ZN(_20812_)
  );
  INV_X1 _56595_ (
    .A(_20812_),
    .ZN(_20813_)
  );
  AND2_X1 _56596_ (
    .A1(is_lui_auipc_jal_jalr_addi_add_sub),
    .A2(_20813_),
    .ZN(_20814_)
  );
  INV_X1 _56597_ (
    .A(_20814_),
    .ZN(_20815_)
  );
  AND2_X1 _56598_ (
    .A1(_22528_),
    .A2(_10951_),
    .ZN(_20816_)
  );
  INV_X1 _56599_ (
    .A(_20816_),
    .ZN(_20817_)
  );
  AND2_X1 _56600_ (
    .A1(_10947_),
    .A2(_20097_),
    .ZN(_20818_)
  );
  INV_X1 _56601_ (
    .A(_20818_),
    .ZN(_20819_)
  );
  AND2_X1 _56602_ (
    .A1(_22532_),
    .A2(_10950_),
    .ZN(_20820_)
  );
  INV_X1 _56603_ (
    .A(_20820_),
    .ZN(_20821_)
  );
  AND2_X1 _56604_ (
    .A1(_20819_),
    .A2(_20821_),
    .ZN(_20822_)
  );
  AND2_X1 _56605_ (
    .A1(_20817_),
    .A2(_20822_),
    .ZN(_20823_)
  );
  AND2_X1 _56606_ (
    .A1(_20815_),
    .A2(_20823_),
    .ZN(_20824_)
  );
  INV_X1 _56607_ (
    .A(_20824_),
    .ZN(alu_out[24])
  );
  AND2_X1 _56608_ (
    .A1(_10556_),
    .A2(_10558_),
    .ZN(_20825_)
  );
  INV_X1 _56609_ (
    .A(_20825_),
    .ZN(_20826_)
  );
  AND2_X1 _56610_ (
    .A1(_10799_),
    .A2(_20826_),
    .ZN(_20827_)
  );
  INV_X1 _56611_ (
    .A(_20827_),
    .ZN(_20828_)
  );
  AND2_X1 _56612_ (
    .A1(_10800_),
    .A2(_20825_),
    .ZN(_20829_)
  );
  INV_X1 _56613_ (
    .A(_20829_),
    .ZN(_20830_)
  );
  AND2_X1 _56614_ (
    .A1(instr_sub),
    .A2(_20830_),
    .ZN(_20831_)
  );
  AND2_X1 _56615_ (
    .A1(_20828_),
    .A2(_20831_),
    .ZN(_20832_)
  );
  INV_X1 _56616_ (
    .A(_20832_),
    .ZN(_20833_)
  );
  AND2_X1 _56617_ (
    .A1(_10948_),
    .A2(_20806_),
    .ZN(_20834_)
  );
  INV_X1 _56618_ (
    .A(_20834_),
    .ZN(_20835_)
  );
  AND2_X1 _56619_ (
    .A1(_11024_),
    .A2(_20834_),
    .ZN(_20836_)
  );
  INV_X1 _56620_ (
    .A(_20836_),
    .ZN(_20837_)
  );
  AND2_X1 _56621_ (
    .A1(_11023_),
    .A2(_20835_),
    .ZN(_20838_)
  );
  INV_X1 _56622_ (
    .A(_20838_),
    .ZN(_20839_)
  );
  AND2_X1 _56623_ (
    .A1(_20837_),
    .A2(_20839_),
    .ZN(_20840_)
  );
  AND2_X1 _56624_ (
    .A1(_21049_),
    .A2(_20840_),
    .ZN(_20841_)
  );
  INV_X1 _56625_ (
    .A(_20841_),
    .ZN(_20842_)
  );
  AND2_X1 _56626_ (
    .A1(_20833_),
    .A2(_20842_),
    .ZN(_20843_)
  );
  INV_X1 _56627_ (
    .A(_20843_),
    .ZN(_20844_)
  );
  AND2_X1 _56628_ (
    .A1(is_lui_auipc_jal_jalr_addi_add_sub),
    .A2(_20844_),
    .ZN(_20845_)
  );
  INV_X1 _56629_ (
    .A(_20845_),
    .ZN(_20846_)
  );
  AND2_X1 _56630_ (
    .A1(_22528_),
    .A2(_11023_),
    .ZN(_20847_)
  );
  INV_X1 _56631_ (
    .A(_20847_),
    .ZN(_20848_)
  );
  AND2_X1 _56632_ (
    .A1(_11019_),
    .A2(_20097_),
    .ZN(_20849_)
  );
  INV_X1 _56633_ (
    .A(_20849_),
    .ZN(_20850_)
  );
  AND2_X1 _56634_ (
    .A1(_22532_),
    .A2(_11022_),
    .ZN(_20851_)
  );
  INV_X1 _56635_ (
    .A(_20851_),
    .ZN(_20852_)
  );
  AND2_X1 _56636_ (
    .A1(_20850_),
    .A2(_20852_),
    .ZN(_20853_)
  );
  AND2_X1 _56637_ (
    .A1(_20848_),
    .A2(_20853_),
    .ZN(_20854_)
  );
  AND2_X1 _56638_ (
    .A1(_20846_),
    .A2(_20854_),
    .ZN(_20855_)
  );
  INV_X1 _56639_ (
    .A(_20855_),
    .ZN(alu_out[25])
  );
  AND2_X1 _56640_ (
    .A1(_10554_),
    .A2(_10805_),
    .ZN(_20856_)
  );
  INV_X1 _56641_ (
    .A(_20856_),
    .ZN(_20857_)
  );
  AND2_X1 _56642_ (
    .A1(instr_sub),
    .A2(_10808_),
    .ZN(_20858_)
  );
  AND2_X1 _56643_ (
    .A1(_20857_),
    .A2(_20858_),
    .ZN(_20859_)
  );
  INV_X1 _56644_ (
    .A(_20859_),
    .ZN(_20860_)
  );
  AND2_X1 _56645_ (
    .A1(_11022_),
    .A2(_20835_),
    .ZN(_20861_)
  );
  INV_X1 _56646_ (
    .A(_20861_),
    .ZN(_20862_)
  );
  AND2_X1 _56647_ (
    .A1(_11020_),
    .A2(_20834_),
    .ZN(_20863_)
  );
  INV_X1 _56648_ (
    .A(_20863_),
    .ZN(_20864_)
  );
  AND2_X1 _56649_ (
    .A1(_11020_),
    .A2(_20862_),
    .ZN(_20865_)
  );
  AND2_X1 _56650_ (
    .A1(_11022_),
    .A2(_20864_),
    .ZN(_20866_)
  );
  AND2_X1 _56651_ (
    .A1(_11017_),
    .A2(_20866_),
    .ZN(_20867_)
  );
  INV_X1 _56652_ (
    .A(_20867_),
    .ZN(_20868_)
  );
  AND2_X1 _56653_ (
    .A1(_11018_),
    .A2(_20865_),
    .ZN(_20869_)
  );
  INV_X1 _56654_ (
    .A(_20869_),
    .ZN(_20870_)
  );
  AND2_X1 _56655_ (
    .A1(_21049_),
    .A2(_20868_),
    .ZN(_20871_)
  );
  AND2_X1 _56656_ (
    .A1(_20870_),
    .A2(_20871_),
    .ZN(_20872_)
  );
  INV_X1 _56657_ (
    .A(_20872_),
    .ZN(_20873_)
  );
  AND2_X1 _56658_ (
    .A1(_20860_),
    .A2(_20873_),
    .ZN(_20874_)
  );
  INV_X1 _56659_ (
    .A(_20874_),
    .ZN(_20875_)
  );
  AND2_X1 _56660_ (
    .A1(is_lui_auipc_jal_jalr_addi_add_sub),
    .A2(_20875_),
    .ZN(_20876_)
  );
  INV_X1 _56661_ (
    .A(_20876_),
    .ZN(_20877_)
  );
  AND2_X1 _56662_ (
    .A1(_22528_),
    .A2(_11017_),
    .ZN(_20878_)
  );
  INV_X1 _56663_ (
    .A(_20878_),
    .ZN(_20879_)
  );
  AND2_X1 _56664_ (
    .A1(_11013_),
    .A2(_20097_),
    .ZN(_20880_)
  );
  INV_X1 _56665_ (
    .A(_20880_),
    .ZN(_20881_)
  );
  AND2_X1 _56666_ (
    .A1(_22532_),
    .A2(_11016_),
    .ZN(_20882_)
  );
  INV_X1 _56667_ (
    .A(_20882_),
    .ZN(_20883_)
  );
  AND2_X1 _56668_ (
    .A1(_20881_),
    .A2(_20883_),
    .ZN(_20884_)
  );
  AND2_X1 _56669_ (
    .A1(_20879_),
    .A2(_20884_),
    .ZN(_20885_)
  );
  AND2_X1 _56670_ (
    .A1(_20877_),
    .A2(_20885_),
    .ZN(_20886_)
  );
  INV_X1 _56671_ (
    .A(_20886_),
    .ZN(alu_out[26])
  );
  AND2_X1 _56672_ (
    .A1(_10546_),
    .A2(_10548_),
    .ZN(_20887_)
  );
  INV_X1 _56673_ (
    .A(_20887_),
    .ZN(_20888_)
  );
  AND2_X1 _56674_ (
    .A1(_10809_),
    .A2(_20888_),
    .ZN(_20889_)
  );
  INV_X1 _56675_ (
    .A(_20889_),
    .ZN(_20890_)
  );
  AND2_X1 _56676_ (
    .A1(_10810_),
    .A2(_20887_),
    .ZN(_20891_)
  );
  INV_X1 _56677_ (
    .A(_20891_),
    .ZN(_20892_)
  );
  AND2_X1 _56678_ (
    .A1(_20890_),
    .A2(_20892_),
    .ZN(_20893_)
  );
  INV_X1 _56679_ (
    .A(_20893_),
    .ZN(_20894_)
  );
  AND2_X1 _56680_ (
    .A1(instr_sub),
    .A2(_20894_),
    .ZN(_20895_)
  );
  INV_X1 _56681_ (
    .A(_20895_),
    .ZN(_20896_)
  );
  AND2_X1 _56682_ (
    .A1(_11014_),
    .A2(_20868_),
    .ZN(_20897_)
  );
  INV_X1 _56683_ (
    .A(_20897_),
    .ZN(_20898_)
  );
  AND2_X1 _56684_ (
    .A1(_10939_),
    .A2(_20897_),
    .ZN(_20899_)
  );
  INV_X1 _56685_ (
    .A(_20899_),
    .ZN(_20900_)
  );
  AND2_X1 _56686_ (
    .A1(_10940_),
    .A2(_20898_),
    .ZN(_20901_)
  );
  INV_X1 _56687_ (
    .A(_20901_),
    .ZN(_20902_)
  );
  AND2_X1 _56688_ (
    .A1(_21049_),
    .A2(_20902_),
    .ZN(_20903_)
  );
  AND2_X1 _56689_ (
    .A1(_20900_),
    .A2(_20903_),
    .ZN(_20904_)
  );
  INV_X1 _56690_ (
    .A(_20904_),
    .ZN(_20905_)
  );
  AND2_X1 _56691_ (
    .A1(is_lui_auipc_jal_jalr_addi_add_sub),
    .A2(_20905_),
    .ZN(_20906_)
  );
  AND2_X1 _56692_ (
    .A1(_20896_),
    .A2(_20906_),
    .ZN(_20907_)
  );
  INV_X1 _56693_ (
    .A(_20907_),
    .ZN(_20908_)
  );
  AND2_X1 _56694_ (
    .A1(_22528_),
    .A2(_10939_),
    .ZN(_20909_)
  );
  INV_X1 _56695_ (
    .A(_20909_),
    .ZN(_20910_)
  );
  AND2_X1 _56696_ (
    .A1(_22532_),
    .A2(_10938_),
    .ZN(_20911_)
  );
  INV_X1 _56697_ (
    .A(_20911_),
    .ZN(_20912_)
  );
  AND2_X1 _56698_ (
    .A1(_10935_),
    .A2(_20097_),
    .ZN(_20913_)
  );
  INV_X1 _56699_ (
    .A(_20913_),
    .ZN(_20914_)
  );
  AND2_X1 _56700_ (
    .A1(_20912_),
    .A2(_20914_),
    .ZN(_20915_)
  );
  AND2_X1 _56701_ (
    .A1(_20910_),
    .A2(_20915_),
    .ZN(_20916_)
  );
  AND2_X1 _56702_ (
    .A1(_20908_),
    .A2(_20916_),
    .ZN(_20917_)
  );
  INV_X1 _56703_ (
    .A(_20917_),
    .ZN(alu_out[27])
  );
  AND2_X1 _56704_ (
    .A1(_10544_),
    .A2(_10815_),
    .ZN(_20918_)
  );
  INV_X1 _56705_ (
    .A(_20918_),
    .ZN(_20919_)
  );
  AND2_X1 _56706_ (
    .A1(instr_sub),
    .A2(_10818_),
    .ZN(_20920_)
  );
  AND2_X1 _56707_ (
    .A1(_20919_),
    .A2(_20920_),
    .ZN(_20921_)
  );
  INV_X1 _56708_ (
    .A(_20921_),
    .ZN(_20922_)
  );
  AND2_X1 _56709_ (
    .A1(_10938_),
    .A2(_20898_),
    .ZN(_20923_)
  );
  INV_X1 _56710_ (
    .A(_20923_),
    .ZN(_20924_)
  );
  AND2_X1 _56711_ (
    .A1(_10936_),
    .A2(_20897_),
    .ZN(_20925_)
  );
  INV_X1 _56712_ (
    .A(_20925_),
    .ZN(_20926_)
  );
  AND2_X1 _56713_ (
    .A1(_10936_),
    .A2(_20924_),
    .ZN(_20927_)
  );
  AND2_X1 _56714_ (
    .A1(_10938_),
    .A2(_20926_),
    .ZN(_20928_)
  );
  AND2_X1 _56715_ (
    .A1(_10988_),
    .A2(_20927_),
    .ZN(_20929_)
  );
  INV_X1 _56716_ (
    .A(_20929_),
    .ZN(_20930_)
  );
  AND2_X1 _56717_ (
    .A1(_10987_),
    .A2(_20928_),
    .ZN(_20931_)
  );
  INV_X1 _56718_ (
    .A(_20931_),
    .ZN(_20932_)
  );
  AND2_X1 _56719_ (
    .A1(_21049_),
    .A2(_20932_),
    .ZN(_20933_)
  );
  AND2_X1 _56720_ (
    .A1(_20930_),
    .A2(_20933_),
    .ZN(_20934_)
  );
  INV_X1 _56721_ (
    .A(_20934_),
    .ZN(_20935_)
  );
  AND2_X1 _56722_ (
    .A1(_20922_),
    .A2(_20935_),
    .ZN(_20936_)
  );
  INV_X1 _56723_ (
    .A(_20936_),
    .ZN(_20937_)
  );
  AND2_X1 _56724_ (
    .A1(is_lui_auipc_jal_jalr_addi_add_sub),
    .A2(_20937_),
    .ZN(_20938_)
  );
  INV_X1 _56725_ (
    .A(_20938_),
    .ZN(_20939_)
  );
  AND2_X1 _56726_ (
    .A1(_22528_),
    .A2(_10987_),
    .ZN(_20940_)
  );
  INV_X1 _56727_ (
    .A(_20940_),
    .ZN(_20941_)
  );
  AND2_X1 _56728_ (
    .A1(_10983_),
    .A2(_20097_),
    .ZN(_20942_)
  );
  INV_X1 _56729_ (
    .A(_20942_),
    .ZN(_20943_)
  );
  AND2_X1 _56730_ (
    .A1(_22532_),
    .A2(_10986_),
    .ZN(_20944_)
  );
  INV_X1 _56731_ (
    .A(_20944_),
    .ZN(_20945_)
  );
  AND2_X1 _56732_ (
    .A1(_20943_),
    .A2(_20945_),
    .ZN(_20946_)
  );
  AND2_X1 _56733_ (
    .A1(_20941_),
    .A2(_20946_),
    .ZN(_20947_)
  );
  AND2_X1 _56734_ (
    .A1(_20939_),
    .A2(_20947_),
    .ZN(_20948_)
  );
  INV_X1 _56735_ (
    .A(_20948_),
    .ZN(alu_out[28])
  );
  AND2_X1 _56736_ (
    .A1(_10984_),
    .A2(_20932_),
    .ZN(_20949_)
  );
  INV_X1 _56737_ (
    .A(_20949_),
    .ZN(_20950_)
  );
  AND2_X1 _56738_ (
    .A1(_10922_),
    .A2(_20949_),
    .ZN(_20951_)
  );
  INV_X1 _56739_ (
    .A(_20951_),
    .ZN(_20952_)
  );
  AND2_X1 _56740_ (
    .A1(_10921_),
    .A2(_20950_),
    .ZN(_20953_)
  );
  INV_X1 _56741_ (
    .A(_20953_),
    .ZN(_20954_)
  );
  AND2_X1 _56742_ (
    .A1(_20952_),
    .A2(_20954_),
    .ZN(_20955_)
  );
  AND2_X1 _56743_ (
    .A1(_21049_),
    .A2(_20955_),
    .ZN(_20956_)
  );
  INV_X1 _56744_ (
    .A(_20956_),
    .ZN(_20957_)
  );
  AND2_X1 _56745_ (
    .A1(_10540_),
    .A2(_10818_),
    .ZN(_20958_)
  );
  INV_X1 _56746_ (
    .A(_20958_),
    .ZN(_20959_)
  );
  AND2_X1 _56747_ (
    .A1(_10824_),
    .A2(_20959_),
    .ZN(_20960_)
  );
  INV_X1 _56748_ (
    .A(_20960_),
    .ZN(_20961_)
  );
  AND2_X1 _56749_ (
    .A1(_10825_),
    .A2(_20958_),
    .ZN(_20962_)
  );
  INV_X1 _56750_ (
    .A(_20962_),
    .ZN(_20963_)
  );
  AND2_X1 _56751_ (
    .A1(instr_sub),
    .A2(_20963_),
    .ZN(_20964_)
  );
  AND2_X1 _56752_ (
    .A1(_20961_),
    .A2(_20964_),
    .ZN(_20965_)
  );
  INV_X1 _56753_ (
    .A(_20965_),
    .ZN(_20966_)
  );
  AND2_X1 _56754_ (
    .A1(_20957_),
    .A2(_20966_),
    .ZN(_20967_)
  );
  INV_X1 _56755_ (
    .A(_20967_),
    .ZN(_20968_)
  );
  AND2_X1 _56756_ (
    .A1(is_lui_auipc_jal_jalr_addi_add_sub),
    .A2(_20968_),
    .ZN(_20969_)
  );
  INV_X1 _56757_ (
    .A(_20969_),
    .ZN(_20970_)
  );
  AND2_X1 _56758_ (
    .A1(_22528_),
    .A2(_10921_),
    .ZN(_20971_)
  );
  INV_X1 _56759_ (
    .A(_20971_),
    .ZN(_20972_)
  );
  AND2_X1 _56760_ (
    .A1(_10917_),
    .A2(_20097_),
    .ZN(_20973_)
  );
  INV_X1 _56761_ (
    .A(_20973_),
    .ZN(_20974_)
  );
  AND2_X1 _56762_ (
    .A1(_22532_),
    .A2(_10920_),
    .ZN(_20975_)
  );
  INV_X1 _56763_ (
    .A(_20975_),
    .ZN(_20976_)
  );
  AND2_X1 _56764_ (
    .A1(_20974_),
    .A2(_20976_),
    .ZN(_20977_)
  );
  AND2_X1 _56765_ (
    .A1(_20972_),
    .A2(_20977_),
    .ZN(_20978_)
  );
  AND2_X1 _56766_ (
    .A1(_20970_),
    .A2(_20978_),
    .ZN(_20979_)
  );
  INV_X1 _56767_ (
    .A(_20979_),
    .ZN(alu_out[29])
  );
  AND2_X1 _56768_ (
    .A1(_10536_),
    .A2(_10827_),
    .ZN(_20980_)
  );
  INV_X1 _56769_ (
    .A(_20980_),
    .ZN(_20981_)
  );
  AND2_X1 _56770_ (
    .A1(_10920_),
    .A2(_20950_),
    .ZN(_20982_)
  );
  INV_X1 _56771_ (
    .A(_20982_),
    .ZN(_20983_)
  );
  AND2_X1 _56772_ (
    .A1(_10918_),
    .A2(_20949_),
    .ZN(_20984_)
  );
  INV_X1 _56773_ (
    .A(_20984_),
    .ZN(_20985_)
  );
  AND2_X1 _56774_ (
    .A1(_10918_),
    .A2(_20983_),
    .ZN(_20986_)
  );
  AND2_X1 _56775_ (
    .A1(_10920_),
    .A2(_20985_),
    .ZN(_20987_)
  );
  AND2_X1 _56776_ (
    .A1(_10880_),
    .A2(_20986_),
    .ZN(_20988_)
  );
  INV_X1 _56777_ (
    .A(_20988_),
    .ZN(_20989_)
  );
  AND2_X1 _56778_ (
    .A1(_10879_),
    .A2(_20987_),
    .ZN(_20990_)
  );
  INV_X1 _56779_ (
    .A(_20990_),
    .ZN(_20991_)
  );
  AND2_X1 _56780_ (
    .A1(instr_sub),
    .A2(_10829_),
    .ZN(_20992_)
  );
  AND2_X1 _56781_ (
    .A1(_20981_),
    .A2(_20992_),
    .ZN(_20993_)
  );
  INV_X1 _56782_ (
    .A(_20993_),
    .ZN(_20994_)
  );
  AND2_X1 _56783_ (
    .A1(_21049_),
    .A2(_20991_),
    .ZN(_20995_)
  );
  AND2_X1 _56784_ (
    .A1(_20989_),
    .A2(_20995_),
    .ZN(_20996_)
  );
  INV_X1 _56785_ (
    .A(_20996_),
    .ZN(_20997_)
  );
  AND2_X1 _56786_ (
    .A1(_20994_),
    .A2(_20997_),
    .ZN(_20998_)
  );
  INV_X1 _56787_ (
    .A(_20998_),
    .ZN(_20999_)
  );
  AND2_X1 _56788_ (
    .A1(is_lui_auipc_jal_jalr_addi_add_sub),
    .A2(_20999_),
    .ZN(_21000_)
  );
  INV_X1 _56789_ (
    .A(_21000_),
    .ZN(_21001_)
  );
  AND2_X1 _56790_ (
    .A1(_22528_),
    .A2(_10879_),
    .ZN(_21002_)
  );
  INV_X1 _56791_ (
    .A(_21002_),
    .ZN(_21003_)
  );
  AND2_X1 _56792_ (
    .A1(_22532_),
    .A2(_10878_),
    .ZN(_21004_)
  );
  INV_X1 _56793_ (
    .A(_21004_),
    .ZN(_21005_)
  );
  AND2_X1 _56794_ (
    .A1(_10875_),
    .A2(_20097_),
    .ZN(_21006_)
  );
  INV_X1 _56795_ (
    .A(_21006_),
    .ZN(_21007_)
  );
  AND2_X1 _56796_ (
    .A1(_21005_),
    .A2(_21007_),
    .ZN(_21008_)
  );
  AND2_X1 _56797_ (
    .A1(_21003_),
    .A2(_21008_),
    .ZN(_21009_)
  );
  AND2_X1 _56798_ (
    .A1(_21001_),
    .A2(_21009_),
    .ZN(_21010_)
  );
  INV_X1 _56799_ (
    .A(_21010_),
    .ZN(alu_out[30])
  );
  AND2_X1 _56800_ (
    .A1(_10530_),
    .A2(_10831_),
    .ZN(_21011_)
  );
  INV_X1 _56801_ (
    .A(_21011_),
    .ZN(_21012_)
  );
  AND2_X1 _56802_ (
    .A1(instr_sub),
    .A2(_10833_),
    .ZN(_21013_)
  );
  AND2_X1 _56803_ (
    .A1(_21012_),
    .A2(_21013_),
    .ZN(_21014_)
  );
  INV_X1 _56804_ (
    .A(_21014_),
    .ZN(_21015_)
  );
  AND2_X1 _56805_ (
    .A1(_10876_),
    .A2(_20991_),
    .ZN(_21016_)
  );
  INV_X1 _56806_ (
    .A(_21016_),
    .ZN(_21017_)
  );
  AND2_X1 _56807_ (
    .A1(_10999_),
    .A2(_21016_),
    .ZN(_21018_)
  );
  INV_X1 _56808_ (
    .A(_21018_),
    .ZN(_21019_)
  );
  AND2_X1 _56809_ (
    .A1(_11000_),
    .A2(_21017_),
    .ZN(_21020_)
  );
  INV_X1 _56810_ (
    .A(_21020_),
    .ZN(_21021_)
  );
  AND2_X1 _56811_ (
    .A1(_21019_),
    .A2(_21021_),
    .ZN(_21022_)
  );
  AND2_X1 _56812_ (
    .A1(_21049_),
    .A2(_21022_),
    .ZN(_21023_)
  );
  INV_X1 _56813_ (
    .A(_21023_),
    .ZN(_21024_)
  );
  AND2_X1 _56814_ (
    .A1(is_lui_auipc_jal_jalr_addi_add_sub),
    .A2(_21024_),
    .ZN(_21025_)
  );
  AND2_X1 _56815_ (
    .A1(_21015_),
    .A2(_21025_),
    .ZN(_21026_)
  );
  INV_X1 _56816_ (
    .A(_21026_),
    .ZN(_21027_)
  );
  AND2_X1 _56817_ (
    .A1(_22528_),
    .A2(_10999_),
    .ZN(_21028_)
  );
  INV_X1 _56818_ (
    .A(_21028_),
    .ZN(_21029_)
  );
  AND2_X1 _56819_ (
    .A1(_10995_),
    .A2(_20097_),
    .ZN(_21030_)
  );
  INV_X1 _56820_ (
    .A(_21030_),
    .ZN(_21031_)
  );
  AND2_X1 _56821_ (
    .A1(_22532_),
    .A2(_10998_),
    .ZN(_21032_)
  );
  INV_X1 _56822_ (
    .A(_21032_),
    .ZN(_21033_)
  );
  AND2_X1 _56823_ (
    .A1(_21031_),
    .A2(_21033_),
    .ZN(_21034_)
  );
  AND2_X1 _56824_ (
    .A1(_21029_),
    .A2(_21034_),
    .ZN(_21035_)
  );
  AND2_X1 _56825_ (
    .A1(_21027_),
    .A2(_21035_),
    .ZN(_21036_)
  );
  INV_X1 _56826_ (
    .A(_21036_),
    .ZN(alu_out[31])
  );
  BUF_X1 _56827_ (
    .A(\cpuregs[0] [31]),
    .Z(_00526_)
  );
  BUF_X1 _56828_ (
    .A(\cpuregs[0] [0]),
    .Z(_01488_)
  );
  BUF_X1 _56829_ (
    .A(\cpuregs[0] [1]),
    .Z(_01489_)
  );
  BUF_X1 _56830_ (
    .A(\cpuregs[0] [2]),
    .Z(_01490_)
  );
  BUF_X1 _56831_ (
    .A(\cpuregs[0] [3]),
    .Z(_01491_)
  );
  BUF_X1 _56832_ (
    .A(\cpuregs[0] [4]),
    .Z(_01492_)
  );
  BUF_X1 _56833_ (
    .A(\cpuregs[0] [5]),
    .Z(_01493_)
  );
  BUF_X1 _56834_ (
    .A(\cpuregs[0] [6]),
    .Z(_01494_)
  );
  BUF_X1 _56835_ (
    .A(\cpuregs[0] [7]),
    .Z(_01495_)
  );
  BUF_X1 _56836_ (
    .A(\cpuregs[0] [8]),
    .Z(_01496_)
  );
  BUF_X1 _56837_ (
    .A(\cpuregs[0] [9]),
    .Z(_01497_)
  );
  BUF_X1 _56838_ (
    .A(\cpuregs[0] [10]),
    .Z(_01498_)
  );
  BUF_X1 _56839_ (
    .A(\cpuregs[0] [11]),
    .Z(_01499_)
  );
  BUF_X1 _56840_ (
    .A(\cpuregs[0] [12]),
    .Z(_01500_)
  );
  BUF_X1 _56841_ (
    .A(\cpuregs[0] [13]),
    .Z(_01501_)
  );
  BUF_X1 _56842_ (
    .A(\cpuregs[0] [14]),
    .Z(_01502_)
  );
  BUF_X1 _56843_ (
    .A(\cpuregs[0] [15]),
    .Z(_01503_)
  );
  BUF_X1 _56844_ (
    .A(\cpuregs[0] [16]),
    .Z(_01504_)
  );
  BUF_X1 _56845_ (
    .A(\cpuregs[0] [17]),
    .Z(_01505_)
  );
  BUF_X1 _56846_ (
    .A(\cpuregs[0] [18]),
    .Z(_01506_)
  );
  BUF_X1 _56847_ (
    .A(\cpuregs[0] [19]),
    .Z(_01507_)
  );
  BUF_X1 _56848_ (
    .A(\cpuregs[0] [20]),
    .Z(_01508_)
  );
  BUF_X1 _56849_ (
    .A(\cpuregs[0] [21]),
    .Z(_01509_)
  );
  BUF_X1 _56850_ (
    .A(\cpuregs[0] [22]),
    .Z(_01510_)
  );
  BUF_X1 _56851_ (
    .A(\cpuregs[0] [23]),
    .Z(_01511_)
  );
  BUF_X1 _56852_ (
    .A(\cpuregs[0] [24]),
    .Z(_01512_)
  );
  BUF_X1 _56853_ (
    .A(\cpuregs[0] [25]),
    .Z(_01513_)
  );
  BUF_X1 _56854_ (
    .A(\cpuregs[0] [26]),
    .Z(_01514_)
  );
  BUF_X1 _56855_ (
    .A(\cpuregs[0] [27]),
    .Z(_01515_)
  );
  BUF_X1 _56856_ (
    .A(\cpuregs[0] [28]),
    .Z(_01516_)
  );
  BUF_X1 _56857_ (
    .A(\cpuregs[0] [29]),
    .Z(_01517_)
  );
  BUF_X1 _56858_ (
    .A(\cpuregs[0] [30]),
    .Z(_01518_)
  );
  AND2_X1 _56859_ (
    .A1(_11664_),
    .A2(_11666_),
    .ZN(_00048_)
  );
  AND2_X1 _56860_ (
    .A1(_11668_),
    .A2(_11670_),
    .ZN(_00049_)
  );
  AND2_X1 _56861_ (
    .A1(_11672_),
    .A2(_11674_),
    .ZN(_00050_)
  );
  AND2_X1 _56862_ (
    .A1(_11676_),
    .A2(_11678_),
    .ZN(_00051_)
  );
  AND2_X1 _56863_ (
    .A1(_18163_),
    .A2(_18165_),
    .ZN(_00052_)
  );
  AND2_X1 _56864_ (
    .A1(_18185_),
    .A2(_18187_),
    .ZN(_00053_)
  );
  AND2_X1 _56865_ (
    .A1(_18189_),
    .A2(_18191_),
    .ZN(_00054_)
  );
  AND2_X1 _56866_ (
    .A1(_18193_),
    .A2(_18195_),
    .ZN(_00055_)
  );
  AND2_X1 _56867_ (
    .A1(_18177_),
    .A2(_18179_),
    .ZN(_00056_)
  );
  AND2_X1 _56868_ (
    .A1(_18181_),
    .A2(_18183_),
    .ZN(_00057_)
  );
  DFF_X1 _56869__reg (
    .CK(clk),
    .D(_00048_),
    .Q(_00007_[0]),
    .QN(_29069_)
  );
  DFF_X1 _56870__reg (
    .CK(clk),
    .D(_00049_),
    .Q(_00007_[1]),
    .QN(_29070_)
  );
  DFF_X1 _56871__reg (
    .CK(clk),
    .D(_00050_),
    .Q(_00007_[2]),
    .QN(_29071_)
  );
  DFF_X1 _56872__reg (
    .CK(clk),
    .D(_00051_),
    .Q(_00007_[3]),
    .QN(_29072_)
  );
  DFF_X1 _56873__reg (
    .CK(clk),
    .D(_00052_),
    .Q(_00007_[4]),
    .QN(_29039_)
  );
  DFF_X1 _56874__reg (
    .CK(clk),
    .D(_00053_),
    .Q(_00008_[0]),
    .QN(_29074_)
  );
  DFF_X1 _56875__reg (
    .CK(clk),
    .D(_00054_),
    .Q(_00008_[1]),
    .QN(_29075_)
  );
  DFF_X1 _56876__reg (
    .CK(clk),
    .D(_00055_),
    .Q(_00008_[2]),
    .QN(_29076_)
  );
  DFF_X1 _56877__reg (
    .CK(clk),
    .D(_00056_),
    .Q(_00008_[3]),
    .QN(_29077_)
  );
  DFF_X1 _56878__reg (
    .CK(clk),
    .D(_00057_),
    .Q(_00008_[4]),
    .QN(_28976_)
  );
  DFF_X1 alu_out_q_reg_0_  (
    .CK(clk),
    .D(alu_out[0]),
    .Q(alu_out_q[0]),
    .QN(_29112_)
  );
  DFF_X1 alu_out_q_reg_10_  (
    .CK(clk),
    .D(alu_out[10]),
    .Q(alu_out_q[10]),
    .QN(_29122_)
  );
  DFF_X1 alu_out_q_reg_11_  (
    .CK(clk),
    .D(alu_out[11]),
    .Q(alu_out_q[11]),
    .QN(_29123_)
  );
  DFF_X1 alu_out_q_reg_12_  (
    .CK(clk),
    .D(alu_out[12]),
    .Q(alu_out_q[12]),
    .QN(_29124_)
  );
  DFF_X1 alu_out_q_reg_13_  (
    .CK(clk),
    .D(alu_out[13]),
    .Q(alu_out_q[13]),
    .QN(_29125_)
  );
  DFF_X1 alu_out_q_reg_14_  (
    .CK(clk),
    .D(alu_out[14]),
    .Q(alu_out_q[14]),
    .QN(_29126_)
  );
  DFF_X1 alu_out_q_reg_15_  (
    .CK(clk),
    .D(alu_out[15]),
    .Q(alu_out_q[15]),
    .QN(_29127_)
  );
  DFF_X1 alu_out_q_reg_16_  (
    .CK(clk),
    .D(alu_out[16]),
    .Q(alu_out_q[16]),
    .QN(_29128_)
  );
  DFF_X1 alu_out_q_reg_17_  (
    .CK(clk),
    .D(alu_out[17]),
    .Q(alu_out_q[17]),
    .QN(_29129_)
  );
  DFF_X1 alu_out_q_reg_18_  (
    .CK(clk),
    .D(alu_out[18]),
    .Q(alu_out_q[18]),
    .QN(_29130_)
  );
  DFF_X1 alu_out_q_reg_19_  (
    .CK(clk),
    .D(alu_out[19]),
    .Q(alu_out_q[19]),
    .QN(_29131_)
  );
  DFF_X1 alu_out_q_reg_1_  (
    .CK(clk),
    .D(alu_out[1]),
    .Q(alu_out_q[1]),
    .QN(_29113_)
  );
  DFF_X1 alu_out_q_reg_20_  (
    .CK(clk),
    .D(alu_out[20]),
    .Q(alu_out_q[20]),
    .QN(_29132_)
  );
  DFF_X1 alu_out_q_reg_21_  (
    .CK(clk),
    .D(alu_out[21]),
    .Q(alu_out_q[21]),
    .QN(_29133_)
  );
  DFF_X1 alu_out_q_reg_22_  (
    .CK(clk),
    .D(alu_out[22]),
    .Q(alu_out_q[22]),
    .QN(_29134_)
  );
  DFF_X1 alu_out_q_reg_23_  (
    .CK(clk),
    .D(alu_out[23]),
    .Q(alu_out_q[23]),
    .QN(_29135_)
  );
  DFF_X1 alu_out_q_reg_24_  (
    .CK(clk),
    .D(alu_out[24]),
    .Q(alu_out_q[24]),
    .QN(_29136_)
  );
  DFF_X1 alu_out_q_reg_25_  (
    .CK(clk),
    .D(alu_out[25]),
    .Q(alu_out_q[25]),
    .QN(_29137_)
  );
  DFF_X1 alu_out_q_reg_26_  (
    .CK(clk),
    .D(alu_out[26]),
    .Q(alu_out_q[26]),
    .QN(_29138_)
  );
  DFF_X1 alu_out_q_reg_27_  (
    .CK(clk),
    .D(alu_out[27]),
    .Q(alu_out_q[27]),
    .QN(_29139_)
  );
  DFF_X1 alu_out_q_reg_28_  (
    .CK(clk),
    .D(alu_out[28]),
    .Q(alu_out_q[28]),
    .QN(_29140_)
  );
  DFF_X1 alu_out_q_reg_29_  (
    .CK(clk),
    .D(alu_out[29]),
    .Q(alu_out_q[29]),
    .QN(_29141_)
  );
  DFF_X1 alu_out_q_reg_2_  (
    .CK(clk),
    .D(alu_out[2]),
    .Q(alu_out_q[2]),
    .QN(_29114_)
  );
  DFF_X1 alu_out_q_reg_30_  (
    .CK(clk),
    .D(alu_out[30]),
    .Q(alu_out_q[30]),
    .QN(_29142_)
  );
  DFF_X1 alu_out_q_reg_31_  (
    .CK(clk),
    .D(alu_out[31]),
    .Q(alu_out_q[31]),
    .QN(_28822_)
  );
  DFF_X1 alu_out_q_reg_3_  (
    .CK(clk),
    .D(alu_out[3]),
    .Q(alu_out_q[3]),
    .QN(_29115_)
  );
  DFF_X1 alu_out_q_reg_4_  (
    .CK(clk),
    .D(alu_out[4]),
    .Q(alu_out_q[4]),
    .QN(_29116_)
  );
  DFF_X1 alu_out_q_reg_5_  (
    .CK(clk),
    .D(alu_out[5]),
    .Q(alu_out_q[5]),
    .QN(_29117_)
  );
  DFF_X1 alu_out_q_reg_6_  (
    .CK(clk),
    .D(alu_out[6]),
    .Q(alu_out_q[6]),
    .QN(_29118_)
  );
  DFF_X1 alu_out_q_reg_7_  (
    .CK(clk),
    .D(alu_out[7]),
    .Q(alu_out_q[7]),
    .QN(_29119_)
  );
  DFF_X1 alu_out_q_reg_8_  (
    .CK(clk),
    .D(alu_out[8]),
    .Q(alu_out_q[8]),
    .QN(_29120_)
  );
  DFF_X1 alu_out_q_reg_9_  (
    .CK(clk),
    .D(alu_out[9]),
    .Q(alu_out_q[9]),
    .QN(_29121_)
  );
  DFF_X1 count_cycle_reg_0_  (
    .CK(clk),
    .D(_00216_),
    .Q(count_cycle[0]),
    .QN(_29147_[0])
  );
  DFF_X1 count_cycle_reg_10_  (
    .CK(clk),
    .D(_00226_),
    .Q(count_cycle[10]),
    .QN(_28903_)
  );
  DFF_X1 count_cycle_reg_11_  (
    .CK(clk),
    .D(_00227_),
    .Q(count_cycle[11]),
    .QN(_28902_)
  );
  DFF_X1 count_cycle_reg_12_  (
    .CK(clk),
    .D(_00228_),
    .Q(count_cycle[12]),
    .QN(_28901_)
  );
  DFF_X1 count_cycle_reg_13_  (
    .CK(clk),
    .D(_00229_),
    .Q(count_cycle[13]),
    .QN(_28900_)
  );
  DFF_X1 count_cycle_reg_14_  (
    .CK(clk),
    .D(_00230_),
    .Q(count_cycle[14]),
    .QN(_28899_)
  );
  DFF_X1 count_cycle_reg_15_  (
    .CK(clk),
    .D(_00231_),
    .Q(count_cycle[15]),
    .QN(_28898_)
  );
  DFF_X1 count_cycle_reg_16_  (
    .CK(clk),
    .D(_00232_),
    .Q(count_cycle[16]),
    .QN(_28897_)
  );
  DFF_X1 count_cycle_reg_17_  (
    .CK(clk),
    .D(_00233_),
    .Q(count_cycle[17]),
    .QN(_28896_)
  );
  DFF_X1 count_cycle_reg_18_  (
    .CK(clk),
    .D(_00234_),
    .Q(count_cycle[18]),
    .QN(_28895_)
  );
  DFF_X1 count_cycle_reg_19_  (
    .CK(clk),
    .D(_00235_),
    .Q(count_cycle[19]),
    .QN(_28894_)
  );
  DFF_X1 count_cycle_reg_1_  (
    .CK(clk),
    .D(_00217_),
    .Q(count_cycle[1]),
    .QN(_28912_)
  );
  DFF_X1 count_cycle_reg_20_  (
    .CK(clk),
    .D(_00236_),
    .Q(count_cycle[20]),
    .QN(_28893_)
  );
  DFF_X1 count_cycle_reg_21_  (
    .CK(clk),
    .D(_00237_),
    .Q(count_cycle[21]),
    .QN(_28892_)
  );
  DFF_X1 count_cycle_reg_22_  (
    .CK(clk),
    .D(_00238_),
    .Q(count_cycle[22]),
    .QN(_28891_)
  );
  DFF_X1 count_cycle_reg_23_  (
    .CK(clk),
    .D(_00239_),
    .Q(count_cycle[23]),
    .QN(_28890_)
  );
  DFF_X1 count_cycle_reg_24_  (
    .CK(clk),
    .D(_00240_),
    .Q(count_cycle[24]),
    .QN(_28889_)
  );
  DFF_X1 count_cycle_reg_25_  (
    .CK(clk),
    .D(_00241_),
    .Q(count_cycle[25]),
    .QN(_28888_)
  );
  DFF_X1 count_cycle_reg_26_  (
    .CK(clk),
    .D(_00242_),
    .Q(count_cycle[26]),
    .QN(_28887_)
  );
  DFF_X1 count_cycle_reg_27_  (
    .CK(clk),
    .D(_00243_),
    .Q(count_cycle[27]),
    .QN(_28886_)
  );
  DFF_X1 count_cycle_reg_28_  (
    .CK(clk),
    .D(_00244_),
    .Q(count_cycle[28]),
    .QN(_28885_)
  );
  DFF_X1 count_cycle_reg_29_  (
    .CK(clk),
    .D(_00245_),
    .Q(count_cycle[29]),
    .QN(_28884_)
  );
  DFF_X1 count_cycle_reg_2_  (
    .CK(clk),
    .D(_00218_),
    .Q(count_cycle[2]),
    .QN(_28911_)
  );
  DFF_X1 count_cycle_reg_30_  (
    .CK(clk),
    .D(_00246_),
    .Q(count_cycle[30]),
    .QN(_28883_)
  );
  DFF_X1 count_cycle_reg_31_  (
    .CK(clk),
    .D(_00247_),
    .Q(count_cycle[31]),
    .QN(_28882_)
  );
  DFF_X1 count_cycle_reg_32_  (
    .CK(clk),
    .D(_00248_),
    .Q(count_cycle[32]),
    .QN(_28881_)
  );
  DFF_X1 count_cycle_reg_33_  (
    .CK(clk),
    .D(_00249_),
    .Q(count_cycle[33]),
    .QN(_28880_)
  );
  DFF_X1 count_cycle_reg_34_  (
    .CK(clk),
    .D(_00250_),
    .Q(count_cycle[34]),
    .QN(_28879_)
  );
  DFF_X1 count_cycle_reg_35_  (
    .CK(clk),
    .D(_00251_),
    .Q(count_cycle[35]),
    .QN(_28878_)
  );
  DFF_X1 count_cycle_reg_36_  (
    .CK(clk),
    .D(_00252_),
    .Q(count_cycle[36]),
    .QN(_28877_)
  );
  DFF_X1 count_cycle_reg_37_  (
    .CK(clk),
    .D(_00253_),
    .Q(count_cycle[37]),
    .QN(_28876_)
  );
  DFF_X1 count_cycle_reg_38_  (
    .CK(clk),
    .D(_00254_),
    .Q(count_cycle[38]),
    .QN(_28875_)
  );
  DFF_X1 count_cycle_reg_39_  (
    .CK(clk),
    .D(_00255_),
    .Q(count_cycle[39]),
    .QN(_28874_)
  );
  DFF_X1 count_cycle_reg_3_  (
    .CK(clk),
    .D(_00219_),
    .Q(count_cycle[3]),
    .QN(_28910_)
  );
  DFF_X1 count_cycle_reg_40_  (
    .CK(clk),
    .D(_00256_),
    .Q(count_cycle[40]),
    .QN(_28873_)
  );
  DFF_X1 count_cycle_reg_41_  (
    .CK(clk),
    .D(_00257_),
    .Q(count_cycle[41]),
    .QN(_28872_)
  );
  DFF_X1 count_cycle_reg_42_  (
    .CK(clk),
    .D(_00258_),
    .Q(count_cycle[42]),
    .QN(_28871_)
  );
  DFF_X1 count_cycle_reg_43_  (
    .CK(clk),
    .D(_00259_),
    .Q(count_cycle[43]),
    .QN(_28870_)
  );
  DFF_X1 count_cycle_reg_44_  (
    .CK(clk),
    .D(_00260_),
    .Q(count_cycle[44]),
    .QN(_28869_)
  );
  DFF_X1 count_cycle_reg_45_  (
    .CK(clk),
    .D(_00261_),
    .Q(count_cycle[45]),
    .QN(_28868_)
  );
  DFF_X1 count_cycle_reg_46_  (
    .CK(clk),
    .D(_00262_),
    .Q(count_cycle[46]),
    .QN(_28867_)
  );
  DFF_X1 count_cycle_reg_47_  (
    .CK(clk),
    .D(_00263_),
    .Q(count_cycle[47]),
    .QN(_28866_)
  );
  DFF_X1 count_cycle_reg_48_  (
    .CK(clk),
    .D(_00264_),
    .Q(count_cycle[48]),
    .QN(_28865_)
  );
  DFF_X1 count_cycle_reg_49_  (
    .CK(clk),
    .D(_00265_),
    .Q(count_cycle[49]),
    .QN(_28864_)
  );
  DFF_X1 count_cycle_reg_4_  (
    .CK(clk),
    .D(_00220_),
    .Q(count_cycle[4]),
    .QN(_28909_)
  );
  DFF_X1 count_cycle_reg_50_  (
    .CK(clk),
    .D(_00266_),
    .Q(count_cycle[50]),
    .QN(_28863_)
  );
  DFF_X1 count_cycle_reg_51_  (
    .CK(clk),
    .D(_00267_),
    .Q(count_cycle[51]),
    .QN(_28862_)
  );
  DFF_X1 count_cycle_reg_52_  (
    .CK(clk),
    .D(_00268_),
    .Q(count_cycle[52]),
    .QN(_28861_)
  );
  DFF_X1 count_cycle_reg_53_  (
    .CK(clk),
    .D(_00269_),
    .Q(count_cycle[53]),
    .QN(_28860_)
  );
  DFF_X1 count_cycle_reg_54_  (
    .CK(clk),
    .D(_00270_),
    .Q(count_cycle[54]),
    .QN(_28859_)
  );
  DFF_X1 count_cycle_reg_55_  (
    .CK(clk),
    .D(_00271_),
    .Q(count_cycle[55]),
    .QN(_28858_)
  );
  DFF_X1 count_cycle_reg_56_  (
    .CK(clk),
    .D(_00272_),
    .Q(count_cycle[56]),
    .QN(_28857_)
  );
  DFF_X1 count_cycle_reg_57_  (
    .CK(clk),
    .D(_00273_),
    .Q(count_cycle[57]),
    .QN(_28856_)
  );
  DFF_X1 count_cycle_reg_58_  (
    .CK(clk),
    .D(_00274_),
    .Q(count_cycle[58]),
    .QN(_28855_)
  );
  DFF_X1 count_cycle_reg_59_  (
    .CK(clk),
    .D(_00275_),
    .Q(count_cycle[59]),
    .QN(_28854_)
  );
  DFF_X1 count_cycle_reg_5_  (
    .CK(clk),
    .D(_00221_),
    .Q(count_cycle[5]),
    .QN(_28908_)
  );
  DFF_X1 count_cycle_reg_60_  (
    .CK(clk),
    .D(_00276_),
    .Q(count_cycle[60]),
    .QN(_28853_)
  );
  DFF_X1 count_cycle_reg_61_  (
    .CK(clk),
    .D(_00277_),
    .Q(count_cycle[61]),
    .QN(_28852_)
  );
  DFF_X1 count_cycle_reg_62_  (
    .CK(clk),
    .D(_00278_),
    .Q(count_cycle[62]),
    .QN(_28851_)
  );
  DFF_X1 count_cycle_reg_63_  (
    .CK(clk),
    .D(_00279_),
    .Q(count_cycle[63]),
    .QN(_28850_)
  );
  DFF_X1 count_cycle_reg_6_  (
    .CK(clk),
    .D(_00222_),
    .Q(count_cycle[6]),
    .QN(_28907_)
  );
  DFF_X1 count_cycle_reg_7_  (
    .CK(clk),
    .D(_00223_),
    .Q(count_cycle[7]),
    .QN(_28906_)
  );
  DFF_X1 count_cycle_reg_8_  (
    .CK(clk),
    .D(_00224_),
    .Q(count_cycle[8]),
    .QN(_28905_)
  );
  DFF_X1 count_cycle_reg_9_  (
    .CK(clk),
    .D(_00225_),
    .Q(count_cycle[9]),
    .QN(_28904_)
  );
  DFF_X1 count_instr_reg_0_  (
    .CK(clk),
    .D(_00088_),
    .Q(count_instr[0]),
    .QN(_29148_[0])
  );
  DFF_X1 count_instr_reg_10_  (
    .CK(clk),
    .D(_00098_),
    .Q(count_instr[10]),
    .QN(_29029_)
  );
  DFF_X1 count_instr_reg_11_  (
    .CK(clk),
    .D(_00099_),
    .Q(count_instr[11]),
    .QN(_29028_)
  );
  DFF_X1 count_instr_reg_12_  (
    .CK(clk),
    .D(_00100_),
    .Q(count_instr[12]),
    .QN(_29027_)
  );
  DFF_X1 count_instr_reg_13_  (
    .CK(clk),
    .D(_00101_),
    .Q(count_instr[13]),
    .QN(_29026_)
  );
  DFF_X1 count_instr_reg_14_  (
    .CK(clk),
    .D(_00102_),
    .Q(count_instr[14]),
    .QN(_29025_)
  );
  DFF_X1 count_instr_reg_15_  (
    .CK(clk),
    .D(_00103_),
    .Q(count_instr[15]),
    .QN(_29024_)
  );
  DFF_X1 count_instr_reg_16_  (
    .CK(clk),
    .D(_00104_),
    .Q(count_instr[16]),
    .QN(_29023_)
  );
  DFF_X1 count_instr_reg_17_  (
    .CK(clk),
    .D(_00105_),
    .Q(count_instr[17]),
    .QN(_29022_)
  );
  DFF_X1 count_instr_reg_18_  (
    .CK(clk),
    .D(_00106_),
    .Q(count_instr[18]),
    .QN(_29021_)
  );
  DFF_X1 count_instr_reg_19_  (
    .CK(clk),
    .D(_00107_),
    .Q(count_instr[19]),
    .QN(_29020_)
  );
  DFF_X1 count_instr_reg_1_  (
    .CK(clk),
    .D(_00089_),
    .Q(count_instr[1]),
    .QN(_29038_)
  );
  DFF_X1 count_instr_reg_20_  (
    .CK(clk),
    .D(_00108_),
    .Q(count_instr[20]),
    .QN(_29019_)
  );
  DFF_X1 count_instr_reg_21_  (
    .CK(clk),
    .D(_00109_),
    .Q(count_instr[21]),
    .QN(_29018_)
  );
  DFF_X1 count_instr_reg_22_  (
    .CK(clk),
    .D(_00110_),
    .Q(count_instr[22]),
    .QN(_29017_)
  );
  DFF_X1 count_instr_reg_23_  (
    .CK(clk),
    .D(_00111_),
    .Q(count_instr[23]),
    .QN(_29016_)
  );
  DFF_X1 count_instr_reg_24_  (
    .CK(clk),
    .D(_00112_),
    .Q(count_instr[24]),
    .QN(_29015_)
  );
  DFF_X1 count_instr_reg_25_  (
    .CK(clk),
    .D(_00113_),
    .Q(count_instr[25]),
    .QN(_29014_)
  );
  DFF_X1 count_instr_reg_26_  (
    .CK(clk),
    .D(_00114_),
    .Q(count_instr[26]),
    .QN(_29013_)
  );
  DFF_X1 count_instr_reg_27_  (
    .CK(clk),
    .D(_00115_),
    .Q(count_instr[27]),
    .QN(_29012_)
  );
  DFF_X1 count_instr_reg_28_  (
    .CK(clk),
    .D(_00116_),
    .Q(count_instr[28]),
    .QN(_29011_)
  );
  DFF_X1 count_instr_reg_29_  (
    .CK(clk),
    .D(_00117_),
    .Q(count_instr[29]),
    .QN(_29010_)
  );
  DFF_X1 count_instr_reg_2_  (
    .CK(clk),
    .D(_00090_),
    .Q(count_instr[2]),
    .QN(_29037_)
  );
  DFF_X1 count_instr_reg_30_  (
    .CK(clk),
    .D(_00118_),
    .Q(count_instr[30]),
    .QN(_29009_)
  );
  DFF_X1 count_instr_reg_31_  (
    .CK(clk),
    .D(_00119_),
    .Q(count_instr[31]),
    .QN(_29008_)
  );
  DFF_X1 count_instr_reg_32_  (
    .CK(clk),
    .D(_00120_),
    .Q(count_instr[32]),
    .QN(_29007_)
  );
  DFF_X1 count_instr_reg_33_  (
    .CK(clk),
    .D(_00121_),
    .Q(count_instr[33]),
    .QN(_29006_)
  );
  DFF_X1 count_instr_reg_34_  (
    .CK(clk),
    .D(_00122_),
    .Q(count_instr[34]),
    .QN(_29005_)
  );
  DFF_X1 count_instr_reg_35_  (
    .CK(clk),
    .D(_00123_),
    .Q(count_instr[35]),
    .QN(_29004_)
  );
  DFF_X1 count_instr_reg_36_  (
    .CK(clk),
    .D(_00124_),
    .Q(count_instr[36]),
    .QN(_29003_)
  );
  DFF_X1 count_instr_reg_37_  (
    .CK(clk),
    .D(_00125_),
    .Q(count_instr[37]),
    .QN(_29002_)
  );
  DFF_X1 count_instr_reg_38_  (
    .CK(clk),
    .D(_00126_),
    .Q(count_instr[38]),
    .QN(_29001_)
  );
  DFF_X1 count_instr_reg_39_  (
    .CK(clk),
    .D(_00127_),
    .Q(count_instr[39]),
    .QN(_29000_)
  );
  DFF_X1 count_instr_reg_3_  (
    .CK(clk),
    .D(_00091_),
    .Q(count_instr[3]),
    .QN(_29036_)
  );
  DFF_X1 count_instr_reg_40_  (
    .CK(clk),
    .D(_00128_),
    .Q(count_instr[40]),
    .QN(_28999_)
  );
  DFF_X1 count_instr_reg_41_  (
    .CK(clk),
    .D(_00129_),
    .Q(count_instr[41]),
    .QN(_28998_)
  );
  DFF_X1 count_instr_reg_42_  (
    .CK(clk),
    .D(_00130_),
    .Q(count_instr[42]),
    .QN(_28997_)
  );
  DFF_X1 count_instr_reg_43_  (
    .CK(clk),
    .D(_00131_),
    .Q(count_instr[43]),
    .QN(_28996_)
  );
  DFF_X1 count_instr_reg_44_  (
    .CK(clk),
    .D(_00132_),
    .Q(count_instr[44]),
    .QN(_28995_)
  );
  DFF_X1 count_instr_reg_45_  (
    .CK(clk),
    .D(_00133_),
    .Q(count_instr[45]),
    .QN(_28994_)
  );
  DFF_X1 count_instr_reg_46_  (
    .CK(clk),
    .D(_00134_),
    .Q(count_instr[46]),
    .QN(_28993_)
  );
  DFF_X1 count_instr_reg_47_  (
    .CK(clk),
    .D(_00135_),
    .Q(count_instr[47]),
    .QN(_28992_)
  );
  DFF_X1 count_instr_reg_48_  (
    .CK(clk),
    .D(_00136_),
    .Q(count_instr[48]),
    .QN(_28991_)
  );
  DFF_X1 count_instr_reg_49_  (
    .CK(clk),
    .D(_00137_),
    .Q(count_instr[49]),
    .QN(_28990_)
  );
  DFF_X1 count_instr_reg_4_  (
    .CK(clk),
    .D(_00092_),
    .Q(count_instr[4]),
    .QN(_29035_)
  );
  DFF_X1 count_instr_reg_50_  (
    .CK(clk),
    .D(_00138_),
    .Q(count_instr[50]),
    .QN(_28989_)
  );
  DFF_X1 count_instr_reg_51_  (
    .CK(clk),
    .D(_00139_),
    .Q(count_instr[51]),
    .QN(_28988_)
  );
  DFF_X1 count_instr_reg_52_  (
    .CK(clk),
    .D(_00140_),
    .Q(count_instr[52]),
    .QN(_28987_)
  );
  DFF_X1 count_instr_reg_53_  (
    .CK(clk),
    .D(_00141_),
    .Q(count_instr[53]),
    .QN(_28986_)
  );
  DFF_X1 count_instr_reg_54_  (
    .CK(clk),
    .D(_00142_),
    .Q(count_instr[54]),
    .QN(_28985_)
  );
  DFF_X1 count_instr_reg_55_  (
    .CK(clk),
    .D(_00143_),
    .Q(count_instr[55]),
    .QN(_28984_)
  );
  DFF_X1 count_instr_reg_56_  (
    .CK(clk),
    .D(_00144_),
    .Q(count_instr[56]),
    .QN(_28983_)
  );
  DFF_X1 count_instr_reg_57_  (
    .CK(clk),
    .D(_00145_),
    .Q(count_instr[57]),
    .QN(_28982_)
  );
  DFF_X1 count_instr_reg_58_  (
    .CK(clk),
    .D(_00146_),
    .Q(count_instr[58]),
    .QN(_28981_)
  );
  DFF_X1 count_instr_reg_59_  (
    .CK(clk),
    .D(_00147_),
    .Q(count_instr[59]),
    .QN(_28980_)
  );
  DFF_X1 count_instr_reg_5_  (
    .CK(clk),
    .D(_00093_),
    .Q(count_instr[5]),
    .QN(_29034_)
  );
  DFF_X1 count_instr_reg_60_  (
    .CK(clk),
    .D(_00148_),
    .Q(count_instr[60]),
    .QN(_28979_)
  );
  DFF_X1 count_instr_reg_61_  (
    .CK(clk),
    .D(_00149_),
    .Q(count_instr[61]),
    .QN(_28978_)
  );
  DFF_X1 count_instr_reg_62_  (
    .CK(clk),
    .D(_00150_),
    .Q(count_instr[62]),
    .QN(_28977_)
  );
  DFF_X1 count_instr_reg_63_  (
    .CK(clk),
    .D(_00151_),
    .Q(count_instr[63]),
    .QN(_29073_)
  );
  DFF_X1 count_instr_reg_6_  (
    .CK(clk),
    .D(_00094_),
    .Q(count_instr[6]),
    .QN(_29033_)
  );
  DFF_X1 count_instr_reg_7_  (
    .CK(clk),
    .D(_00095_),
    .Q(count_instr[7]),
    .QN(_29032_)
  );
  DFF_X1 count_instr_reg_8_  (
    .CK(clk),
    .D(_00096_),
    .Q(count_instr[8]),
    .QN(_29031_)
  );
  DFF_X1 count_instr_reg_9_  (
    .CK(clk),
    .D(_00097_),
    .Q(count_instr[9]),
    .QN(_29030_)
  );
  DFF_X1 cpu_state_reg_0_  (
    .CK(clk),
    .D(_01567_),
    .Q(cpu_state[0]),
    .QN(_00016_)
  );
  DFF_X1 cpu_state_reg_1_  (
    .CK(clk),
    .D(_01568_),
    .Q(cpu_state[1]),
    .QN(_00015_)
  );
  DFF_X1 cpu_state_reg_2_  (
    .CK(clk),
    .D(_01569_),
    .Q(cpu_state[2]),
    .QN(_00014_)
  );
  DFF_X1 cpu_state_reg_3_  (
    .CK(clk),
    .D(_01570_),
    .Q(cpu_state[3]),
    .QN(_00013_)
  );
  DFF_X1 cpu_state_reg_4_  (
    .CK(clk),
    .D(_01571_),
    .Q(cpu_state[4]),
    .QN(_00012_)
  );
  DFF_X1 cpu_state_reg_5_  (
    .CK(clk),
    .D(_01572_),
    .Q(cpu_state[5]),
    .QN(_00011_)
  );
  DFF_X1 cpu_state_reg_6_  (
    .CK(clk),
    .D(_01573_),
    .Q(cpu_state[6]),
    .QN(_00010_)
  );
  DFF_X1 cpu_state_reg_7_  (
    .CK(clk),
    .D(_01574_),
    .Q(cpu_state[7]),
    .QN(_00009_)
  );
  DFF_X1 cpuregs_reg_0__0_  (
    .CK(clk),
    .D(_01488_),
    .Q(\cpuregs[0] [0]),
    .QN(_27700_)
  );
  DFF_X1 cpuregs_reg_0__10_  (
    .CK(clk),
    .D(_01498_),
    .Q(\cpuregs[0] [10]),
    .QN(_27690_)
  );
  DFF_X1 cpuregs_reg_0__11_  (
    .CK(clk),
    .D(_01499_),
    .Q(\cpuregs[0] [11]),
    .QN(_27689_)
  );
  DFF_X1 cpuregs_reg_0__12_  (
    .CK(clk),
    .D(_01500_),
    .Q(\cpuregs[0] [12]),
    .QN(_27688_)
  );
  DFF_X1 cpuregs_reg_0__13_  (
    .CK(clk),
    .D(_01501_),
    .Q(\cpuregs[0] [13]),
    .QN(_27687_)
  );
  DFF_X1 cpuregs_reg_0__14_  (
    .CK(clk),
    .D(_01502_),
    .Q(\cpuregs[0] [14]),
    .QN(_27686_)
  );
  DFF_X1 cpuregs_reg_0__15_  (
    .CK(clk),
    .D(_01503_),
    .Q(\cpuregs[0] [15]),
    .QN(_27685_)
  );
  DFF_X1 cpuregs_reg_0__16_  (
    .CK(clk),
    .D(_01504_),
    .Q(\cpuregs[0] [16]),
    .QN(_27684_)
  );
  DFF_X1 cpuregs_reg_0__17_  (
    .CK(clk),
    .D(_01505_),
    .Q(\cpuregs[0] [17]),
    .QN(_27683_)
  );
  DFF_X1 cpuregs_reg_0__18_  (
    .CK(clk),
    .D(_01506_),
    .Q(\cpuregs[0] [18]),
    .QN(_27682_)
  );
  DFF_X1 cpuregs_reg_0__19_  (
    .CK(clk),
    .D(_01507_),
    .Q(\cpuregs[0] [19]),
    .QN(_27681_)
  );
  DFF_X1 cpuregs_reg_0__1_  (
    .CK(clk),
    .D(_01489_),
    .Q(\cpuregs[0] [1]),
    .QN(_27699_)
  );
  DFF_X1 cpuregs_reg_0__20_  (
    .CK(clk),
    .D(_01508_),
    .Q(\cpuregs[0] [20]),
    .QN(_27680_)
  );
  DFF_X1 cpuregs_reg_0__21_  (
    .CK(clk),
    .D(_01509_),
    .Q(\cpuregs[0] [21]),
    .QN(_27679_)
  );
  DFF_X1 cpuregs_reg_0__22_  (
    .CK(clk),
    .D(_01510_),
    .Q(\cpuregs[0] [22]),
    .QN(_27678_)
  );
  DFF_X1 cpuregs_reg_0__23_  (
    .CK(clk),
    .D(_01511_),
    .Q(\cpuregs[0] [23]),
    .QN(_27677_)
  );
  DFF_X1 cpuregs_reg_0__24_  (
    .CK(clk),
    .D(_01512_),
    .Q(\cpuregs[0] [24]),
    .QN(_27676_)
  );
  DFF_X1 cpuregs_reg_0__25_  (
    .CK(clk),
    .D(_01513_),
    .Q(\cpuregs[0] [25]),
    .QN(_27675_)
  );
  DFF_X1 cpuregs_reg_0__26_  (
    .CK(clk),
    .D(_01514_),
    .Q(\cpuregs[0] [26]),
    .QN(_27674_)
  );
  DFF_X1 cpuregs_reg_0__27_  (
    .CK(clk),
    .D(_01515_),
    .Q(\cpuregs[0] [27]),
    .QN(_27673_)
  );
  DFF_X1 cpuregs_reg_0__28_  (
    .CK(clk),
    .D(_01516_),
    .Q(\cpuregs[0] [28]),
    .QN(_27672_)
  );
  DFF_X1 cpuregs_reg_0__29_  (
    .CK(clk),
    .D(_01517_),
    .Q(\cpuregs[0] [29]),
    .QN(_27671_)
  );
  DFF_X1 cpuregs_reg_0__2_  (
    .CK(clk),
    .D(_01490_),
    .Q(\cpuregs[0] [2]),
    .QN(_27698_)
  );
  DFF_X1 cpuregs_reg_0__30_  (
    .CK(clk),
    .D(_01518_),
    .Q(\cpuregs[0] [30]),
    .QN(_27670_)
  );
  DFF_X1 cpuregs_reg_0__31_  (
    .CK(clk),
    .D(_00526_),
    .Q(\cpuregs[0] [31]),
    .QN(_28662_)
  );
  DFF_X1 cpuregs_reg_0__3_  (
    .CK(clk),
    .D(_01491_),
    .Q(\cpuregs[0] [3]),
    .QN(_27697_)
  );
  DFF_X1 cpuregs_reg_0__4_  (
    .CK(clk),
    .D(_01492_),
    .Q(\cpuregs[0] [4]),
    .QN(_27696_)
  );
  DFF_X1 cpuregs_reg_0__5_  (
    .CK(clk),
    .D(_01493_),
    .Q(\cpuregs[0] [5]),
    .QN(_27695_)
  );
  DFF_X1 cpuregs_reg_0__6_  (
    .CK(clk),
    .D(_01494_),
    .Q(\cpuregs[0] [6]),
    .QN(_27694_)
  );
  DFF_X1 cpuregs_reg_0__7_  (
    .CK(clk),
    .D(_01495_),
    .Q(\cpuregs[0] [7]),
    .QN(_27693_)
  );
  DFF_X1 cpuregs_reg_0__8_  (
    .CK(clk),
    .D(_01496_),
    .Q(\cpuregs[0] [8]),
    .QN(_27692_)
  );
  DFF_X1 cpuregs_reg_0__9_  (
    .CK(clk),
    .D(_01497_),
    .Q(\cpuregs[0] [9]),
    .QN(_27691_)
  );
  DFF_X1 cpuregs_reg_10__0_  (
    .CK(clk),
    .D(_01054_),
    .Q(\cpuregs[10] [0]),
    .QN(_28134_)
  );
  DFF_X1 cpuregs_reg_10__10_  (
    .CK(clk),
    .D(_01064_),
    .Q(\cpuregs[10] [10]),
    .QN(_28124_)
  );
  DFF_X1 cpuregs_reg_10__11_  (
    .CK(clk),
    .D(_01065_),
    .Q(\cpuregs[10] [11]),
    .QN(_28123_)
  );
  DFF_X1 cpuregs_reg_10__12_  (
    .CK(clk),
    .D(_01066_),
    .Q(\cpuregs[10] [12]),
    .QN(_28122_)
  );
  DFF_X1 cpuregs_reg_10__13_  (
    .CK(clk),
    .D(_01067_),
    .Q(\cpuregs[10] [13]),
    .QN(_28121_)
  );
  DFF_X1 cpuregs_reg_10__14_  (
    .CK(clk),
    .D(_01068_),
    .Q(\cpuregs[10] [14]),
    .QN(_28120_)
  );
  DFF_X1 cpuregs_reg_10__15_  (
    .CK(clk),
    .D(_01069_),
    .Q(\cpuregs[10] [15]),
    .QN(_28119_)
  );
  DFF_X1 cpuregs_reg_10__16_  (
    .CK(clk),
    .D(_01070_),
    .Q(\cpuregs[10] [16]),
    .QN(_28118_)
  );
  DFF_X1 cpuregs_reg_10__17_  (
    .CK(clk),
    .D(_01071_),
    .Q(\cpuregs[10] [17]),
    .QN(_28117_)
  );
  DFF_X1 cpuregs_reg_10__18_  (
    .CK(clk),
    .D(_01072_),
    .Q(\cpuregs[10] [18]),
    .QN(_28116_)
  );
  DFF_X1 cpuregs_reg_10__19_  (
    .CK(clk),
    .D(_01073_),
    .Q(\cpuregs[10] [19]),
    .QN(_28115_)
  );
  DFF_X1 cpuregs_reg_10__1_  (
    .CK(clk),
    .D(_01055_),
    .Q(\cpuregs[10] [1]),
    .QN(_28133_)
  );
  DFF_X1 cpuregs_reg_10__20_  (
    .CK(clk),
    .D(_01074_),
    .Q(\cpuregs[10] [20]),
    .QN(_28114_)
  );
  DFF_X1 cpuregs_reg_10__21_  (
    .CK(clk),
    .D(_01075_),
    .Q(\cpuregs[10] [21]),
    .QN(_28113_)
  );
  DFF_X1 cpuregs_reg_10__22_  (
    .CK(clk),
    .D(_01076_),
    .Q(\cpuregs[10] [22]),
    .QN(_28112_)
  );
  DFF_X1 cpuregs_reg_10__23_  (
    .CK(clk),
    .D(_01077_),
    .Q(\cpuregs[10] [23]),
    .QN(_28111_)
  );
  DFF_X1 cpuregs_reg_10__24_  (
    .CK(clk),
    .D(_01078_),
    .Q(\cpuregs[10] [24]),
    .QN(_28110_)
  );
  DFF_X1 cpuregs_reg_10__25_  (
    .CK(clk),
    .D(_01079_),
    .Q(\cpuregs[10] [25]),
    .QN(_28109_)
  );
  DFF_X1 cpuregs_reg_10__26_  (
    .CK(clk),
    .D(_01080_),
    .Q(\cpuregs[10] [26]),
    .QN(_28108_)
  );
  DFF_X1 cpuregs_reg_10__27_  (
    .CK(clk),
    .D(_01081_),
    .Q(\cpuregs[10] [27]),
    .QN(_28107_)
  );
  DFF_X1 cpuregs_reg_10__28_  (
    .CK(clk),
    .D(_01082_),
    .Q(\cpuregs[10] [28]),
    .QN(_28106_)
  );
  DFF_X1 cpuregs_reg_10__29_  (
    .CK(clk),
    .D(_01083_),
    .Q(\cpuregs[10] [29]),
    .QN(_28105_)
  );
  DFF_X1 cpuregs_reg_10__2_  (
    .CK(clk),
    .D(_01056_),
    .Q(\cpuregs[10] [2]),
    .QN(_28132_)
  );
  DFF_X1 cpuregs_reg_10__30_  (
    .CK(clk),
    .D(_01084_),
    .Q(\cpuregs[10] [30]),
    .QN(_28104_)
  );
  DFF_X1 cpuregs_reg_10__31_  (
    .CK(clk),
    .D(_00525_),
    .Q(\cpuregs[10] [31]),
    .QN(_28663_)
  );
  DFF_X1 cpuregs_reg_10__3_  (
    .CK(clk),
    .D(_01057_),
    .Q(\cpuregs[10] [3]),
    .QN(_28131_)
  );
  DFF_X1 cpuregs_reg_10__4_  (
    .CK(clk),
    .D(_01058_),
    .Q(\cpuregs[10] [4]),
    .QN(_28130_)
  );
  DFF_X1 cpuregs_reg_10__5_  (
    .CK(clk),
    .D(_01059_),
    .Q(\cpuregs[10] [5]),
    .QN(_28129_)
  );
  DFF_X1 cpuregs_reg_10__6_  (
    .CK(clk),
    .D(_01060_),
    .Q(\cpuregs[10] [6]),
    .QN(_28128_)
  );
  DFF_X1 cpuregs_reg_10__7_  (
    .CK(clk),
    .D(_01061_),
    .Q(\cpuregs[10] [7]),
    .QN(_28127_)
  );
  DFF_X1 cpuregs_reg_10__8_  (
    .CK(clk),
    .D(_01062_),
    .Q(\cpuregs[10] [8]),
    .QN(_28126_)
  );
  DFF_X1 cpuregs_reg_10__9_  (
    .CK(clk),
    .D(_01063_),
    .Q(\cpuregs[10] [9]),
    .QN(_28125_)
  );
  DFF_X1 cpuregs_reg_11__0_  (
    .CK(clk),
    .D(_00868_),
    .Q(\cpuregs[11] [0]),
    .QN(_28320_)
  );
  DFF_X1 cpuregs_reg_11__10_  (
    .CK(clk),
    .D(_00878_),
    .Q(\cpuregs[11] [10]),
    .QN(_28310_)
  );
  DFF_X1 cpuregs_reg_11__11_  (
    .CK(clk),
    .D(_00879_),
    .Q(\cpuregs[11] [11]),
    .QN(_28309_)
  );
  DFF_X1 cpuregs_reg_11__12_  (
    .CK(clk),
    .D(_00880_),
    .Q(\cpuregs[11] [12]),
    .QN(_28308_)
  );
  DFF_X1 cpuregs_reg_11__13_  (
    .CK(clk),
    .D(_00881_),
    .Q(\cpuregs[11] [13]),
    .QN(_28307_)
  );
  DFF_X1 cpuregs_reg_11__14_  (
    .CK(clk),
    .D(_00882_),
    .Q(\cpuregs[11] [14]),
    .QN(_28306_)
  );
  DFF_X1 cpuregs_reg_11__15_  (
    .CK(clk),
    .D(_00883_),
    .Q(\cpuregs[11] [15]),
    .QN(_28305_)
  );
  DFF_X1 cpuregs_reg_11__16_  (
    .CK(clk),
    .D(_00884_),
    .Q(\cpuregs[11] [16]),
    .QN(_28304_)
  );
  DFF_X1 cpuregs_reg_11__17_  (
    .CK(clk),
    .D(_00885_),
    .Q(\cpuregs[11] [17]),
    .QN(_28303_)
  );
  DFF_X1 cpuregs_reg_11__18_  (
    .CK(clk),
    .D(_00886_),
    .Q(\cpuregs[11] [18]),
    .QN(_28302_)
  );
  DFF_X1 cpuregs_reg_11__19_  (
    .CK(clk),
    .D(_00887_),
    .Q(\cpuregs[11] [19]),
    .QN(_28301_)
  );
  DFF_X1 cpuregs_reg_11__1_  (
    .CK(clk),
    .D(_00869_),
    .Q(\cpuregs[11] [1]),
    .QN(_28319_)
  );
  DFF_X1 cpuregs_reg_11__20_  (
    .CK(clk),
    .D(_00888_),
    .Q(\cpuregs[11] [20]),
    .QN(_28300_)
  );
  DFF_X1 cpuregs_reg_11__21_  (
    .CK(clk),
    .D(_00889_),
    .Q(\cpuregs[11] [21]),
    .QN(_28299_)
  );
  DFF_X1 cpuregs_reg_11__22_  (
    .CK(clk),
    .D(_00890_),
    .Q(\cpuregs[11] [22]),
    .QN(_28298_)
  );
  DFF_X1 cpuregs_reg_11__23_  (
    .CK(clk),
    .D(_00891_),
    .Q(\cpuregs[11] [23]),
    .QN(_28297_)
  );
  DFF_X1 cpuregs_reg_11__24_  (
    .CK(clk),
    .D(_00892_),
    .Q(\cpuregs[11] [24]),
    .QN(_28296_)
  );
  DFF_X1 cpuregs_reg_11__25_  (
    .CK(clk),
    .D(_00893_),
    .Q(\cpuregs[11] [25]),
    .QN(_28295_)
  );
  DFF_X1 cpuregs_reg_11__26_  (
    .CK(clk),
    .D(_00894_),
    .Q(\cpuregs[11] [26]),
    .QN(_28294_)
  );
  DFF_X1 cpuregs_reg_11__27_  (
    .CK(clk),
    .D(_00895_),
    .Q(\cpuregs[11] [27]),
    .QN(_28293_)
  );
  DFF_X1 cpuregs_reg_11__28_  (
    .CK(clk),
    .D(_00896_),
    .Q(\cpuregs[11] [28]),
    .QN(_28292_)
  );
  DFF_X1 cpuregs_reg_11__29_  (
    .CK(clk),
    .D(_00897_),
    .Q(\cpuregs[11] [29]),
    .QN(_28291_)
  );
  DFF_X1 cpuregs_reg_11__2_  (
    .CK(clk),
    .D(_00870_),
    .Q(\cpuregs[11] [2]),
    .QN(_28318_)
  );
  DFF_X1 cpuregs_reg_11__30_  (
    .CK(clk),
    .D(_00898_),
    .Q(\cpuregs[11] [30]),
    .QN(_28290_)
  );
  DFF_X1 cpuregs_reg_11__31_  (
    .CK(clk),
    .D(_00524_),
    .Q(\cpuregs[11] [31]),
    .QN(_28664_)
  );
  DFF_X1 cpuregs_reg_11__3_  (
    .CK(clk),
    .D(_00871_),
    .Q(\cpuregs[11] [3]),
    .QN(_28317_)
  );
  DFF_X1 cpuregs_reg_11__4_  (
    .CK(clk),
    .D(_00872_),
    .Q(\cpuregs[11] [4]),
    .QN(_28316_)
  );
  DFF_X1 cpuregs_reg_11__5_  (
    .CK(clk),
    .D(_00873_),
    .Q(\cpuregs[11] [5]),
    .QN(_28315_)
  );
  DFF_X1 cpuregs_reg_11__6_  (
    .CK(clk),
    .D(_00874_),
    .Q(\cpuregs[11] [6]),
    .QN(_28314_)
  );
  DFF_X1 cpuregs_reg_11__7_  (
    .CK(clk),
    .D(_00875_),
    .Q(\cpuregs[11] [7]),
    .QN(_28313_)
  );
  DFF_X1 cpuregs_reg_11__8_  (
    .CK(clk),
    .D(_00876_),
    .Q(\cpuregs[11] [8]),
    .QN(_28312_)
  );
  DFF_X1 cpuregs_reg_11__9_  (
    .CK(clk),
    .D(_00877_),
    .Q(\cpuregs[11] [9]),
    .QN(_28311_)
  );
  DFF_X1 cpuregs_reg_12__0_  (
    .CK(clk),
    .D(_00713_),
    .Q(\cpuregs[12] [0]),
    .QN(_28475_)
  );
  DFF_X1 cpuregs_reg_12__10_  (
    .CK(clk),
    .D(_00723_),
    .Q(\cpuregs[12] [10]),
    .QN(_28465_)
  );
  DFF_X1 cpuregs_reg_12__11_  (
    .CK(clk),
    .D(_00724_),
    .Q(\cpuregs[12] [11]),
    .QN(_28464_)
  );
  DFF_X1 cpuregs_reg_12__12_  (
    .CK(clk),
    .D(_00725_),
    .Q(\cpuregs[12] [12]),
    .QN(_28463_)
  );
  DFF_X1 cpuregs_reg_12__13_  (
    .CK(clk),
    .D(_00726_),
    .Q(\cpuregs[12] [13]),
    .QN(_28462_)
  );
  DFF_X1 cpuregs_reg_12__14_  (
    .CK(clk),
    .D(_00727_),
    .Q(\cpuregs[12] [14]),
    .QN(_28461_)
  );
  DFF_X1 cpuregs_reg_12__15_  (
    .CK(clk),
    .D(_00728_),
    .Q(\cpuregs[12] [15]),
    .QN(_28460_)
  );
  DFF_X1 cpuregs_reg_12__16_  (
    .CK(clk),
    .D(_00729_),
    .Q(\cpuregs[12] [16]),
    .QN(_28459_)
  );
  DFF_X1 cpuregs_reg_12__17_  (
    .CK(clk),
    .D(_00730_),
    .Q(\cpuregs[12] [17]),
    .QN(_28458_)
  );
  DFF_X1 cpuregs_reg_12__18_  (
    .CK(clk),
    .D(_00731_),
    .Q(\cpuregs[12] [18]),
    .QN(_28457_)
  );
  DFF_X1 cpuregs_reg_12__19_  (
    .CK(clk),
    .D(_00732_),
    .Q(\cpuregs[12] [19]),
    .QN(_28456_)
  );
  DFF_X1 cpuregs_reg_12__1_  (
    .CK(clk),
    .D(_00714_),
    .Q(\cpuregs[12] [1]),
    .QN(_28474_)
  );
  DFF_X1 cpuregs_reg_12__20_  (
    .CK(clk),
    .D(_00733_),
    .Q(\cpuregs[12] [20]),
    .QN(_28455_)
  );
  DFF_X1 cpuregs_reg_12__21_  (
    .CK(clk),
    .D(_00734_),
    .Q(\cpuregs[12] [21]),
    .QN(_28454_)
  );
  DFF_X1 cpuregs_reg_12__22_  (
    .CK(clk),
    .D(_00735_),
    .Q(\cpuregs[12] [22]),
    .QN(_28453_)
  );
  DFF_X1 cpuregs_reg_12__23_  (
    .CK(clk),
    .D(_00736_),
    .Q(\cpuregs[12] [23]),
    .QN(_28452_)
  );
  DFF_X1 cpuregs_reg_12__24_  (
    .CK(clk),
    .D(_00737_),
    .Q(\cpuregs[12] [24]),
    .QN(_28451_)
  );
  DFF_X1 cpuregs_reg_12__25_  (
    .CK(clk),
    .D(_00738_),
    .Q(\cpuregs[12] [25]),
    .QN(_28450_)
  );
  DFF_X1 cpuregs_reg_12__26_  (
    .CK(clk),
    .D(_00739_),
    .Q(\cpuregs[12] [26]),
    .QN(_28449_)
  );
  DFF_X1 cpuregs_reg_12__27_  (
    .CK(clk),
    .D(_00740_),
    .Q(\cpuregs[12] [27]),
    .QN(_28448_)
  );
  DFF_X1 cpuregs_reg_12__28_  (
    .CK(clk),
    .D(_00741_),
    .Q(\cpuregs[12] [28]),
    .QN(_28447_)
  );
  DFF_X1 cpuregs_reg_12__29_  (
    .CK(clk),
    .D(_00742_),
    .Q(\cpuregs[12] [29]),
    .QN(_28446_)
  );
  DFF_X1 cpuregs_reg_12__2_  (
    .CK(clk),
    .D(_00715_),
    .Q(\cpuregs[12] [2]),
    .QN(_28473_)
  );
  DFF_X1 cpuregs_reg_12__30_  (
    .CK(clk),
    .D(_00743_),
    .Q(\cpuregs[12] [30]),
    .QN(_28445_)
  );
  DFF_X1 cpuregs_reg_12__31_  (
    .CK(clk),
    .D(_00523_),
    .Q(\cpuregs[12] [31]),
    .QN(_28665_)
  );
  DFF_X1 cpuregs_reg_12__3_  (
    .CK(clk),
    .D(_00716_),
    .Q(\cpuregs[12] [3]),
    .QN(_28472_)
  );
  DFF_X1 cpuregs_reg_12__4_  (
    .CK(clk),
    .D(_00717_),
    .Q(\cpuregs[12] [4]),
    .QN(_28471_)
  );
  DFF_X1 cpuregs_reg_12__5_  (
    .CK(clk),
    .D(_00718_),
    .Q(\cpuregs[12] [5]),
    .QN(_28470_)
  );
  DFF_X1 cpuregs_reg_12__6_  (
    .CK(clk),
    .D(_00719_),
    .Q(\cpuregs[12] [6]),
    .QN(_28469_)
  );
  DFF_X1 cpuregs_reg_12__7_  (
    .CK(clk),
    .D(_00720_),
    .Q(\cpuregs[12] [7]),
    .QN(_28468_)
  );
  DFF_X1 cpuregs_reg_12__8_  (
    .CK(clk),
    .D(_00721_),
    .Q(\cpuregs[12] [8]),
    .QN(_28467_)
  );
  DFF_X1 cpuregs_reg_12__9_  (
    .CK(clk),
    .D(_00722_),
    .Q(\cpuregs[12] [9]),
    .QN(_28466_)
  );
  DFF_X1 cpuregs_reg_13__0_  (
    .CK(clk),
    .D(_00961_),
    .Q(\cpuregs[13] [0]),
    .QN(_28227_)
  );
  DFF_X1 cpuregs_reg_13__10_  (
    .CK(clk),
    .D(_00971_),
    .Q(\cpuregs[13] [10]),
    .QN(_28217_)
  );
  DFF_X1 cpuregs_reg_13__11_  (
    .CK(clk),
    .D(_00972_),
    .Q(\cpuregs[13] [11]),
    .QN(_28216_)
  );
  DFF_X1 cpuregs_reg_13__12_  (
    .CK(clk),
    .D(_00973_),
    .Q(\cpuregs[13] [12]),
    .QN(_28215_)
  );
  DFF_X1 cpuregs_reg_13__13_  (
    .CK(clk),
    .D(_00974_),
    .Q(\cpuregs[13] [13]),
    .QN(_28214_)
  );
  DFF_X1 cpuregs_reg_13__14_  (
    .CK(clk),
    .D(_00975_),
    .Q(\cpuregs[13] [14]),
    .QN(_28213_)
  );
  DFF_X1 cpuregs_reg_13__15_  (
    .CK(clk),
    .D(_00976_),
    .Q(\cpuregs[13] [15]),
    .QN(_28212_)
  );
  DFF_X1 cpuregs_reg_13__16_  (
    .CK(clk),
    .D(_00977_),
    .Q(\cpuregs[13] [16]),
    .QN(_28211_)
  );
  DFF_X1 cpuregs_reg_13__17_  (
    .CK(clk),
    .D(_00978_),
    .Q(\cpuregs[13] [17]),
    .QN(_28210_)
  );
  DFF_X1 cpuregs_reg_13__18_  (
    .CK(clk),
    .D(_00979_),
    .Q(\cpuregs[13] [18]),
    .QN(_28209_)
  );
  DFF_X1 cpuregs_reg_13__19_  (
    .CK(clk),
    .D(_00980_),
    .Q(\cpuregs[13] [19]),
    .QN(_28208_)
  );
  DFF_X1 cpuregs_reg_13__1_  (
    .CK(clk),
    .D(_00962_),
    .Q(\cpuregs[13] [1]),
    .QN(_28226_)
  );
  DFF_X1 cpuregs_reg_13__20_  (
    .CK(clk),
    .D(_00981_),
    .Q(\cpuregs[13] [20]),
    .QN(_28207_)
  );
  DFF_X1 cpuregs_reg_13__21_  (
    .CK(clk),
    .D(_00982_),
    .Q(\cpuregs[13] [21]),
    .QN(_28206_)
  );
  DFF_X1 cpuregs_reg_13__22_  (
    .CK(clk),
    .D(_00983_),
    .Q(\cpuregs[13] [22]),
    .QN(_28205_)
  );
  DFF_X1 cpuregs_reg_13__23_  (
    .CK(clk),
    .D(_00984_),
    .Q(\cpuregs[13] [23]),
    .QN(_28204_)
  );
  DFF_X1 cpuregs_reg_13__24_  (
    .CK(clk),
    .D(_00985_),
    .Q(\cpuregs[13] [24]),
    .QN(_28203_)
  );
  DFF_X1 cpuregs_reg_13__25_  (
    .CK(clk),
    .D(_00986_),
    .Q(\cpuregs[13] [25]),
    .QN(_28202_)
  );
  DFF_X1 cpuregs_reg_13__26_  (
    .CK(clk),
    .D(_00987_),
    .Q(\cpuregs[13] [26]),
    .QN(_28201_)
  );
  DFF_X1 cpuregs_reg_13__27_  (
    .CK(clk),
    .D(_00988_),
    .Q(\cpuregs[13] [27]),
    .QN(_28200_)
  );
  DFF_X1 cpuregs_reg_13__28_  (
    .CK(clk),
    .D(_00989_),
    .Q(\cpuregs[13] [28]),
    .QN(_28199_)
  );
  DFF_X1 cpuregs_reg_13__29_  (
    .CK(clk),
    .D(_00990_),
    .Q(\cpuregs[13] [29]),
    .QN(_28198_)
  );
  DFF_X1 cpuregs_reg_13__2_  (
    .CK(clk),
    .D(_00963_),
    .Q(\cpuregs[13] [2]),
    .QN(_28225_)
  );
  DFF_X1 cpuregs_reg_13__30_  (
    .CK(clk),
    .D(_00991_),
    .Q(\cpuregs[13] [30]),
    .QN(_28197_)
  );
  DFF_X1 cpuregs_reg_13__31_  (
    .CK(clk),
    .D(_00522_),
    .Q(\cpuregs[13] [31]),
    .QN(_28666_)
  );
  DFF_X1 cpuregs_reg_13__3_  (
    .CK(clk),
    .D(_00964_),
    .Q(\cpuregs[13] [3]),
    .QN(_28224_)
  );
  DFF_X1 cpuregs_reg_13__4_  (
    .CK(clk),
    .D(_00965_),
    .Q(\cpuregs[13] [4]),
    .QN(_28223_)
  );
  DFF_X1 cpuregs_reg_13__5_  (
    .CK(clk),
    .D(_00966_),
    .Q(\cpuregs[13] [5]),
    .QN(_28222_)
  );
  DFF_X1 cpuregs_reg_13__6_  (
    .CK(clk),
    .D(_00967_),
    .Q(\cpuregs[13] [6]),
    .QN(_28221_)
  );
  DFF_X1 cpuregs_reg_13__7_  (
    .CK(clk),
    .D(_00968_),
    .Q(\cpuregs[13] [7]),
    .QN(_28220_)
  );
  DFF_X1 cpuregs_reg_13__8_  (
    .CK(clk),
    .D(_00969_),
    .Q(\cpuregs[13] [8]),
    .QN(_28219_)
  );
  DFF_X1 cpuregs_reg_13__9_  (
    .CK(clk),
    .D(_00970_),
    .Q(\cpuregs[13] [9]),
    .QN(_28218_)
  );
  DFF_X1 cpuregs_reg_14__0_  (
    .CK(clk),
    .D(_00558_),
    .Q(\cpuregs[14] [0]),
    .QN(_28630_)
  );
  DFF_X1 cpuregs_reg_14__10_  (
    .CK(clk),
    .D(_00568_),
    .Q(\cpuregs[14] [10]),
    .QN(_28620_)
  );
  DFF_X1 cpuregs_reg_14__11_  (
    .CK(clk),
    .D(_00569_),
    .Q(\cpuregs[14] [11]),
    .QN(_28619_)
  );
  DFF_X1 cpuregs_reg_14__12_  (
    .CK(clk),
    .D(_00570_),
    .Q(\cpuregs[14] [12]),
    .QN(_28618_)
  );
  DFF_X1 cpuregs_reg_14__13_  (
    .CK(clk),
    .D(_00571_),
    .Q(\cpuregs[14] [13]),
    .QN(_28617_)
  );
  DFF_X1 cpuregs_reg_14__14_  (
    .CK(clk),
    .D(_00572_),
    .Q(\cpuregs[14] [14]),
    .QN(_28616_)
  );
  DFF_X1 cpuregs_reg_14__15_  (
    .CK(clk),
    .D(_00573_),
    .Q(\cpuregs[14] [15]),
    .QN(_28615_)
  );
  DFF_X1 cpuregs_reg_14__16_  (
    .CK(clk),
    .D(_00574_),
    .Q(\cpuregs[14] [16]),
    .QN(_28614_)
  );
  DFF_X1 cpuregs_reg_14__17_  (
    .CK(clk),
    .D(_00575_),
    .Q(\cpuregs[14] [17]),
    .QN(_28613_)
  );
  DFF_X1 cpuregs_reg_14__18_  (
    .CK(clk),
    .D(_00576_),
    .Q(\cpuregs[14] [18]),
    .QN(_28612_)
  );
  DFF_X1 cpuregs_reg_14__19_  (
    .CK(clk),
    .D(_00577_),
    .Q(\cpuregs[14] [19]),
    .QN(_28611_)
  );
  DFF_X1 cpuregs_reg_14__1_  (
    .CK(clk),
    .D(_00559_),
    .Q(\cpuregs[14] [1]),
    .QN(_28629_)
  );
  DFF_X1 cpuregs_reg_14__20_  (
    .CK(clk),
    .D(_00578_),
    .Q(\cpuregs[14] [20]),
    .QN(_28610_)
  );
  DFF_X1 cpuregs_reg_14__21_  (
    .CK(clk),
    .D(_00579_),
    .Q(\cpuregs[14] [21]),
    .QN(_28609_)
  );
  DFF_X1 cpuregs_reg_14__22_  (
    .CK(clk),
    .D(_00580_),
    .Q(\cpuregs[14] [22]),
    .QN(_28608_)
  );
  DFF_X1 cpuregs_reg_14__23_  (
    .CK(clk),
    .D(_00581_),
    .Q(\cpuregs[14] [23]),
    .QN(_28607_)
  );
  DFF_X1 cpuregs_reg_14__24_  (
    .CK(clk),
    .D(_00582_),
    .Q(\cpuregs[14] [24]),
    .QN(_28606_)
  );
  DFF_X1 cpuregs_reg_14__25_  (
    .CK(clk),
    .D(_00583_),
    .Q(\cpuregs[14] [25]),
    .QN(_28605_)
  );
  DFF_X1 cpuregs_reg_14__26_  (
    .CK(clk),
    .D(_00584_),
    .Q(\cpuregs[14] [26]),
    .QN(_28604_)
  );
  DFF_X1 cpuregs_reg_14__27_  (
    .CK(clk),
    .D(_00585_),
    .Q(\cpuregs[14] [27]),
    .QN(_28603_)
  );
  DFF_X1 cpuregs_reg_14__28_  (
    .CK(clk),
    .D(_00586_),
    .Q(\cpuregs[14] [28]),
    .QN(_28602_)
  );
  DFF_X1 cpuregs_reg_14__29_  (
    .CK(clk),
    .D(_00587_),
    .Q(\cpuregs[14] [29]),
    .QN(_28601_)
  );
  DFF_X1 cpuregs_reg_14__2_  (
    .CK(clk),
    .D(_00560_),
    .Q(\cpuregs[14] [2]),
    .QN(_28628_)
  );
  DFF_X1 cpuregs_reg_14__30_  (
    .CK(clk),
    .D(_00588_),
    .Q(\cpuregs[14] [30]),
    .QN(_28600_)
  );
  DFF_X1 cpuregs_reg_14__31_  (
    .CK(clk),
    .D(_00521_),
    .Q(\cpuregs[14] [31]),
    .QN(_28667_)
  );
  DFF_X1 cpuregs_reg_14__3_  (
    .CK(clk),
    .D(_00561_),
    .Q(\cpuregs[14] [3]),
    .QN(_28627_)
  );
  DFF_X1 cpuregs_reg_14__4_  (
    .CK(clk),
    .D(_00562_),
    .Q(\cpuregs[14] [4]),
    .QN(_28626_)
  );
  DFF_X1 cpuregs_reg_14__5_  (
    .CK(clk),
    .D(_00563_),
    .Q(\cpuregs[14] [5]),
    .QN(_28625_)
  );
  DFF_X1 cpuregs_reg_14__6_  (
    .CK(clk),
    .D(_00564_),
    .Q(\cpuregs[14] [6]),
    .QN(_28624_)
  );
  DFF_X1 cpuregs_reg_14__7_  (
    .CK(clk),
    .D(_00565_),
    .Q(\cpuregs[14] [7]),
    .QN(_28623_)
  );
  DFF_X1 cpuregs_reg_14__8_  (
    .CK(clk),
    .D(_00566_),
    .Q(\cpuregs[14] [8]),
    .QN(_28622_)
  );
  DFF_X1 cpuregs_reg_14__9_  (
    .CK(clk),
    .D(_00567_),
    .Q(\cpuregs[14] [9]),
    .QN(_28621_)
  );
  DFF_X1 cpuregs_reg_15__0_  (
    .CK(clk),
    .D(_00589_),
    .Q(\cpuregs[15] [0]),
    .QN(_28599_)
  );
  DFF_X1 cpuregs_reg_15__10_  (
    .CK(clk),
    .D(_00599_),
    .Q(\cpuregs[15] [10]),
    .QN(_28589_)
  );
  DFF_X1 cpuregs_reg_15__11_  (
    .CK(clk),
    .D(_00600_),
    .Q(\cpuregs[15] [11]),
    .QN(_28588_)
  );
  DFF_X1 cpuregs_reg_15__12_  (
    .CK(clk),
    .D(_00601_),
    .Q(\cpuregs[15] [12]),
    .QN(_28587_)
  );
  DFF_X1 cpuregs_reg_15__13_  (
    .CK(clk),
    .D(_00602_),
    .Q(\cpuregs[15] [13]),
    .QN(_28586_)
  );
  DFF_X1 cpuregs_reg_15__14_  (
    .CK(clk),
    .D(_00603_),
    .Q(\cpuregs[15] [14]),
    .QN(_28585_)
  );
  DFF_X1 cpuregs_reg_15__15_  (
    .CK(clk),
    .D(_00604_),
    .Q(\cpuregs[15] [15]),
    .QN(_28584_)
  );
  DFF_X1 cpuregs_reg_15__16_  (
    .CK(clk),
    .D(_00605_),
    .Q(\cpuregs[15] [16]),
    .QN(_28583_)
  );
  DFF_X1 cpuregs_reg_15__17_  (
    .CK(clk),
    .D(_00606_),
    .Q(\cpuregs[15] [17]),
    .QN(_28582_)
  );
  DFF_X1 cpuregs_reg_15__18_  (
    .CK(clk),
    .D(_00607_),
    .Q(\cpuregs[15] [18]),
    .QN(_28581_)
  );
  DFF_X1 cpuregs_reg_15__19_  (
    .CK(clk),
    .D(_00608_),
    .Q(\cpuregs[15] [19]),
    .QN(_28580_)
  );
  DFF_X1 cpuregs_reg_15__1_  (
    .CK(clk),
    .D(_00590_),
    .Q(\cpuregs[15] [1]),
    .QN(_28598_)
  );
  DFF_X1 cpuregs_reg_15__20_  (
    .CK(clk),
    .D(_00609_),
    .Q(\cpuregs[15] [20]),
    .QN(_28579_)
  );
  DFF_X1 cpuregs_reg_15__21_  (
    .CK(clk),
    .D(_00610_),
    .Q(\cpuregs[15] [21]),
    .QN(_28578_)
  );
  DFF_X1 cpuregs_reg_15__22_  (
    .CK(clk),
    .D(_00611_),
    .Q(\cpuregs[15] [22]),
    .QN(_28577_)
  );
  DFF_X1 cpuregs_reg_15__23_  (
    .CK(clk),
    .D(_00612_),
    .Q(\cpuregs[15] [23]),
    .QN(_28576_)
  );
  DFF_X1 cpuregs_reg_15__24_  (
    .CK(clk),
    .D(_00613_),
    .Q(\cpuregs[15] [24]),
    .QN(_28575_)
  );
  DFF_X1 cpuregs_reg_15__25_  (
    .CK(clk),
    .D(_00614_),
    .Q(\cpuregs[15] [25]),
    .QN(_28574_)
  );
  DFF_X1 cpuregs_reg_15__26_  (
    .CK(clk),
    .D(_00615_),
    .Q(\cpuregs[15] [26]),
    .QN(_28573_)
  );
  DFF_X1 cpuregs_reg_15__27_  (
    .CK(clk),
    .D(_00616_),
    .Q(\cpuregs[15] [27]),
    .QN(_28572_)
  );
  DFF_X1 cpuregs_reg_15__28_  (
    .CK(clk),
    .D(_00617_),
    .Q(\cpuregs[15] [28]),
    .QN(_28571_)
  );
  DFF_X1 cpuregs_reg_15__29_  (
    .CK(clk),
    .D(_00618_),
    .Q(\cpuregs[15] [29]),
    .QN(_28570_)
  );
  DFF_X1 cpuregs_reg_15__2_  (
    .CK(clk),
    .D(_00591_),
    .Q(\cpuregs[15] [2]),
    .QN(_28597_)
  );
  DFF_X1 cpuregs_reg_15__30_  (
    .CK(clk),
    .D(_00619_),
    .Q(\cpuregs[15] [30]),
    .QN(_28569_)
  );
  DFF_X1 cpuregs_reg_15__31_  (
    .CK(clk),
    .D(_00520_),
    .Q(\cpuregs[15] [31]),
    .QN(_28668_)
  );
  DFF_X1 cpuregs_reg_15__3_  (
    .CK(clk),
    .D(_00592_),
    .Q(\cpuregs[15] [3]),
    .QN(_28596_)
  );
  DFF_X1 cpuregs_reg_15__4_  (
    .CK(clk),
    .D(_00593_),
    .Q(\cpuregs[15] [4]),
    .QN(_28595_)
  );
  DFF_X1 cpuregs_reg_15__5_  (
    .CK(clk),
    .D(_00594_),
    .Q(\cpuregs[15] [5]),
    .QN(_28594_)
  );
  DFF_X1 cpuregs_reg_15__6_  (
    .CK(clk),
    .D(_00595_),
    .Q(\cpuregs[15] [6]),
    .QN(_28593_)
  );
  DFF_X1 cpuregs_reg_15__7_  (
    .CK(clk),
    .D(_00596_),
    .Q(\cpuregs[15] [7]),
    .QN(_28592_)
  );
  DFF_X1 cpuregs_reg_15__8_  (
    .CK(clk),
    .D(_00597_),
    .Q(\cpuregs[15] [8]),
    .QN(_28591_)
  );
  DFF_X1 cpuregs_reg_15__9_  (
    .CK(clk),
    .D(_00598_),
    .Q(\cpuregs[15] [9]),
    .QN(_28590_)
  );
  DFF_X1 cpuregs_reg_16__0_  (
    .CK(clk),
    .D(_00651_),
    .Q(\cpuregs[16] [0]),
    .QN(_28537_)
  );
  DFF_X1 cpuregs_reg_16__10_  (
    .CK(clk),
    .D(_00661_),
    .Q(\cpuregs[16] [10]),
    .QN(_28527_)
  );
  DFF_X1 cpuregs_reg_16__11_  (
    .CK(clk),
    .D(_00662_),
    .Q(\cpuregs[16] [11]),
    .QN(_28526_)
  );
  DFF_X1 cpuregs_reg_16__12_  (
    .CK(clk),
    .D(_00663_),
    .Q(\cpuregs[16] [12]),
    .QN(_28525_)
  );
  DFF_X1 cpuregs_reg_16__13_  (
    .CK(clk),
    .D(_00664_),
    .Q(\cpuregs[16] [13]),
    .QN(_28524_)
  );
  DFF_X1 cpuregs_reg_16__14_  (
    .CK(clk),
    .D(_00665_),
    .Q(\cpuregs[16] [14]),
    .QN(_28523_)
  );
  DFF_X1 cpuregs_reg_16__15_  (
    .CK(clk),
    .D(_00666_),
    .Q(\cpuregs[16] [15]),
    .QN(_28522_)
  );
  DFF_X1 cpuregs_reg_16__16_  (
    .CK(clk),
    .D(_00667_),
    .Q(\cpuregs[16] [16]),
    .QN(_28521_)
  );
  DFF_X1 cpuregs_reg_16__17_  (
    .CK(clk),
    .D(_00668_),
    .Q(\cpuregs[16] [17]),
    .QN(_28520_)
  );
  DFF_X1 cpuregs_reg_16__18_  (
    .CK(clk),
    .D(_00669_),
    .Q(\cpuregs[16] [18]),
    .QN(_28519_)
  );
  DFF_X1 cpuregs_reg_16__19_  (
    .CK(clk),
    .D(_00670_),
    .Q(\cpuregs[16] [19]),
    .QN(_28518_)
  );
  DFF_X1 cpuregs_reg_16__1_  (
    .CK(clk),
    .D(_00652_),
    .Q(\cpuregs[16] [1]),
    .QN(_28536_)
  );
  DFF_X1 cpuregs_reg_16__20_  (
    .CK(clk),
    .D(_00671_),
    .Q(\cpuregs[16] [20]),
    .QN(_28517_)
  );
  DFF_X1 cpuregs_reg_16__21_  (
    .CK(clk),
    .D(_00672_),
    .Q(\cpuregs[16] [21]),
    .QN(_28516_)
  );
  DFF_X1 cpuregs_reg_16__22_  (
    .CK(clk),
    .D(_00673_),
    .Q(\cpuregs[16] [22]),
    .QN(_28515_)
  );
  DFF_X1 cpuregs_reg_16__23_  (
    .CK(clk),
    .D(_00674_),
    .Q(\cpuregs[16] [23]),
    .QN(_28514_)
  );
  DFF_X1 cpuregs_reg_16__24_  (
    .CK(clk),
    .D(_00675_),
    .Q(\cpuregs[16] [24]),
    .QN(_28513_)
  );
  DFF_X1 cpuregs_reg_16__25_  (
    .CK(clk),
    .D(_00676_),
    .Q(\cpuregs[16] [25]),
    .QN(_28512_)
  );
  DFF_X1 cpuregs_reg_16__26_  (
    .CK(clk),
    .D(_00677_),
    .Q(\cpuregs[16] [26]),
    .QN(_28511_)
  );
  DFF_X1 cpuregs_reg_16__27_  (
    .CK(clk),
    .D(_00678_),
    .Q(\cpuregs[16] [27]),
    .QN(_28510_)
  );
  DFF_X1 cpuregs_reg_16__28_  (
    .CK(clk),
    .D(_00679_),
    .Q(\cpuregs[16] [28]),
    .QN(_28509_)
  );
  DFF_X1 cpuregs_reg_16__29_  (
    .CK(clk),
    .D(_00680_),
    .Q(\cpuregs[16] [29]),
    .QN(_28508_)
  );
  DFF_X1 cpuregs_reg_16__2_  (
    .CK(clk),
    .D(_00653_),
    .Q(\cpuregs[16] [2]),
    .QN(_28535_)
  );
  DFF_X1 cpuregs_reg_16__30_  (
    .CK(clk),
    .D(_00681_),
    .Q(\cpuregs[16] [30]),
    .QN(_28507_)
  );
  DFF_X1 cpuregs_reg_16__31_  (
    .CK(clk),
    .D(_00519_),
    .Q(\cpuregs[16] [31]),
    .QN(_28669_)
  );
  DFF_X1 cpuregs_reg_16__3_  (
    .CK(clk),
    .D(_00654_),
    .Q(\cpuregs[16] [3]),
    .QN(_28534_)
  );
  DFF_X1 cpuregs_reg_16__4_  (
    .CK(clk),
    .D(_00655_),
    .Q(\cpuregs[16] [4]),
    .QN(_28533_)
  );
  DFF_X1 cpuregs_reg_16__5_  (
    .CK(clk),
    .D(_00656_),
    .Q(\cpuregs[16] [5]),
    .QN(_28532_)
  );
  DFF_X1 cpuregs_reg_16__6_  (
    .CK(clk),
    .D(_00657_),
    .Q(\cpuregs[16] [6]),
    .QN(_28531_)
  );
  DFF_X1 cpuregs_reg_16__7_  (
    .CK(clk),
    .D(_00658_),
    .Q(\cpuregs[16] [7]),
    .QN(_28530_)
  );
  DFF_X1 cpuregs_reg_16__8_  (
    .CK(clk),
    .D(_00659_),
    .Q(\cpuregs[16] [8]),
    .QN(_28529_)
  );
  DFF_X1 cpuregs_reg_16__9_  (
    .CK(clk),
    .D(_00660_),
    .Q(\cpuregs[16] [9]),
    .QN(_28528_)
  );
  DFF_X1 cpuregs_reg_17__0_  (
    .CK(clk),
    .D(_00682_),
    .Q(\cpuregs[17] [0]),
    .QN(_28506_)
  );
  DFF_X1 cpuregs_reg_17__10_  (
    .CK(clk),
    .D(_00692_),
    .Q(\cpuregs[17] [10]),
    .QN(_28496_)
  );
  DFF_X1 cpuregs_reg_17__11_  (
    .CK(clk),
    .D(_00693_),
    .Q(\cpuregs[17] [11]),
    .QN(_28495_)
  );
  DFF_X1 cpuregs_reg_17__12_  (
    .CK(clk),
    .D(_00694_),
    .Q(\cpuregs[17] [12]),
    .QN(_28494_)
  );
  DFF_X1 cpuregs_reg_17__13_  (
    .CK(clk),
    .D(_00695_),
    .Q(\cpuregs[17] [13]),
    .QN(_28493_)
  );
  DFF_X1 cpuregs_reg_17__14_  (
    .CK(clk),
    .D(_00696_),
    .Q(\cpuregs[17] [14]),
    .QN(_28492_)
  );
  DFF_X1 cpuregs_reg_17__15_  (
    .CK(clk),
    .D(_00697_),
    .Q(\cpuregs[17] [15]),
    .QN(_28491_)
  );
  DFF_X1 cpuregs_reg_17__16_  (
    .CK(clk),
    .D(_00698_),
    .Q(\cpuregs[17] [16]),
    .QN(_28490_)
  );
  DFF_X1 cpuregs_reg_17__17_  (
    .CK(clk),
    .D(_00699_),
    .Q(\cpuregs[17] [17]),
    .QN(_28489_)
  );
  DFF_X1 cpuregs_reg_17__18_  (
    .CK(clk),
    .D(_00700_),
    .Q(\cpuregs[17] [18]),
    .QN(_28488_)
  );
  DFF_X1 cpuregs_reg_17__19_  (
    .CK(clk),
    .D(_00701_),
    .Q(\cpuregs[17] [19]),
    .QN(_28487_)
  );
  DFF_X1 cpuregs_reg_17__1_  (
    .CK(clk),
    .D(_00683_),
    .Q(\cpuregs[17] [1]),
    .QN(_28505_)
  );
  DFF_X1 cpuregs_reg_17__20_  (
    .CK(clk),
    .D(_00702_),
    .Q(\cpuregs[17] [20]),
    .QN(_28486_)
  );
  DFF_X1 cpuregs_reg_17__21_  (
    .CK(clk),
    .D(_00703_),
    .Q(\cpuregs[17] [21]),
    .QN(_28485_)
  );
  DFF_X1 cpuregs_reg_17__22_  (
    .CK(clk),
    .D(_00704_),
    .Q(\cpuregs[17] [22]),
    .QN(_28484_)
  );
  DFF_X1 cpuregs_reg_17__23_  (
    .CK(clk),
    .D(_00705_),
    .Q(\cpuregs[17] [23]),
    .QN(_28483_)
  );
  DFF_X1 cpuregs_reg_17__24_  (
    .CK(clk),
    .D(_00706_),
    .Q(\cpuregs[17] [24]),
    .QN(_28482_)
  );
  DFF_X1 cpuregs_reg_17__25_  (
    .CK(clk),
    .D(_00707_),
    .Q(\cpuregs[17] [25]),
    .QN(_28481_)
  );
  DFF_X1 cpuregs_reg_17__26_  (
    .CK(clk),
    .D(_00708_),
    .Q(\cpuregs[17] [26]),
    .QN(_28480_)
  );
  DFF_X1 cpuregs_reg_17__27_  (
    .CK(clk),
    .D(_00709_),
    .Q(\cpuregs[17] [27]),
    .QN(_28479_)
  );
  DFF_X1 cpuregs_reg_17__28_  (
    .CK(clk),
    .D(_00710_),
    .Q(\cpuregs[17] [28]),
    .QN(_28478_)
  );
  DFF_X1 cpuregs_reg_17__29_  (
    .CK(clk),
    .D(_00711_),
    .Q(\cpuregs[17] [29]),
    .QN(_28477_)
  );
  DFF_X1 cpuregs_reg_17__2_  (
    .CK(clk),
    .D(_00684_),
    .Q(\cpuregs[17] [2]),
    .QN(_28504_)
  );
  DFF_X1 cpuregs_reg_17__30_  (
    .CK(clk),
    .D(_00712_),
    .Q(\cpuregs[17] [30]),
    .QN(_28476_)
  );
  DFF_X1 cpuregs_reg_17__31_  (
    .CK(clk),
    .D(_00518_),
    .Q(\cpuregs[17] [31]),
    .QN(_28670_)
  );
  DFF_X1 cpuregs_reg_17__3_  (
    .CK(clk),
    .D(_00685_),
    .Q(\cpuregs[17] [3]),
    .QN(_28503_)
  );
  DFF_X1 cpuregs_reg_17__4_  (
    .CK(clk),
    .D(_00686_),
    .Q(\cpuregs[17] [4]),
    .QN(_28502_)
  );
  DFF_X1 cpuregs_reg_17__5_  (
    .CK(clk),
    .D(_00687_),
    .Q(\cpuregs[17] [5]),
    .QN(_28501_)
  );
  DFF_X1 cpuregs_reg_17__6_  (
    .CK(clk),
    .D(_00688_),
    .Q(\cpuregs[17] [6]),
    .QN(_28500_)
  );
  DFF_X1 cpuregs_reg_17__7_  (
    .CK(clk),
    .D(_00689_),
    .Q(\cpuregs[17] [7]),
    .QN(_28499_)
  );
  DFF_X1 cpuregs_reg_17__8_  (
    .CK(clk),
    .D(_00690_),
    .Q(\cpuregs[17] [8]),
    .QN(_28498_)
  );
  DFF_X1 cpuregs_reg_17__9_  (
    .CK(clk),
    .D(_00691_),
    .Q(\cpuregs[17] [9]),
    .QN(_28497_)
  );
  DFF_X1 cpuregs_reg_18__0_  (
    .CK(clk),
    .D(_00899_),
    .Q(\cpuregs[18] [0]),
    .QN(_28289_)
  );
  DFF_X1 cpuregs_reg_18__10_  (
    .CK(clk),
    .D(_00909_),
    .Q(\cpuregs[18] [10]),
    .QN(_28279_)
  );
  DFF_X1 cpuregs_reg_18__11_  (
    .CK(clk),
    .D(_00910_),
    .Q(\cpuregs[18] [11]),
    .QN(_28278_)
  );
  DFF_X1 cpuregs_reg_18__12_  (
    .CK(clk),
    .D(_00911_),
    .Q(\cpuregs[18] [12]),
    .QN(_28277_)
  );
  DFF_X1 cpuregs_reg_18__13_  (
    .CK(clk),
    .D(_00912_),
    .Q(\cpuregs[18] [13]),
    .QN(_28276_)
  );
  DFF_X1 cpuregs_reg_18__14_  (
    .CK(clk),
    .D(_00913_),
    .Q(\cpuregs[18] [14]),
    .QN(_28275_)
  );
  DFF_X1 cpuregs_reg_18__15_  (
    .CK(clk),
    .D(_00914_),
    .Q(\cpuregs[18] [15]),
    .QN(_28274_)
  );
  DFF_X1 cpuregs_reg_18__16_  (
    .CK(clk),
    .D(_00915_),
    .Q(\cpuregs[18] [16]),
    .QN(_28273_)
  );
  DFF_X1 cpuregs_reg_18__17_  (
    .CK(clk),
    .D(_00916_),
    .Q(\cpuregs[18] [17]),
    .QN(_28272_)
  );
  DFF_X1 cpuregs_reg_18__18_  (
    .CK(clk),
    .D(_00917_),
    .Q(\cpuregs[18] [18]),
    .QN(_28271_)
  );
  DFF_X1 cpuregs_reg_18__19_  (
    .CK(clk),
    .D(_00918_),
    .Q(\cpuregs[18] [19]),
    .QN(_28270_)
  );
  DFF_X1 cpuregs_reg_18__1_  (
    .CK(clk),
    .D(_00900_),
    .Q(\cpuregs[18] [1]),
    .QN(_28288_)
  );
  DFF_X1 cpuregs_reg_18__20_  (
    .CK(clk),
    .D(_00919_),
    .Q(\cpuregs[18] [20]),
    .QN(_28269_)
  );
  DFF_X1 cpuregs_reg_18__21_  (
    .CK(clk),
    .D(_00920_),
    .Q(\cpuregs[18] [21]),
    .QN(_28268_)
  );
  DFF_X1 cpuregs_reg_18__22_  (
    .CK(clk),
    .D(_00921_),
    .Q(\cpuregs[18] [22]),
    .QN(_28267_)
  );
  DFF_X1 cpuregs_reg_18__23_  (
    .CK(clk),
    .D(_00922_),
    .Q(\cpuregs[18] [23]),
    .QN(_28266_)
  );
  DFF_X1 cpuregs_reg_18__24_  (
    .CK(clk),
    .D(_00923_),
    .Q(\cpuregs[18] [24]),
    .QN(_28265_)
  );
  DFF_X1 cpuregs_reg_18__25_  (
    .CK(clk),
    .D(_00924_),
    .Q(\cpuregs[18] [25]),
    .QN(_28264_)
  );
  DFF_X1 cpuregs_reg_18__26_  (
    .CK(clk),
    .D(_00925_),
    .Q(\cpuregs[18] [26]),
    .QN(_28263_)
  );
  DFF_X1 cpuregs_reg_18__27_  (
    .CK(clk),
    .D(_00926_),
    .Q(\cpuregs[18] [27]),
    .QN(_28262_)
  );
  DFF_X1 cpuregs_reg_18__28_  (
    .CK(clk),
    .D(_00927_),
    .Q(\cpuregs[18] [28]),
    .QN(_28261_)
  );
  DFF_X1 cpuregs_reg_18__29_  (
    .CK(clk),
    .D(_00928_),
    .Q(\cpuregs[18] [29]),
    .QN(_28260_)
  );
  DFF_X1 cpuregs_reg_18__2_  (
    .CK(clk),
    .D(_00901_),
    .Q(\cpuregs[18] [2]),
    .QN(_28287_)
  );
  DFF_X1 cpuregs_reg_18__30_  (
    .CK(clk),
    .D(_00929_),
    .Q(\cpuregs[18] [30]),
    .QN(_28259_)
  );
  DFF_X1 cpuregs_reg_18__31_  (
    .CK(clk),
    .D(_00517_),
    .Q(\cpuregs[18] [31]),
    .QN(_28671_)
  );
  DFF_X1 cpuregs_reg_18__3_  (
    .CK(clk),
    .D(_00902_),
    .Q(\cpuregs[18] [3]),
    .QN(_28286_)
  );
  DFF_X1 cpuregs_reg_18__4_  (
    .CK(clk),
    .D(_00903_),
    .Q(\cpuregs[18] [4]),
    .QN(_28285_)
  );
  DFF_X1 cpuregs_reg_18__5_  (
    .CK(clk),
    .D(_00904_),
    .Q(\cpuregs[18] [5]),
    .QN(_28284_)
  );
  DFF_X1 cpuregs_reg_18__6_  (
    .CK(clk),
    .D(_00905_),
    .Q(\cpuregs[18] [6]),
    .QN(_28283_)
  );
  DFF_X1 cpuregs_reg_18__7_  (
    .CK(clk),
    .D(_00906_),
    .Q(\cpuregs[18] [7]),
    .QN(_28282_)
  );
  DFF_X1 cpuregs_reg_18__8_  (
    .CK(clk),
    .D(_00907_),
    .Q(\cpuregs[18] [8]),
    .QN(_28281_)
  );
  DFF_X1 cpuregs_reg_18__9_  (
    .CK(clk),
    .D(_00908_),
    .Q(\cpuregs[18] [9]),
    .QN(_28280_)
  );
  DFF_X1 cpuregs_reg_19__0_  (
    .CK(clk),
    .D(_00930_),
    .Q(\cpuregs[19] [0]),
    .QN(_28258_)
  );
  DFF_X1 cpuregs_reg_19__10_  (
    .CK(clk),
    .D(_00940_),
    .Q(\cpuregs[19] [10]),
    .QN(_28248_)
  );
  DFF_X1 cpuregs_reg_19__11_  (
    .CK(clk),
    .D(_00941_),
    .Q(\cpuregs[19] [11]),
    .QN(_28247_)
  );
  DFF_X1 cpuregs_reg_19__12_  (
    .CK(clk),
    .D(_00942_),
    .Q(\cpuregs[19] [12]),
    .QN(_28246_)
  );
  DFF_X1 cpuregs_reg_19__13_  (
    .CK(clk),
    .D(_00943_),
    .Q(\cpuregs[19] [13]),
    .QN(_28245_)
  );
  DFF_X1 cpuregs_reg_19__14_  (
    .CK(clk),
    .D(_00944_),
    .Q(\cpuregs[19] [14]),
    .QN(_28244_)
  );
  DFF_X1 cpuregs_reg_19__15_  (
    .CK(clk),
    .D(_00945_),
    .Q(\cpuregs[19] [15]),
    .QN(_28243_)
  );
  DFF_X1 cpuregs_reg_19__16_  (
    .CK(clk),
    .D(_00946_),
    .Q(\cpuregs[19] [16]),
    .QN(_28242_)
  );
  DFF_X1 cpuregs_reg_19__17_  (
    .CK(clk),
    .D(_00947_),
    .Q(\cpuregs[19] [17]),
    .QN(_28241_)
  );
  DFF_X1 cpuregs_reg_19__18_  (
    .CK(clk),
    .D(_00948_),
    .Q(\cpuregs[19] [18]),
    .QN(_28240_)
  );
  DFF_X1 cpuregs_reg_19__19_  (
    .CK(clk),
    .D(_00949_),
    .Q(\cpuregs[19] [19]),
    .QN(_28239_)
  );
  DFF_X1 cpuregs_reg_19__1_  (
    .CK(clk),
    .D(_00931_),
    .Q(\cpuregs[19] [1]),
    .QN(_28257_)
  );
  DFF_X1 cpuregs_reg_19__20_  (
    .CK(clk),
    .D(_00950_),
    .Q(\cpuregs[19] [20]),
    .QN(_28238_)
  );
  DFF_X1 cpuregs_reg_19__21_  (
    .CK(clk),
    .D(_00951_),
    .Q(\cpuregs[19] [21]),
    .QN(_28237_)
  );
  DFF_X1 cpuregs_reg_19__22_  (
    .CK(clk),
    .D(_00952_),
    .Q(\cpuregs[19] [22]),
    .QN(_28236_)
  );
  DFF_X1 cpuregs_reg_19__23_  (
    .CK(clk),
    .D(_00953_),
    .Q(\cpuregs[19] [23]),
    .QN(_28235_)
  );
  DFF_X1 cpuregs_reg_19__24_  (
    .CK(clk),
    .D(_00954_),
    .Q(\cpuregs[19] [24]),
    .QN(_28234_)
  );
  DFF_X1 cpuregs_reg_19__25_  (
    .CK(clk),
    .D(_00955_),
    .Q(\cpuregs[19] [25]),
    .QN(_28233_)
  );
  DFF_X1 cpuregs_reg_19__26_  (
    .CK(clk),
    .D(_00956_),
    .Q(\cpuregs[19] [26]),
    .QN(_28232_)
  );
  DFF_X1 cpuregs_reg_19__27_  (
    .CK(clk),
    .D(_00957_),
    .Q(\cpuregs[19] [27]),
    .QN(_28231_)
  );
  DFF_X1 cpuregs_reg_19__28_  (
    .CK(clk),
    .D(_00958_),
    .Q(\cpuregs[19] [28]),
    .QN(_28230_)
  );
  DFF_X1 cpuregs_reg_19__29_  (
    .CK(clk),
    .D(_00959_),
    .Q(\cpuregs[19] [29]),
    .QN(_28229_)
  );
  DFF_X1 cpuregs_reg_19__2_  (
    .CK(clk),
    .D(_00932_),
    .Q(\cpuregs[19] [2]),
    .QN(_28256_)
  );
  DFF_X1 cpuregs_reg_19__30_  (
    .CK(clk),
    .D(_00960_),
    .Q(\cpuregs[19] [30]),
    .QN(_28228_)
  );
  DFF_X1 cpuregs_reg_19__31_  (
    .CK(clk),
    .D(_00516_),
    .Q(\cpuregs[19] [31]),
    .QN(_28672_)
  );
  DFF_X1 cpuregs_reg_19__3_  (
    .CK(clk),
    .D(_00933_),
    .Q(\cpuregs[19] [3]),
    .QN(_28255_)
  );
  DFF_X1 cpuregs_reg_19__4_  (
    .CK(clk),
    .D(_00934_),
    .Q(\cpuregs[19] [4]),
    .QN(_28254_)
  );
  DFF_X1 cpuregs_reg_19__5_  (
    .CK(clk),
    .D(_00935_),
    .Q(\cpuregs[19] [5]),
    .QN(_28253_)
  );
  DFF_X1 cpuregs_reg_19__6_  (
    .CK(clk),
    .D(_00936_),
    .Q(\cpuregs[19] [6]),
    .QN(_28252_)
  );
  DFF_X1 cpuregs_reg_19__7_  (
    .CK(clk),
    .D(_00937_),
    .Q(\cpuregs[19] [7]),
    .QN(_28251_)
  );
  DFF_X1 cpuregs_reg_19__8_  (
    .CK(clk),
    .D(_00938_),
    .Q(\cpuregs[19] [8]),
    .QN(_28250_)
  );
  DFF_X1 cpuregs_reg_19__9_  (
    .CK(clk),
    .D(_00939_),
    .Q(\cpuregs[19] [9]),
    .QN(_28249_)
  );
  DFF_X1 cpuregs_reg_1__0_  (
    .CK(clk),
    .D(_00775_),
    .Q(\cpuregs[1] [0]),
    .QN(_28413_)
  );
  DFF_X1 cpuregs_reg_1__10_  (
    .CK(clk),
    .D(_00785_),
    .Q(\cpuregs[1] [10]),
    .QN(_28403_)
  );
  DFF_X1 cpuregs_reg_1__11_  (
    .CK(clk),
    .D(_00786_),
    .Q(\cpuregs[1] [11]),
    .QN(_28402_)
  );
  DFF_X1 cpuregs_reg_1__12_  (
    .CK(clk),
    .D(_00787_),
    .Q(\cpuregs[1] [12]),
    .QN(_28401_)
  );
  DFF_X1 cpuregs_reg_1__13_  (
    .CK(clk),
    .D(_00788_),
    .Q(\cpuregs[1] [13]),
    .QN(_28400_)
  );
  DFF_X1 cpuregs_reg_1__14_  (
    .CK(clk),
    .D(_00789_),
    .Q(\cpuregs[1] [14]),
    .QN(_28399_)
  );
  DFF_X1 cpuregs_reg_1__15_  (
    .CK(clk),
    .D(_00790_),
    .Q(\cpuregs[1] [15]),
    .QN(_28398_)
  );
  DFF_X1 cpuregs_reg_1__16_  (
    .CK(clk),
    .D(_00791_),
    .Q(\cpuregs[1] [16]),
    .QN(_28397_)
  );
  DFF_X1 cpuregs_reg_1__17_  (
    .CK(clk),
    .D(_00792_),
    .Q(\cpuregs[1] [17]),
    .QN(_28396_)
  );
  DFF_X1 cpuregs_reg_1__18_  (
    .CK(clk),
    .D(_00793_),
    .Q(\cpuregs[1] [18]),
    .QN(_28395_)
  );
  DFF_X1 cpuregs_reg_1__19_  (
    .CK(clk),
    .D(_00794_),
    .Q(\cpuregs[1] [19]),
    .QN(_28394_)
  );
  DFF_X1 cpuregs_reg_1__1_  (
    .CK(clk),
    .D(_00776_),
    .Q(\cpuregs[1] [1]),
    .QN(_28412_)
  );
  DFF_X1 cpuregs_reg_1__20_  (
    .CK(clk),
    .D(_00795_),
    .Q(\cpuregs[1] [20]),
    .QN(_28393_)
  );
  DFF_X1 cpuregs_reg_1__21_  (
    .CK(clk),
    .D(_00796_),
    .Q(\cpuregs[1] [21]),
    .QN(_28392_)
  );
  DFF_X1 cpuregs_reg_1__22_  (
    .CK(clk),
    .D(_00797_),
    .Q(\cpuregs[1] [22]),
    .QN(_28391_)
  );
  DFF_X1 cpuregs_reg_1__23_  (
    .CK(clk),
    .D(_00798_),
    .Q(\cpuregs[1] [23]),
    .QN(_28390_)
  );
  DFF_X1 cpuregs_reg_1__24_  (
    .CK(clk),
    .D(_00799_),
    .Q(\cpuregs[1] [24]),
    .QN(_28389_)
  );
  DFF_X1 cpuregs_reg_1__25_  (
    .CK(clk),
    .D(_00800_),
    .Q(\cpuregs[1] [25]),
    .QN(_28388_)
  );
  DFF_X1 cpuregs_reg_1__26_  (
    .CK(clk),
    .D(_00801_),
    .Q(\cpuregs[1] [26]),
    .QN(_28387_)
  );
  DFF_X1 cpuregs_reg_1__27_  (
    .CK(clk),
    .D(_00802_),
    .Q(\cpuregs[1] [27]),
    .QN(_28386_)
  );
  DFF_X1 cpuregs_reg_1__28_  (
    .CK(clk),
    .D(_00803_),
    .Q(\cpuregs[1] [28]),
    .QN(_28385_)
  );
  DFF_X1 cpuregs_reg_1__29_  (
    .CK(clk),
    .D(_00804_),
    .Q(\cpuregs[1] [29]),
    .QN(_28384_)
  );
  DFF_X1 cpuregs_reg_1__2_  (
    .CK(clk),
    .D(_00777_),
    .Q(\cpuregs[1] [2]),
    .QN(_28411_)
  );
  DFF_X1 cpuregs_reg_1__30_  (
    .CK(clk),
    .D(_00805_),
    .Q(\cpuregs[1] [30]),
    .QN(_28383_)
  );
  DFF_X1 cpuregs_reg_1__31_  (
    .CK(clk),
    .D(_00515_),
    .Q(\cpuregs[1] [31]),
    .QN(_28673_)
  );
  DFF_X1 cpuregs_reg_1__3_  (
    .CK(clk),
    .D(_00778_),
    .Q(\cpuregs[1] [3]),
    .QN(_28410_)
  );
  DFF_X1 cpuregs_reg_1__4_  (
    .CK(clk),
    .D(_00779_),
    .Q(\cpuregs[1] [4]),
    .QN(_28409_)
  );
  DFF_X1 cpuregs_reg_1__5_  (
    .CK(clk),
    .D(_00780_),
    .Q(\cpuregs[1] [5]),
    .QN(_28408_)
  );
  DFF_X1 cpuregs_reg_1__6_  (
    .CK(clk),
    .D(_00781_),
    .Q(\cpuregs[1] [6]),
    .QN(_28407_)
  );
  DFF_X1 cpuregs_reg_1__7_  (
    .CK(clk),
    .D(_00782_),
    .Q(\cpuregs[1] [7]),
    .QN(_28406_)
  );
  DFF_X1 cpuregs_reg_1__8_  (
    .CK(clk),
    .D(_00783_),
    .Q(\cpuregs[1] [8]),
    .QN(_28405_)
  );
  DFF_X1 cpuregs_reg_1__9_  (
    .CK(clk),
    .D(_00784_),
    .Q(\cpuregs[1] [9]),
    .QN(_28404_)
  );
  DFF_X1 cpuregs_reg_20__0_  (
    .CK(clk),
    .D(_00992_),
    .Q(\cpuregs[20] [0]),
    .QN(_28196_)
  );
  DFF_X1 cpuregs_reg_20__10_  (
    .CK(clk),
    .D(_01002_),
    .Q(\cpuregs[20] [10]),
    .QN(_28186_)
  );
  DFF_X1 cpuregs_reg_20__11_  (
    .CK(clk),
    .D(_01003_),
    .Q(\cpuregs[20] [11]),
    .QN(_28185_)
  );
  DFF_X1 cpuregs_reg_20__12_  (
    .CK(clk),
    .D(_01004_),
    .Q(\cpuregs[20] [12]),
    .QN(_28184_)
  );
  DFF_X1 cpuregs_reg_20__13_  (
    .CK(clk),
    .D(_01005_),
    .Q(\cpuregs[20] [13]),
    .QN(_28183_)
  );
  DFF_X1 cpuregs_reg_20__14_  (
    .CK(clk),
    .D(_01006_),
    .Q(\cpuregs[20] [14]),
    .QN(_28182_)
  );
  DFF_X1 cpuregs_reg_20__15_  (
    .CK(clk),
    .D(_01007_),
    .Q(\cpuregs[20] [15]),
    .QN(_28181_)
  );
  DFF_X1 cpuregs_reg_20__16_  (
    .CK(clk),
    .D(_01008_),
    .Q(\cpuregs[20] [16]),
    .QN(_28180_)
  );
  DFF_X1 cpuregs_reg_20__17_  (
    .CK(clk),
    .D(_01009_),
    .Q(\cpuregs[20] [17]),
    .QN(_28179_)
  );
  DFF_X1 cpuregs_reg_20__18_  (
    .CK(clk),
    .D(_01010_),
    .Q(\cpuregs[20] [18]),
    .QN(_28178_)
  );
  DFF_X1 cpuregs_reg_20__19_  (
    .CK(clk),
    .D(_01011_),
    .Q(\cpuregs[20] [19]),
    .QN(_28177_)
  );
  DFF_X1 cpuregs_reg_20__1_  (
    .CK(clk),
    .D(_00993_),
    .Q(\cpuregs[20] [1]),
    .QN(_28195_)
  );
  DFF_X1 cpuregs_reg_20__20_  (
    .CK(clk),
    .D(_01012_),
    .Q(\cpuregs[20] [20]),
    .QN(_28176_)
  );
  DFF_X1 cpuregs_reg_20__21_  (
    .CK(clk),
    .D(_01013_),
    .Q(\cpuregs[20] [21]),
    .QN(_28175_)
  );
  DFF_X1 cpuregs_reg_20__22_  (
    .CK(clk),
    .D(_01014_),
    .Q(\cpuregs[20] [22]),
    .QN(_28174_)
  );
  DFF_X1 cpuregs_reg_20__23_  (
    .CK(clk),
    .D(_01015_),
    .Q(\cpuregs[20] [23]),
    .QN(_28173_)
  );
  DFF_X1 cpuregs_reg_20__24_  (
    .CK(clk),
    .D(_01016_),
    .Q(\cpuregs[20] [24]),
    .QN(_28172_)
  );
  DFF_X1 cpuregs_reg_20__25_  (
    .CK(clk),
    .D(_01017_),
    .Q(\cpuregs[20] [25]),
    .QN(_28171_)
  );
  DFF_X1 cpuregs_reg_20__26_  (
    .CK(clk),
    .D(_01018_),
    .Q(\cpuregs[20] [26]),
    .QN(_28170_)
  );
  DFF_X1 cpuregs_reg_20__27_  (
    .CK(clk),
    .D(_01019_),
    .Q(\cpuregs[20] [27]),
    .QN(_28169_)
  );
  DFF_X1 cpuregs_reg_20__28_  (
    .CK(clk),
    .D(_01020_),
    .Q(\cpuregs[20] [28]),
    .QN(_28168_)
  );
  DFF_X1 cpuregs_reg_20__29_  (
    .CK(clk),
    .D(_01021_),
    .Q(\cpuregs[20] [29]),
    .QN(_28167_)
  );
  DFF_X1 cpuregs_reg_20__2_  (
    .CK(clk),
    .D(_00994_),
    .Q(\cpuregs[20] [2]),
    .QN(_28194_)
  );
  DFF_X1 cpuregs_reg_20__30_  (
    .CK(clk),
    .D(_01022_),
    .Q(\cpuregs[20] [30]),
    .QN(_28166_)
  );
  DFF_X1 cpuregs_reg_20__31_  (
    .CK(clk),
    .D(_00514_),
    .Q(\cpuregs[20] [31]),
    .QN(_28674_)
  );
  DFF_X1 cpuregs_reg_20__3_  (
    .CK(clk),
    .D(_00995_),
    .Q(\cpuregs[20] [3]),
    .QN(_28193_)
  );
  DFF_X1 cpuregs_reg_20__4_  (
    .CK(clk),
    .D(_00996_),
    .Q(\cpuregs[20] [4]),
    .QN(_28192_)
  );
  DFF_X1 cpuregs_reg_20__5_  (
    .CK(clk),
    .D(_00997_),
    .Q(\cpuregs[20] [5]),
    .QN(_28191_)
  );
  DFF_X1 cpuregs_reg_20__6_  (
    .CK(clk),
    .D(_00998_),
    .Q(\cpuregs[20] [6]),
    .QN(_28190_)
  );
  DFF_X1 cpuregs_reg_20__7_  (
    .CK(clk),
    .D(_00999_),
    .Q(\cpuregs[20] [7]),
    .QN(_28189_)
  );
  DFF_X1 cpuregs_reg_20__8_  (
    .CK(clk),
    .D(_01000_),
    .Q(\cpuregs[20] [8]),
    .QN(_28188_)
  );
  DFF_X1 cpuregs_reg_20__9_  (
    .CK(clk),
    .D(_01001_),
    .Q(\cpuregs[20] [9]),
    .QN(_28187_)
  );
  DFF_X1 cpuregs_reg_21__0_  (
    .CK(clk),
    .D(_01178_),
    .Q(\cpuregs[21] [0]),
    .QN(_28010_)
  );
  DFF_X1 cpuregs_reg_21__10_  (
    .CK(clk),
    .D(_01188_),
    .Q(\cpuregs[21] [10]),
    .QN(_28000_)
  );
  DFF_X1 cpuregs_reg_21__11_  (
    .CK(clk),
    .D(_01189_),
    .Q(\cpuregs[21] [11]),
    .QN(_27999_)
  );
  DFF_X1 cpuregs_reg_21__12_  (
    .CK(clk),
    .D(_01190_),
    .Q(\cpuregs[21] [12]),
    .QN(_27998_)
  );
  DFF_X1 cpuregs_reg_21__13_  (
    .CK(clk),
    .D(_01191_),
    .Q(\cpuregs[21] [13]),
    .QN(_27997_)
  );
  DFF_X1 cpuregs_reg_21__14_  (
    .CK(clk),
    .D(_01192_),
    .Q(\cpuregs[21] [14]),
    .QN(_27996_)
  );
  DFF_X1 cpuregs_reg_21__15_  (
    .CK(clk),
    .D(_01193_),
    .Q(\cpuregs[21] [15]),
    .QN(_27995_)
  );
  DFF_X1 cpuregs_reg_21__16_  (
    .CK(clk),
    .D(_01194_),
    .Q(\cpuregs[21] [16]),
    .QN(_27994_)
  );
  DFF_X1 cpuregs_reg_21__17_  (
    .CK(clk),
    .D(_01195_),
    .Q(\cpuregs[21] [17]),
    .QN(_27993_)
  );
  DFF_X1 cpuregs_reg_21__18_  (
    .CK(clk),
    .D(_01196_),
    .Q(\cpuregs[21] [18]),
    .QN(_27992_)
  );
  DFF_X1 cpuregs_reg_21__19_  (
    .CK(clk),
    .D(_01197_),
    .Q(\cpuregs[21] [19]),
    .QN(_27991_)
  );
  DFF_X1 cpuregs_reg_21__1_  (
    .CK(clk),
    .D(_01179_),
    .Q(\cpuregs[21] [1]),
    .QN(_28009_)
  );
  DFF_X1 cpuregs_reg_21__20_  (
    .CK(clk),
    .D(_01198_),
    .Q(\cpuregs[21] [20]),
    .QN(_27990_)
  );
  DFF_X1 cpuregs_reg_21__21_  (
    .CK(clk),
    .D(_01199_),
    .Q(\cpuregs[21] [21]),
    .QN(_27989_)
  );
  DFF_X1 cpuregs_reg_21__22_  (
    .CK(clk),
    .D(_01200_),
    .Q(\cpuregs[21] [22]),
    .QN(_27988_)
  );
  DFF_X1 cpuregs_reg_21__23_  (
    .CK(clk),
    .D(_01201_),
    .Q(\cpuregs[21] [23]),
    .QN(_27987_)
  );
  DFF_X1 cpuregs_reg_21__24_  (
    .CK(clk),
    .D(_01202_),
    .Q(\cpuregs[21] [24]),
    .QN(_27986_)
  );
  DFF_X1 cpuregs_reg_21__25_  (
    .CK(clk),
    .D(_01203_),
    .Q(\cpuregs[21] [25]),
    .QN(_27985_)
  );
  DFF_X1 cpuregs_reg_21__26_  (
    .CK(clk),
    .D(_01204_),
    .Q(\cpuregs[21] [26]),
    .QN(_27984_)
  );
  DFF_X1 cpuregs_reg_21__27_  (
    .CK(clk),
    .D(_01205_),
    .Q(\cpuregs[21] [27]),
    .QN(_27983_)
  );
  DFF_X1 cpuregs_reg_21__28_  (
    .CK(clk),
    .D(_01206_),
    .Q(\cpuregs[21] [28]),
    .QN(_27982_)
  );
  DFF_X1 cpuregs_reg_21__29_  (
    .CK(clk),
    .D(_01207_),
    .Q(\cpuregs[21] [29]),
    .QN(_27981_)
  );
  DFF_X1 cpuregs_reg_21__2_  (
    .CK(clk),
    .D(_01180_),
    .Q(\cpuregs[21] [2]),
    .QN(_28008_)
  );
  DFF_X1 cpuregs_reg_21__30_  (
    .CK(clk),
    .D(_01208_),
    .Q(\cpuregs[21] [30]),
    .QN(_27980_)
  );
  DFF_X1 cpuregs_reg_21__31_  (
    .CK(clk),
    .D(_00513_),
    .Q(\cpuregs[21] [31]),
    .QN(_28675_)
  );
  DFF_X1 cpuregs_reg_21__3_  (
    .CK(clk),
    .D(_01181_),
    .Q(\cpuregs[21] [3]),
    .QN(_28007_)
  );
  DFF_X1 cpuregs_reg_21__4_  (
    .CK(clk),
    .D(_01182_),
    .Q(\cpuregs[21] [4]),
    .QN(_28006_)
  );
  DFF_X1 cpuregs_reg_21__5_  (
    .CK(clk),
    .D(_01183_),
    .Q(\cpuregs[21] [5]),
    .QN(_28005_)
  );
  DFF_X1 cpuregs_reg_21__6_  (
    .CK(clk),
    .D(_01184_),
    .Q(\cpuregs[21] [6]),
    .QN(_28004_)
  );
  DFF_X1 cpuregs_reg_21__7_  (
    .CK(clk),
    .D(_01185_),
    .Q(\cpuregs[21] [7]),
    .QN(_28003_)
  );
  DFF_X1 cpuregs_reg_21__8_  (
    .CK(clk),
    .D(_01186_),
    .Q(\cpuregs[21] [8]),
    .QN(_28002_)
  );
  DFF_X1 cpuregs_reg_21__9_  (
    .CK(clk),
    .D(_01187_),
    .Q(\cpuregs[21] [9]),
    .QN(_28001_)
  );
  DFF_X1 cpuregs_reg_22__0_  (
    .CK(clk),
    .D(_00620_),
    .Q(\cpuregs[22] [0]),
    .QN(_28568_)
  );
  DFF_X1 cpuregs_reg_22__10_  (
    .CK(clk),
    .D(_00630_),
    .Q(\cpuregs[22] [10]),
    .QN(_28558_)
  );
  DFF_X1 cpuregs_reg_22__11_  (
    .CK(clk),
    .D(_00631_),
    .Q(\cpuregs[22] [11]),
    .QN(_28557_)
  );
  DFF_X1 cpuregs_reg_22__12_  (
    .CK(clk),
    .D(_00632_),
    .Q(\cpuregs[22] [12]),
    .QN(_28556_)
  );
  DFF_X1 cpuregs_reg_22__13_  (
    .CK(clk),
    .D(_00633_),
    .Q(\cpuregs[22] [13]),
    .QN(_28555_)
  );
  DFF_X1 cpuregs_reg_22__14_  (
    .CK(clk),
    .D(_00634_),
    .Q(\cpuregs[22] [14]),
    .QN(_28554_)
  );
  DFF_X1 cpuregs_reg_22__15_  (
    .CK(clk),
    .D(_00635_),
    .Q(\cpuregs[22] [15]),
    .QN(_28553_)
  );
  DFF_X1 cpuregs_reg_22__16_  (
    .CK(clk),
    .D(_00636_),
    .Q(\cpuregs[22] [16]),
    .QN(_28552_)
  );
  DFF_X1 cpuregs_reg_22__17_  (
    .CK(clk),
    .D(_00637_),
    .Q(\cpuregs[22] [17]),
    .QN(_28551_)
  );
  DFF_X1 cpuregs_reg_22__18_  (
    .CK(clk),
    .D(_00638_),
    .Q(\cpuregs[22] [18]),
    .QN(_28550_)
  );
  DFF_X1 cpuregs_reg_22__19_  (
    .CK(clk),
    .D(_00639_),
    .Q(\cpuregs[22] [19]),
    .QN(_28549_)
  );
  DFF_X1 cpuregs_reg_22__1_  (
    .CK(clk),
    .D(_00621_),
    .Q(\cpuregs[22] [1]),
    .QN(_28567_)
  );
  DFF_X1 cpuregs_reg_22__20_  (
    .CK(clk),
    .D(_00640_),
    .Q(\cpuregs[22] [20]),
    .QN(_28548_)
  );
  DFF_X1 cpuregs_reg_22__21_  (
    .CK(clk),
    .D(_00641_),
    .Q(\cpuregs[22] [21]),
    .QN(_28547_)
  );
  DFF_X1 cpuregs_reg_22__22_  (
    .CK(clk),
    .D(_00642_),
    .Q(\cpuregs[22] [22]),
    .QN(_28546_)
  );
  DFF_X1 cpuregs_reg_22__23_  (
    .CK(clk),
    .D(_00643_),
    .Q(\cpuregs[22] [23]),
    .QN(_28545_)
  );
  DFF_X1 cpuregs_reg_22__24_  (
    .CK(clk),
    .D(_00644_),
    .Q(\cpuregs[22] [24]),
    .QN(_28544_)
  );
  DFF_X1 cpuregs_reg_22__25_  (
    .CK(clk),
    .D(_00645_),
    .Q(\cpuregs[22] [25]),
    .QN(_28543_)
  );
  DFF_X1 cpuregs_reg_22__26_  (
    .CK(clk),
    .D(_00646_),
    .Q(\cpuregs[22] [26]),
    .QN(_28542_)
  );
  DFF_X1 cpuregs_reg_22__27_  (
    .CK(clk),
    .D(_00647_),
    .Q(\cpuregs[22] [27]),
    .QN(_28541_)
  );
  DFF_X1 cpuregs_reg_22__28_  (
    .CK(clk),
    .D(_00648_),
    .Q(\cpuregs[22] [28]),
    .QN(_28540_)
  );
  DFF_X1 cpuregs_reg_22__29_  (
    .CK(clk),
    .D(_00649_),
    .Q(\cpuregs[22] [29]),
    .QN(_28539_)
  );
  DFF_X1 cpuregs_reg_22__2_  (
    .CK(clk),
    .D(_00622_),
    .Q(\cpuregs[22] [2]),
    .QN(_28566_)
  );
  DFF_X1 cpuregs_reg_22__30_  (
    .CK(clk),
    .D(_00650_),
    .Q(\cpuregs[22] [30]),
    .QN(_28538_)
  );
  DFF_X1 cpuregs_reg_22__31_  (
    .CK(clk),
    .D(_00512_),
    .Q(\cpuregs[22] [31]),
    .QN(_28676_)
  );
  DFF_X1 cpuregs_reg_22__3_  (
    .CK(clk),
    .D(_00623_),
    .Q(\cpuregs[22] [3]),
    .QN(_28565_)
  );
  DFF_X1 cpuregs_reg_22__4_  (
    .CK(clk),
    .D(_00624_),
    .Q(\cpuregs[22] [4]),
    .QN(_28564_)
  );
  DFF_X1 cpuregs_reg_22__5_  (
    .CK(clk),
    .D(_00625_),
    .Q(\cpuregs[22] [5]),
    .QN(_28563_)
  );
  DFF_X1 cpuregs_reg_22__6_  (
    .CK(clk),
    .D(_00626_),
    .Q(\cpuregs[22] [6]),
    .QN(_28562_)
  );
  DFF_X1 cpuregs_reg_22__7_  (
    .CK(clk),
    .D(_00627_),
    .Q(\cpuregs[22] [7]),
    .QN(_28561_)
  );
  DFF_X1 cpuregs_reg_22__8_  (
    .CK(clk),
    .D(_00628_),
    .Q(\cpuregs[22] [8]),
    .QN(_28560_)
  );
  DFF_X1 cpuregs_reg_22__9_  (
    .CK(clk),
    .D(_00629_),
    .Q(\cpuregs[22] [9]),
    .QN(_28559_)
  );
  DFF_X1 cpuregs_reg_23__0_  (
    .CK(clk),
    .D(_00527_),
    .Q(\cpuregs[23] [0]),
    .QN(_28661_)
  );
  DFF_X1 cpuregs_reg_23__10_  (
    .CK(clk),
    .D(_00537_),
    .Q(\cpuregs[23] [10]),
    .QN(_28651_)
  );
  DFF_X1 cpuregs_reg_23__11_  (
    .CK(clk),
    .D(_00538_),
    .Q(\cpuregs[23] [11]),
    .QN(_28650_)
  );
  DFF_X1 cpuregs_reg_23__12_  (
    .CK(clk),
    .D(_00539_),
    .Q(\cpuregs[23] [12]),
    .QN(_28649_)
  );
  DFF_X1 cpuregs_reg_23__13_  (
    .CK(clk),
    .D(_00540_),
    .Q(\cpuregs[23] [13]),
    .QN(_28648_)
  );
  DFF_X1 cpuregs_reg_23__14_  (
    .CK(clk),
    .D(_00541_),
    .Q(\cpuregs[23] [14]),
    .QN(_28647_)
  );
  DFF_X1 cpuregs_reg_23__15_  (
    .CK(clk),
    .D(_00542_),
    .Q(\cpuregs[23] [15]),
    .QN(_28646_)
  );
  DFF_X1 cpuregs_reg_23__16_  (
    .CK(clk),
    .D(_00543_),
    .Q(\cpuregs[23] [16]),
    .QN(_28645_)
  );
  DFF_X1 cpuregs_reg_23__17_  (
    .CK(clk),
    .D(_00544_),
    .Q(\cpuregs[23] [17]),
    .QN(_28644_)
  );
  DFF_X1 cpuregs_reg_23__18_  (
    .CK(clk),
    .D(_00545_),
    .Q(\cpuregs[23] [18]),
    .QN(_28643_)
  );
  DFF_X1 cpuregs_reg_23__19_  (
    .CK(clk),
    .D(_00546_),
    .Q(\cpuregs[23] [19]),
    .QN(_28642_)
  );
  DFF_X1 cpuregs_reg_23__1_  (
    .CK(clk),
    .D(_00528_),
    .Q(\cpuregs[23] [1]),
    .QN(_28660_)
  );
  DFF_X1 cpuregs_reg_23__20_  (
    .CK(clk),
    .D(_00547_),
    .Q(\cpuregs[23] [20]),
    .QN(_28641_)
  );
  DFF_X1 cpuregs_reg_23__21_  (
    .CK(clk),
    .D(_00548_),
    .Q(\cpuregs[23] [21]),
    .QN(_28640_)
  );
  DFF_X1 cpuregs_reg_23__22_  (
    .CK(clk),
    .D(_00549_),
    .Q(\cpuregs[23] [22]),
    .QN(_28639_)
  );
  DFF_X1 cpuregs_reg_23__23_  (
    .CK(clk),
    .D(_00550_),
    .Q(\cpuregs[23] [23]),
    .QN(_28638_)
  );
  DFF_X1 cpuregs_reg_23__24_  (
    .CK(clk),
    .D(_00551_),
    .Q(\cpuregs[23] [24]),
    .QN(_28637_)
  );
  DFF_X1 cpuregs_reg_23__25_  (
    .CK(clk),
    .D(_00552_),
    .Q(\cpuregs[23] [25]),
    .QN(_28636_)
  );
  DFF_X1 cpuregs_reg_23__26_  (
    .CK(clk),
    .D(_00553_),
    .Q(\cpuregs[23] [26]),
    .QN(_28635_)
  );
  DFF_X1 cpuregs_reg_23__27_  (
    .CK(clk),
    .D(_00554_),
    .Q(\cpuregs[23] [27]),
    .QN(_28634_)
  );
  DFF_X1 cpuregs_reg_23__28_  (
    .CK(clk),
    .D(_00555_),
    .Q(\cpuregs[23] [28]),
    .QN(_28633_)
  );
  DFF_X1 cpuregs_reg_23__29_  (
    .CK(clk),
    .D(_00556_),
    .Q(\cpuregs[23] [29]),
    .QN(_28632_)
  );
  DFF_X1 cpuregs_reg_23__2_  (
    .CK(clk),
    .D(_00529_),
    .Q(\cpuregs[23] [2]),
    .QN(_28659_)
  );
  DFF_X1 cpuregs_reg_23__30_  (
    .CK(clk),
    .D(_00557_),
    .Q(\cpuregs[23] [30]),
    .QN(_28631_)
  );
  DFF_X1 cpuregs_reg_23__31_  (
    .CK(clk),
    .D(_00511_),
    .Q(\cpuregs[23] [31]),
    .QN(_28677_)
  );
  DFF_X1 cpuregs_reg_23__3_  (
    .CK(clk),
    .D(_00530_),
    .Q(\cpuregs[23] [3]),
    .QN(_28658_)
  );
  DFF_X1 cpuregs_reg_23__4_  (
    .CK(clk),
    .D(_00531_),
    .Q(\cpuregs[23] [4]),
    .QN(_28657_)
  );
  DFF_X1 cpuregs_reg_23__5_  (
    .CK(clk),
    .D(_00532_),
    .Q(\cpuregs[23] [5]),
    .QN(_28656_)
  );
  DFF_X1 cpuregs_reg_23__6_  (
    .CK(clk),
    .D(_00533_),
    .Q(\cpuregs[23] [6]),
    .QN(_28655_)
  );
  DFF_X1 cpuregs_reg_23__7_  (
    .CK(clk),
    .D(_00534_),
    .Q(\cpuregs[23] [7]),
    .QN(_28654_)
  );
  DFF_X1 cpuregs_reg_23__8_  (
    .CK(clk),
    .D(_00535_),
    .Q(\cpuregs[23] [8]),
    .QN(_28653_)
  );
  DFF_X1 cpuregs_reg_23__9_  (
    .CK(clk),
    .D(_00536_),
    .Q(\cpuregs[23] [9]),
    .QN(_28652_)
  );
  DFF_X1 cpuregs_reg_24__0_  (
    .CK(clk),
    .D(_00837_),
    .Q(\cpuregs[24] [0]),
    .QN(_28351_)
  );
  DFF_X1 cpuregs_reg_24__10_  (
    .CK(clk),
    .D(_00847_),
    .Q(\cpuregs[24] [10]),
    .QN(_28341_)
  );
  DFF_X1 cpuregs_reg_24__11_  (
    .CK(clk),
    .D(_00848_),
    .Q(\cpuregs[24] [11]),
    .QN(_28340_)
  );
  DFF_X1 cpuregs_reg_24__12_  (
    .CK(clk),
    .D(_00849_),
    .Q(\cpuregs[24] [12]),
    .QN(_28339_)
  );
  DFF_X1 cpuregs_reg_24__13_  (
    .CK(clk),
    .D(_00850_),
    .Q(\cpuregs[24] [13]),
    .QN(_28338_)
  );
  DFF_X1 cpuregs_reg_24__14_  (
    .CK(clk),
    .D(_00851_),
    .Q(\cpuregs[24] [14]),
    .QN(_28337_)
  );
  DFF_X1 cpuregs_reg_24__15_  (
    .CK(clk),
    .D(_00852_),
    .Q(\cpuregs[24] [15]),
    .QN(_28336_)
  );
  DFF_X1 cpuregs_reg_24__16_  (
    .CK(clk),
    .D(_00853_),
    .Q(\cpuregs[24] [16]),
    .QN(_28335_)
  );
  DFF_X1 cpuregs_reg_24__17_  (
    .CK(clk),
    .D(_00854_),
    .Q(\cpuregs[24] [17]),
    .QN(_28334_)
  );
  DFF_X1 cpuregs_reg_24__18_  (
    .CK(clk),
    .D(_00855_),
    .Q(\cpuregs[24] [18]),
    .QN(_28333_)
  );
  DFF_X1 cpuregs_reg_24__19_  (
    .CK(clk),
    .D(_00856_),
    .Q(\cpuregs[24] [19]),
    .QN(_28332_)
  );
  DFF_X1 cpuregs_reg_24__1_  (
    .CK(clk),
    .D(_00838_),
    .Q(\cpuregs[24] [1]),
    .QN(_28350_)
  );
  DFF_X1 cpuregs_reg_24__20_  (
    .CK(clk),
    .D(_00857_),
    .Q(\cpuregs[24] [20]),
    .QN(_28331_)
  );
  DFF_X1 cpuregs_reg_24__21_  (
    .CK(clk),
    .D(_00858_),
    .Q(\cpuregs[24] [21]),
    .QN(_28330_)
  );
  DFF_X1 cpuregs_reg_24__22_  (
    .CK(clk),
    .D(_00859_),
    .Q(\cpuregs[24] [22]),
    .QN(_28329_)
  );
  DFF_X1 cpuregs_reg_24__23_  (
    .CK(clk),
    .D(_00860_),
    .Q(\cpuregs[24] [23]),
    .QN(_28328_)
  );
  DFF_X1 cpuregs_reg_24__24_  (
    .CK(clk),
    .D(_00861_),
    .Q(\cpuregs[24] [24]),
    .QN(_28327_)
  );
  DFF_X1 cpuregs_reg_24__25_  (
    .CK(clk),
    .D(_00862_),
    .Q(\cpuregs[24] [25]),
    .QN(_28326_)
  );
  DFF_X1 cpuregs_reg_24__26_  (
    .CK(clk),
    .D(_00863_),
    .Q(\cpuregs[24] [26]),
    .QN(_28325_)
  );
  DFF_X1 cpuregs_reg_24__27_  (
    .CK(clk),
    .D(_00864_),
    .Q(\cpuregs[24] [27]),
    .QN(_28324_)
  );
  DFF_X1 cpuregs_reg_24__28_  (
    .CK(clk),
    .D(_00865_),
    .Q(\cpuregs[24] [28]),
    .QN(_28323_)
  );
  DFF_X1 cpuregs_reg_24__29_  (
    .CK(clk),
    .D(_00866_),
    .Q(\cpuregs[24] [29]),
    .QN(_28322_)
  );
  DFF_X1 cpuregs_reg_24__2_  (
    .CK(clk),
    .D(_00839_),
    .Q(\cpuregs[24] [2]),
    .QN(_28349_)
  );
  DFF_X1 cpuregs_reg_24__30_  (
    .CK(clk),
    .D(_00867_),
    .Q(\cpuregs[24] [30]),
    .QN(_28321_)
  );
  DFF_X1 cpuregs_reg_24__31_  (
    .CK(clk),
    .D(_00510_),
    .Q(\cpuregs[24] [31]),
    .QN(_28678_)
  );
  DFF_X1 cpuregs_reg_24__3_  (
    .CK(clk),
    .D(_00840_),
    .Q(\cpuregs[24] [3]),
    .QN(_28348_)
  );
  DFF_X1 cpuregs_reg_24__4_  (
    .CK(clk),
    .D(_00841_),
    .Q(\cpuregs[24] [4]),
    .QN(_28347_)
  );
  DFF_X1 cpuregs_reg_24__5_  (
    .CK(clk),
    .D(_00842_),
    .Q(\cpuregs[24] [5]),
    .QN(_28346_)
  );
  DFF_X1 cpuregs_reg_24__6_  (
    .CK(clk),
    .D(_00843_),
    .Q(\cpuregs[24] [6]),
    .QN(_28345_)
  );
  DFF_X1 cpuregs_reg_24__7_  (
    .CK(clk),
    .D(_00844_),
    .Q(\cpuregs[24] [7]),
    .QN(_28344_)
  );
  DFF_X1 cpuregs_reg_24__8_  (
    .CK(clk),
    .D(_00845_),
    .Q(\cpuregs[24] [8]),
    .QN(_28343_)
  );
  DFF_X1 cpuregs_reg_24__9_  (
    .CK(clk),
    .D(_00846_),
    .Q(\cpuregs[24] [9]),
    .QN(_28342_)
  );
  DFF_X1 cpuregs_reg_25__0_  (
    .CK(clk),
    .D(_01271_),
    .Q(\cpuregs[25] [0]),
    .QN(_27917_)
  );
  DFF_X1 cpuregs_reg_25__10_  (
    .CK(clk),
    .D(_01281_),
    .Q(\cpuregs[25] [10]),
    .QN(_27907_)
  );
  DFF_X1 cpuregs_reg_25__11_  (
    .CK(clk),
    .D(_01282_),
    .Q(\cpuregs[25] [11]),
    .QN(_27906_)
  );
  DFF_X1 cpuregs_reg_25__12_  (
    .CK(clk),
    .D(_01283_),
    .Q(\cpuregs[25] [12]),
    .QN(_27905_)
  );
  DFF_X1 cpuregs_reg_25__13_  (
    .CK(clk),
    .D(_01284_),
    .Q(\cpuregs[25] [13]),
    .QN(_27904_)
  );
  DFF_X1 cpuregs_reg_25__14_  (
    .CK(clk),
    .D(_01285_),
    .Q(\cpuregs[25] [14]),
    .QN(_27903_)
  );
  DFF_X1 cpuregs_reg_25__15_  (
    .CK(clk),
    .D(_01286_),
    .Q(\cpuregs[25] [15]),
    .QN(_27902_)
  );
  DFF_X1 cpuregs_reg_25__16_  (
    .CK(clk),
    .D(_01287_),
    .Q(\cpuregs[25] [16]),
    .QN(_27901_)
  );
  DFF_X1 cpuregs_reg_25__17_  (
    .CK(clk),
    .D(_01288_),
    .Q(\cpuregs[25] [17]),
    .QN(_27900_)
  );
  DFF_X1 cpuregs_reg_25__18_  (
    .CK(clk),
    .D(_01289_),
    .Q(\cpuregs[25] [18]),
    .QN(_27899_)
  );
  DFF_X1 cpuregs_reg_25__19_  (
    .CK(clk),
    .D(_01290_),
    .Q(\cpuregs[25] [19]),
    .QN(_27898_)
  );
  DFF_X1 cpuregs_reg_25__1_  (
    .CK(clk),
    .D(_01272_),
    .Q(\cpuregs[25] [1]),
    .QN(_27916_)
  );
  DFF_X1 cpuregs_reg_25__20_  (
    .CK(clk),
    .D(_01291_),
    .Q(\cpuregs[25] [20]),
    .QN(_27897_)
  );
  DFF_X1 cpuregs_reg_25__21_  (
    .CK(clk),
    .D(_01292_),
    .Q(\cpuregs[25] [21]),
    .QN(_27896_)
  );
  DFF_X1 cpuregs_reg_25__22_  (
    .CK(clk),
    .D(_01293_),
    .Q(\cpuregs[25] [22]),
    .QN(_27895_)
  );
  DFF_X1 cpuregs_reg_25__23_  (
    .CK(clk),
    .D(_01294_),
    .Q(\cpuregs[25] [23]),
    .QN(_27894_)
  );
  DFF_X1 cpuregs_reg_25__24_  (
    .CK(clk),
    .D(_01295_),
    .Q(\cpuregs[25] [24]),
    .QN(_27893_)
  );
  DFF_X1 cpuregs_reg_25__25_  (
    .CK(clk),
    .D(_01296_),
    .Q(\cpuregs[25] [25]),
    .QN(_27892_)
  );
  DFF_X1 cpuregs_reg_25__26_  (
    .CK(clk),
    .D(_01297_),
    .Q(\cpuregs[25] [26]),
    .QN(_27891_)
  );
  DFF_X1 cpuregs_reg_25__27_  (
    .CK(clk),
    .D(_01298_),
    .Q(\cpuregs[25] [27]),
    .QN(_27890_)
  );
  DFF_X1 cpuregs_reg_25__28_  (
    .CK(clk),
    .D(_01299_),
    .Q(\cpuregs[25] [28]),
    .QN(_27889_)
  );
  DFF_X1 cpuregs_reg_25__29_  (
    .CK(clk),
    .D(_01300_),
    .Q(\cpuregs[25] [29]),
    .QN(_27888_)
  );
  DFF_X1 cpuregs_reg_25__2_  (
    .CK(clk),
    .D(_01273_),
    .Q(\cpuregs[25] [2]),
    .QN(_27915_)
  );
  DFF_X1 cpuregs_reg_25__30_  (
    .CK(clk),
    .D(_01301_),
    .Q(\cpuregs[25] [30]),
    .QN(_27887_)
  );
  DFF_X1 cpuregs_reg_25__31_  (
    .CK(clk),
    .D(_00509_),
    .Q(\cpuregs[25] [31]),
    .QN(_28679_)
  );
  DFF_X1 cpuregs_reg_25__3_  (
    .CK(clk),
    .D(_01274_),
    .Q(\cpuregs[25] [3]),
    .QN(_27914_)
  );
  DFF_X1 cpuregs_reg_25__4_  (
    .CK(clk),
    .D(_01275_),
    .Q(\cpuregs[25] [4]),
    .QN(_27913_)
  );
  DFF_X1 cpuregs_reg_25__5_  (
    .CK(clk),
    .D(_01276_),
    .Q(\cpuregs[25] [5]),
    .QN(_27912_)
  );
  DFF_X1 cpuregs_reg_25__6_  (
    .CK(clk),
    .D(_01277_),
    .Q(\cpuregs[25] [6]),
    .QN(_27911_)
  );
  DFF_X1 cpuregs_reg_25__7_  (
    .CK(clk),
    .D(_01278_),
    .Q(\cpuregs[25] [7]),
    .QN(_27910_)
  );
  DFF_X1 cpuregs_reg_25__8_  (
    .CK(clk),
    .D(_01279_),
    .Q(\cpuregs[25] [8]),
    .QN(_27909_)
  );
  DFF_X1 cpuregs_reg_25__9_  (
    .CK(clk),
    .D(_01280_),
    .Q(\cpuregs[25] [9]),
    .QN(_27908_)
  );
  DFF_X1 cpuregs_reg_26__0_  (
    .CK(clk),
    .D(_01333_),
    .Q(\cpuregs[26] [0]),
    .QN(_27855_)
  );
  DFF_X1 cpuregs_reg_26__10_  (
    .CK(clk),
    .D(_01343_),
    .Q(\cpuregs[26] [10]),
    .QN(_27845_)
  );
  DFF_X1 cpuregs_reg_26__11_  (
    .CK(clk),
    .D(_01344_),
    .Q(\cpuregs[26] [11]),
    .QN(_27844_)
  );
  DFF_X1 cpuregs_reg_26__12_  (
    .CK(clk),
    .D(_01345_),
    .Q(\cpuregs[26] [12]),
    .QN(_27843_)
  );
  DFF_X1 cpuregs_reg_26__13_  (
    .CK(clk),
    .D(_01346_),
    .Q(\cpuregs[26] [13]),
    .QN(_27842_)
  );
  DFF_X1 cpuregs_reg_26__14_  (
    .CK(clk),
    .D(_01347_),
    .Q(\cpuregs[26] [14]),
    .QN(_27841_)
  );
  DFF_X1 cpuregs_reg_26__15_  (
    .CK(clk),
    .D(_01348_),
    .Q(\cpuregs[26] [15]),
    .QN(_27840_)
  );
  DFF_X1 cpuregs_reg_26__16_  (
    .CK(clk),
    .D(_01349_),
    .Q(\cpuregs[26] [16]),
    .QN(_27839_)
  );
  DFF_X1 cpuregs_reg_26__17_  (
    .CK(clk),
    .D(_01350_),
    .Q(\cpuregs[26] [17]),
    .QN(_27838_)
  );
  DFF_X1 cpuregs_reg_26__18_  (
    .CK(clk),
    .D(_01351_),
    .Q(\cpuregs[26] [18]),
    .QN(_27837_)
  );
  DFF_X1 cpuregs_reg_26__19_  (
    .CK(clk),
    .D(_01352_),
    .Q(\cpuregs[26] [19]),
    .QN(_27836_)
  );
  DFF_X1 cpuregs_reg_26__1_  (
    .CK(clk),
    .D(_01334_),
    .Q(\cpuregs[26] [1]),
    .QN(_27854_)
  );
  DFF_X1 cpuregs_reg_26__20_  (
    .CK(clk),
    .D(_01353_),
    .Q(\cpuregs[26] [20]),
    .QN(_27835_)
  );
  DFF_X1 cpuregs_reg_26__21_  (
    .CK(clk),
    .D(_01354_),
    .Q(\cpuregs[26] [21]),
    .QN(_27834_)
  );
  DFF_X1 cpuregs_reg_26__22_  (
    .CK(clk),
    .D(_01355_),
    .Q(\cpuregs[26] [22]),
    .QN(_27833_)
  );
  DFF_X1 cpuregs_reg_26__23_  (
    .CK(clk),
    .D(_01356_),
    .Q(\cpuregs[26] [23]),
    .QN(_27832_)
  );
  DFF_X1 cpuregs_reg_26__24_  (
    .CK(clk),
    .D(_01357_),
    .Q(\cpuregs[26] [24]),
    .QN(_27831_)
  );
  DFF_X1 cpuregs_reg_26__25_  (
    .CK(clk),
    .D(_01358_),
    .Q(\cpuregs[26] [25]),
    .QN(_27830_)
  );
  DFF_X1 cpuregs_reg_26__26_  (
    .CK(clk),
    .D(_01359_),
    .Q(\cpuregs[26] [26]),
    .QN(_27829_)
  );
  DFF_X1 cpuregs_reg_26__27_  (
    .CK(clk),
    .D(_01360_),
    .Q(\cpuregs[26] [27]),
    .QN(_27828_)
  );
  DFF_X1 cpuregs_reg_26__28_  (
    .CK(clk),
    .D(_01361_),
    .Q(\cpuregs[26] [28]),
    .QN(_27827_)
  );
  DFF_X1 cpuregs_reg_26__29_  (
    .CK(clk),
    .D(_01362_),
    .Q(\cpuregs[26] [29]),
    .QN(_27826_)
  );
  DFF_X1 cpuregs_reg_26__2_  (
    .CK(clk),
    .D(_01335_),
    .Q(\cpuregs[26] [2]),
    .QN(_27853_)
  );
  DFF_X1 cpuregs_reg_26__30_  (
    .CK(clk),
    .D(_01363_),
    .Q(\cpuregs[26] [30]),
    .QN(_27825_)
  );
  DFF_X1 cpuregs_reg_26__31_  (
    .CK(clk),
    .D(_00508_),
    .Q(\cpuregs[26] [31]),
    .QN(_28680_)
  );
  DFF_X1 cpuregs_reg_26__3_  (
    .CK(clk),
    .D(_01336_),
    .Q(\cpuregs[26] [3]),
    .QN(_27852_)
  );
  DFF_X1 cpuregs_reg_26__4_  (
    .CK(clk),
    .D(_01337_),
    .Q(\cpuregs[26] [4]),
    .QN(_27851_)
  );
  DFF_X1 cpuregs_reg_26__5_  (
    .CK(clk),
    .D(_01338_),
    .Q(\cpuregs[26] [5]),
    .QN(_27850_)
  );
  DFF_X1 cpuregs_reg_26__6_  (
    .CK(clk),
    .D(_01339_),
    .Q(\cpuregs[26] [6]),
    .QN(_27849_)
  );
  DFF_X1 cpuregs_reg_26__7_  (
    .CK(clk),
    .D(_01340_),
    .Q(\cpuregs[26] [7]),
    .QN(_27848_)
  );
  DFF_X1 cpuregs_reg_26__8_  (
    .CK(clk),
    .D(_01341_),
    .Q(\cpuregs[26] [8]),
    .QN(_27847_)
  );
  DFF_X1 cpuregs_reg_26__9_  (
    .CK(clk),
    .D(_01342_),
    .Q(\cpuregs[26] [9]),
    .QN(_27846_)
  );
  DFF_X1 cpuregs_reg_27__0_  (
    .CK(clk),
    .D(_01426_),
    .Q(\cpuregs[27] [0]),
    .QN(_27762_)
  );
  DFF_X1 cpuregs_reg_27__10_  (
    .CK(clk),
    .D(_01436_),
    .Q(\cpuregs[27] [10]),
    .QN(_27752_)
  );
  DFF_X1 cpuregs_reg_27__11_  (
    .CK(clk),
    .D(_01437_),
    .Q(\cpuregs[27] [11]),
    .QN(_27751_)
  );
  DFF_X1 cpuregs_reg_27__12_  (
    .CK(clk),
    .D(_01438_),
    .Q(\cpuregs[27] [12]),
    .QN(_27750_)
  );
  DFF_X1 cpuregs_reg_27__13_  (
    .CK(clk),
    .D(_01439_),
    .Q(\cpuregs[27] [13]),
    .QN(_27749_)
  );
  DFF_X1 cpuregs_reg_27__14_  (
    .CK(clk),
    .D(_01440_),
    .Q(\cpuregs[27] [14]),
    .QN(_27748_)
  );
  DFF_X1 cpuregs_reg_27__15_  (
    .CK(clk),
    .D(_01441_),
    .Q(\cpuregs[27] [15]),
    .QN(_27747_)
  );
  DFF_X1 cpuregs_reg_27__16_  (
    .CK(clk),
    .D(_01442_),
    .Q(\cpuregs[27] [16]),
    .QN(_27746_)
  );
  DFF_X1 cpuregs_reg_27__17_  (
    .CK(clk),
    .D(_01443_),
    .Q(\cpuregs[27] [17]),
    .QN(_27745_)
  );
  DFF_X1 cpuregs_reg_27__18_  (
    .CK(clk),
    .D(_01444_),
    .Q(\cpuregs[27] [18]),
    .QN(_27744_)
  );
  DFF_X1 cpuregs_reg_27__19_  (
    .CK(clk),
    .D(_01445_),
    .Q(\cpuregs[27] [19]),
    .QN(_27743_)
  );
  DFF_X1 cpuregs_reg_27__1_  (
    .CK(clk),
    .D(_01427_),
    .Q(\cpuregs[27] [1]),
    .QN(_27761_)
  );
  DFF_X1 cpuregs_reg_27__20_  (
    .CK(clk),
    .D(_01446_),
    .Q(\cpuregs[27] [20]),
    .QN(_27742_)
  );
  DFF_X1 cpuregs_reg_27__21_  (
    .CK(clk),
    .D(_01447_),
    .Q(\cpuregs[27] [21]),
    .QN(_27741_)
  );
  DFF_X1 cpuregs_reg_27__22_  (
    .CK(clk),
    .D(_01448_),
    .Q(\cpuregs[27] [22]),
    .QN(_27740_)
  );
  DFF_X1 cpuregs_reg_27__23_  (
    .CK(clk),
    .D(_01449_),
    .Q(\cpuregs[27] [23]),
    .QN(_27739_)
  );
  DFF_X1 cpuregs_reg_27__24_  (
    .CK(clk),
    .D(_01450_),
    .Q(\cpuregs[27] [24]),
    .QN(_27738_)
  );
  DFF_X1 cpuregs_reg_27__25_  (
    .CK(clk),
    .D(_01451_),
    .Q(\cpuregs[27] [25]),
    .QN(_27737_)
  );
  DFF_X1 cpuregs_reg_27__26_  (
    .CK(clk),
    .D(_01452_),
    .Q(\cpuregs[27] [26]),
    .QN(_27736_)
  );
  DFF_X1 cpuregs_reg_27__27_  (
    .CK(clk),
    .D(_01453_),
    .Q(\cpuregs[27] [27]),
    .QN(_27735_)
  );
  DFF_X1 cpuregs_reg_27__28_  (
    .CK(clk),
    .D(_01454_),
    .Q(\cpuregs[27] [28]),
    .QN(_27734_)
  );
  DFF_X1 cpuregs_reg_27__29_  (
    .CK(clk),
    .D(_01455_),
    .Q(\cpuregs[27] [29]),
    .QN(_27733_)
  );
  DFF_X1 cpuregs_reg_27__2_  (
    .CK(clk),
    .D(_01428_),
    .Q(\cpuregs[27] [2]),
    .QN(_27760_)
  );
  DFF_X1 cpuregs_reg_27__30_  (
    .CK(clk),
    .D(_01456_),
    .Q(\cpuregs[27] [30]),
    .QN(_27732_)
  );
  DFF_X1 cpuregs_reg_27__31_  (
    .CK(clk),
    .D(_00507_),
    .Q(\cpuregs[27] [31]),
    .QN(_28681_)
  );
  DFF_X1 cpuregs_reg_27__3_  (
    .CK(clk),
    .D(_01429_),
    .Q(\cpuregs[27] [3]),
    .QN(_27759_)
  );
  DFF_X1 cpuregs_reg_27__4_  (
    .CK(clk),
    .D(_01430_),
    .Q(\cpuregs[27] [4]),
    .QN(_27758_)
  );
  DFF_X1 cpuregs_reg_27__5_  (
    .CK(clk),
    .D(_01431_),
    .Q(\cpuregs[27] [5]),
    .QN(_27757_)
  );
  DFF_X1 cpuregs_reg_27__6_  (
    .CK(clk),
    .D(_01432_),
    .Q(\cpuregs[27] [6]),
    .QN(_27756_)
  );
  DFF_X1 cpuregs_reg_27__7_  (
    .CK(clk),
    .D(_01433_),
    .Q(\cpuregs[27] [7]),
    .QN(_27755_)
  );
  DFF_X1 cpuregs_reg_27__8_  (
    .CK(clk),
    .D(_01434_),
    .Q(\cpuregs[27] [8]),
    .QN(_27754_)
  );
  DFF_X1 cpuregs_reg_27__9_  (
    .CK(clk),
    .D(_01435_),
    .Q(\cpuregs[27] [9]),
    .QN(_27753_)
  );
  DFF_X1 cpuregs_reg_28__0_  (
    .CK(clk),
    .D(_01395_),
    .Q(\cpuregs[28] [0]),
    .QN(_27793_)
  );
  DFF_X1 cpuregs_reg_28__10_  (
    .CK(clk),
    .D(_01405_),
    .Q(\cpuregs[28] [10]),
    .QN(_27783_)
  );
  DFF_X1 cpuregs_reg_28__11_  (
    .CK(clk),
    .D(_01406_),
    .Q(\cpuregs[28] [11]),
    .QN(_27782_)
  );
  DFF_X1 cpuregs_reg_28__12_  (
    .CK(clk),
    .D(_01407_),
    .Q(\cpuregs[28] [12]),
    .QN(_27781_)
  );
  DFF_X1 cpuregs_reg_28__13_  (
    .CK(clk),
    .D(_01408_),
    .Q(\cpuregs[28] [13]),
    .QN(_27780_)
  );
  DFF_X1 cpuregs_reg_28__14_  (
    .CK(clk),
    .D(_01409_),
    .Q(\cpuregs[28] [14]),
    .QN(_27779_)
  );
  DFF_X1 cpuregs_reg_28__15_  (
    .CK(clk),
    .D(_01410_),
    .Q(\cpuregs[28] [15]),
    .QN(_27778_)
  );
  DFF_X1 cpuregs_reg_28__16_  (
    .CK(clk),
    .D(_01411_),
    .Q(\cpuregs[28] [16]),
    .QN(_27777_)
  );
  DFF_X1 cpuregs_reg_28__17_  (
    .CK(clk),
    .D(_01412_),
    .Q(\cpuregs[28] [17]),
    .QN(_27776_)
  );
  DFF_X1 cpuregs_reg_28__18_  (
    .CK(clk),
    .D(_01413_),
    .Q(\cpuregs[28] [18]),
    .QN(_27775_)
  );
  DFF_X1 cpuregs_reg_28__19_  (
    .CK(clk),
    .D(_01414_),
    .Q(\cpuregs[28] [19]),
    .QN(_27774_)
  );
  DFF_X1 cpuregs_reg_28__1_  (
    .CK(clk),
    .D(_01396_),
    .Q(\cpuregs[28] [1]),
    .QN(_27792_)
  );
  DFF_X1 cpuregs_reg_28__20_  (
    .CK(clk),
    .D(_01415_),
    .Q(\cpuregs[28] [20]),
    .QN(_27773_)
  );
  DFF_X1 cpuregs_reg_28__21_  (
    .CK(clk),
    .D(_01416_),
    .Q(\cpuregs[28] [21]),
    .QN(_27772_)
  );
  DFF_X1 cpuregs_reg_28__22_  (
    .CK(clk),
    .D(_01417_),
    .Q(\cpuregs[28] [22]),
    .QN(_27771_)
  );
  DFF_X1 cpuregs_reg_28__23_  (
    .CK(clk),
    .D(_01418_),
    .Q(\cpuregs[28] [23]),
    .QN(_27770_)
  );
  DFF_X1 cpuregs_reg_28__24_  (
    .CK(clk),
    .D(_01419_),
    .Q(\cpuregs[28] [24]),
    .QN(_27769_)
  );
  DFF_X1 cpuregs_reg_28__25_  (
    .CK(clk),
    .D(_01420_),
    .Q(\cpuregs[28] [25]),
    .QN(_27768_)
  );
  DFF_X1 cpuregs_reg_28__26_  (
    .CK(clk),
    .D(_01421_),
    .Q(\cpuregs[28] [26]),
    .QN(_27767_)
  );
  DFF_X1 cpuregs_reg_28__27_  (
    .CK(clk),
    .D(_01422_),
    .Q(\cpuregs[28] [27]),
    .QN(_27766_)
  );
  DFF_X1 cpuregs_reg_28__28_  (
    .CK(clk),
    .D(_01423_),
    .Q(\cpuregs[28] [28]),
    .QN(_27765_)
  );
  DFF_X1 cpuregs_reg_28__29_  (
    .CK(clk),
    .D(_01424_),
    .Q(\cpuregs[28] [29]),
    .QN(_27764_)
  );
  DFF_X1 cpuregs_reg_28__2_  (
    .CK(clk),
    .D(_01397_),
    .Q(\cpuregs[28] [2]),
    .QN(_27791_)
  );
  DFF_X1 cpuregs_reg_28__30_  (
    .CK(clk),
    .D(_01425_),
    .Q(\cpuregs[28] [30]),
    .QN(_27763_)
  );
  DFF_X1 cpuregs_reg_28__31_  (
    .CK(clk),
    .D(_00506_),
    .Q(\cpuregs[28] [31]),
    .QN(_28682_)
  );
  DFF_X1 cpuregs_reg_28__3_  (
    .CK(clk),
    .D(_01398_),
    .Q(\cpuregs[28] [3]),
    .QN(_27790_)
  );
  DFF_X1 cpuregs_reg_28__4_  (
    .CK(clk),
    .D(_01399_),
    .Q(\cpuregs[28] [4]),
    .QN(_27789_)
  );
  DFF_X1 cpuregs_reg_28__5_  (
    .CK(clk),
    .D(_01400_),
    .Q(\cpuregs[28] [5]),
    .QN(_27788_)
  );
  DFF_X1 cpuregs_reg_28__6_  (
    .CK(clk),
    .D(_01401_),
    .Q(\cpuregs[28] [6]),
    .QN(_27787_)
  );
  DFF_X1 cpuregs_reg_28__7_  (
    .CK(clk),
    .D(_01402_),
    .Q(\cpuregs[28] [7]),
    .QN(_27786_)
  );
  DFF_X1 cpuregs_reg_28__8_  (
    .CK(clk),
    .D(_01403_),
    .Q(\cpuregs[28] [8]),
    .QN(_27785_)
  );
  DFF_X1 cpuregs_reg_28__9_  (
    .CK(clk),
    .D(_01404_),
    .Q(\cpuregs[28] [9]),
    .QN(_27784_)
  );
  DFF_X1 cpuregs_reg_29__0_  (
    .CK(clk),
    .D(_01364_),
    .Q(\cpuregs[29] [0]),
    .QN(_27824_)
  );
  DFF_X1 cpuregs_reg_29__10_  (
    .CK(clk),
    .D(_01374_),
    .Q(\cpuregs[29] [10]),
    .QN(_27814_)
  );
  DFF_X1 cpuregs_reg_29__11_  (
    .CK(clk),
    .D(_01375_),
    .Q(\cpuregs[29] [11]),
    .QN(_27813_)
  );
  DFF_X1 cpuregs_reg_29__12_  (
    .CK(clk),
    .D(_01376_),
    .Q(\cpuregs[29] [12]),
    .QN(_27812_)
  );
  DFF_X1 cpuregs_reg_29__13_  (
    .CK(clk),
    .D(_01377_),
    .Q(\cpuregs[29] [13]),
    .QN(_27811_)
  );
  DFF_X1 cpuregs_reg_29__14_  (
    .CK(clk),
    .D(_01378_),
    .Q(\cpuregs[29] [14]),
    .QN(_27810_)
  );
  DFF_X1 cpuregs_reg_29__15_  (
    .CK(clk),
    .D(_01379_),
    .Q(\cpuregs[29] [15]),
    .QN(_27809_)
  );
  DFF_X1 cpuregs_reg_29__16_  (
    .CK(clk),
    .D(_01380_),
    .Q(\cpuregs[29] [16]),
    .QN(_27808_)
  );
  DFF_X1 cpuregs_reg_29__17_  (
    .CK(clk),
    .D(_01381_),
    .Q(\cpuregs[29] [17]),
    .QN(_27807_)
  );
  DFF_X1 cpuregs_reg_29__18_  (
    .CK(clk),
    .D(_01382_),
    .Q(\cpuregs[29] [18]),
    .QN(_27806_)
  );
  DFF_X1 cpuregs_reg_29__19_  (
    .CK(clk),
    .D(_01383_),
    .Q(\cpuregs[29] [19]),
    .QN(_27805_)
  );
  DFF_X1 cpuregs_reg_29__1_  (
    .CK(clk),
    .D(_01365_),
    .Q(\cpuregs[29] [1]),
    .QN(_27823_)
  );
  DFF_X1 cpuregs_reg_29__20_  (
    .CK(clk),
    .D(_01384_),
    .Q(\cpuregs[29] [20]),
    .QN(_27804_)
  );
  DFF_X1 cpuregs_reg_29__21_  (
    .CK(clk),
    .D(_01385_),
    .Q(\cpuregs[29] [21]),
    .QN(_27803_)
  );
  DFF_X1 cpuregs_reg_29__22_  (
    .CK(clk),
    .D(_01386_),
    .Q(\cpuregs[29] [22]),
    .QN(_27802_)
  );
  DFF_X1 cpuregs_reg_29__23_  (
    .CK(clk),
    .D(_01387_),
    .Q(\cpuregs[29] [23]),
    .QN(_27801_)
  );
  DFF_X1 cpuregs_reg_29__24_  (
    .CK(clk),
    .D(_01388_),
    .Q(\cpuregs[29] [24]),
    .QN(_27800_)
  );
  DFF_X1 cpuregs_reg_29__25_  (
    .CK(clk),
    .D(_01389_),
    .Q(\cpuregs[29] [25]),
    .QN(_27799_)
  );
  DFF_X1 cpuregs_reg_29__26_  (
    .CK(clk),
    .D(_01390_),
    .Q(\cpuregs[29] [26]),
    .QN(_27798_)
  );
  DFF_X1 cpuregs_reg_29__27_  (
    .CK(clk),
    .D(_01391_),
    .Q(\cpuregs[29] [27]),
    .QN(_27797_)
  );
  DFF_X1 cpuregs_reg_29__28_  (
    .CK(clk),
    .D(_01392_),
    .Q(\cpuregs[29] [28]),
    .QN(_27796_)
  );
  DFF_X1 cpuregs_reg_29__29_  (
    .CK(clk),
    .D(_01393_),
    .Q(\cpuregs[29] [29]),
    .QN(_27795_)
  );
  DFF_X1 cpuregs_reg_29__2_  (
    .CK(clk),
    .D(_01366_),
    .Q(\cpuregs[29] [2]),
    .QN(_27822_)
  );
  DFF_X1 cpuregs_reg_29__30_  (
    .CK(clk),
    .D(_01394_),
    .Q(\cpuregs[29] [30]),
    .QN(_27794_)
  );
  DFF_X1 cpuregs_reg_29__31_  (
    .CK(clk),
    .D(_00505_),
    .Q(\cpuregs[29] [31]),
    .QN(_28683_)
  );
  DFF_X1 cpuregs_reg_29__3_  (
    .CK(clk),
    .D(_01367_),
    .Q(\cpuregs[29] [3]),
    .QN(_27821_)
  );
  DFF_X1 cpuregs_reg_29__4_  (
    .CK(clk),
    .D(_01368_),
    .Q(\cpuregs[29] [4]),
    .QN(_27820_)
  );
  DFF_X1 cpuregs_reg_29__5_  (
    .CK(clk),
    .D(_01369_),
    .Q(\cpuregs[29] [5]),
    .QN(_27819_)
  );
  DFF_X1 cpuregs_reg_29__6_  (
    .CK(clk),
    .D(_01370_),
    .Q(\cpuregs[29] [6]),
    .QN(_27818_)
  );
  DFF_X1 cpuregs_reg_29__7_  (
    .CK(clk),
    .D(_01371_),
    .Q(\cpuregs[29] [7]),
    .QN(_27817_)
  );
  DFF_X1 cpuregs_reg_29__8_  (
    .CK(clk),
    .D(_01372_),
    .Q(\cpuregs[29] [8]),
    .QN(_27816_)
  );
  DFF_X1 cpuregs_reg_29__9_  (
    .CK(clk),
    .D(_01373_),
    .Q(\cpuregs[29] [9]),
    .QN(_27815_)
  );
  DFF_X1 cpuregs_reg_2__0_  (
    .CK(clk),
    .D(_00806_),
    .Q(\cpuregs[2] [0]),
    .QN(_28382_)
  );
  DFF_X1 cpuregs_reg_2__10_  (
    .CK(clk),
    .D(_00816_),
    .Q(\cpuregs[2] [10]),
    .QN(_28372_)
  );
  DFF_X1 cpuregs_reg_2__11_  (
    .CK(clk),
    .D(_00817_),
    .Q(\cpuregs[2] [11]),
    .QN(_28371_)
  );
  DFF_X1 cpuregs_reg_2__12_  (
    .CK(clk),
    .D(_00818_),
    .Q(\cpuregs[2] [12]),
    .QN(_28370_)
  );
  DFF_X1 cpuregs_reg_2__13_  (
    .CK(clk),
    .D(_00819_),
    .Q(\cpuregs[2] [13]),
    .QN(_28369_)
  );
  DFF_X1 cpuregs_reg_2__14_  (
    .CK(clk),
    .D(_00820_),
    .Q(\cpuregs[2] [14]),
    .QN(_28368_)
  );
  DFF_X1 cpuregs_reg_2__15_  (
    .CK(clk),
    .D(_00821_),
    .Q(\cpuregs[2] [15]),
    .QN(_28367_)
  );
  DFF_X1 cpuregs_reg_2__16_  (
    .CK(clk),
    .D(_00822_),
    .Q(\cpuregs[2] [16]),
    .QN(_28366_)
  );
  DFF_X1 cpuregs_reg_2__17_  (
    .CK(clk),
    .D(_00823_),
    .Q(\cpuregs[2] [17]),
    .QN(_28365_)
  );
  DFF_X1 cpuregs_reg_2__18_  (
    .CK(clk),
    .D(_00824_),
    .Q(\cpuregs[2] [18]),
    .QN(_28364_)
  );
  DFF_X1 cpuregs_reg_2__19_  (
    .CK(clk),
    .D(_00825_),
    .Q(\cpuregs[2] [19]),
    .QN(_28363_)
  );
  DFF_X1 cpuregs_reg_2__1_  (
    .CK(clk),
    .D(_00807_),
    .Q(\cpuregs[2] [1]),
    .QN(_28381_)
  );
  DFF_X1 cpuregs_reg_2__20_  (
    .CK(clk),
    .D(_00826_),
    .Q(\cpuregs[2] [20]),
    .QN(_28362_)
  );
  DFF_X1 cpuregs_reg_2__21_  (
    .CK(clk),
    .D(_00827_),
    .Q(\cpuregs[2] [21]),
    .QN(_28361_)
  );
  DFF_X1 cpuregs_reg_2__22_  (
    .CK(clk),
    .D(_00828_),
    .Q(\cpuregs[2] [22]),
    .QN(_28360_)
  );
  DFF_X1 cpuregs_reg_2__23_  (
    .CK(clk),
    .D(_00829_),
    .Q(\cpuregs[2] [23]),
    .QN(_28359_)
  );
  DFF_X1 cpuregs_reg_2__24_  (
    .CK(clk),
    .D(_00830_),
    .Q(\cpuregs[2] [24]),
    .QN(_28358_)
  );
  DFF_X1 cpuregs_reg_2__25_  (
    .CK(clk),
    .D(_00831_),
    .Q(\cpuregs[2] [25]),
    .QN(_28357_)
  );
  DFF_X1 cpuregs_reg_2__26_  (
    .CK(clk),
    .D(_00832_),
    .Q(\cpuregs[2] [26]),
    .QN(_28356_)
  );
  DFF_X1 cpuregs_reg_2__27_  (
    .CK(clk),
    .D(_00833_),
    .Q(\cpuregs[2] [27]),
    .QN(_28355_)
  );
  DFF_X1 cpuregs_reg_2__28_  (
    .CK(clk),
    .D(_00834_),
    .Q(\cpuregs[2] [28]),
    .QN(_28354_)
  );
  DFF_X1 cpuregs_reg_2__29_  (
    .CK(clk),
    .D(_00835_),
    .Q(\cpuregs[2] [29]),
    .QN(_28353_)
  );
  DFF_X1 cpuregs_reg_2__2_  (
    .CK(clk),
    .D(_00808_),
    .Q(\cpuregs[2] [2]),
    .QN(_28380_)
  );
  DFF_X1 cpuregs_reg_2__30_  (
    .CK(clk),
    .D(_00836_),
    .Q(\cpuregs[2] [30]),
    .QN(_28352_)
  );
  DFF_X1 cpuregs_reg_2__31_  (
    .CK(clk),
    .D(_00504_),
    .Q(\cpuregs[2] [31]),
    .QN(_28684_)
  );
  DFF_X1 cpuregs_reg_2__3_  (
    .CK(clk),
    .D(_00809_),
    .Q(\cpuregs[2] [3]),
    .QN(_28379_)
  );
  DFF_X1 cpuregs_reg_2__4_  (
    .CK(clk),
    .D(_00810_),
    .Q(\cpuregs[2] [4]),
    .QN(_28378_)
  );
  DFF_X1 cpuregs_reg_2__5_  (
    .CK(clk),
    .D(_00811_),
    .Q(\cpuregs[2] [5]),
    .QN(_28377_)
  );
  DFF_X1 cpuregs_reg_2__6_  (
    .CK(clk),
    .D(_00812_),
    .Q(\cpuregs[2] [6]),
    .QN(_28376_)
  );
  DFF_X1 cpuregs_reg_2__7_  (
    .CK(clk),
    .D(_00813_),
    .Q(\cpuregs[2] [7]),
    .QN(_28375_)
  );
  DFF_X1 cpuregs_reg_2__8_  (
    .CK(clk),
    .D(_00814_),
    .Q(\cpuregs[2] [8]),
    .QN(_28374_)
  );
  DFF_X1 cpuregs_reg_2__9_  (
    .CK(clk),
    .D(_00815_),
    .Q(\cpuregs[2] [9]),
    .QN(_28373_)
  );
  DFF_X1 cpuregs_reg_30__0_  (
    .CK(clk),
    .D(_01302_),
    .Q(\cpuregs[30] [0]),
    .QN(_27886_)
  );
  DFF_X1 cpuregs_reg_30__10_  (
    .CK(clk),
    .D(_01312_),
    .Q(\cpuregs[30] [10]),
    .QN(_27876_)
  );
  DFF_X1 cpuregs_reg_30__11_  (
    .CK(clk),
    .D(_01313_),
    .Q(\cpuregs[30] [11]),
    .QN(_27875_)
  );
  DFF_X1 cpuregs_reg_30__12_  (
    .CK(clk),
    .D(_01314_),
    .Q(\cpuregs[30] [12]),
    .QN(_27874_)
  );
  DFF_X1 cpuregs_reg_30__13_  (
    .CK(clk),
    .D(_01315_),
    .Q(\cpuregs[30] [13]),
    .QN(_27873_)
  );
  DFF_X1 cpuregs_reg_30__14_  (
    .CK(clk),
    .D(_01316_),
    .Q(\cpuregs[30] [14]),
    .QN(_27872_)
  );
  DFF_X1 cpuregs_reg_30__15_  (
    .CK(clk),
    .D(_01317_),
    .Q(\cpuregs[30] [15]),
    .QN(_27871_)
  );
  DFF_X1 cpuregs_reg_30__16_  (
    .CK(clk),
    .D(_01318_),
    .Q(\cpuregs[30] [16]),
    .QN(_27870_)
  );
  DFF_X1 cpuregs_reg_30__17_  (
    .CK(clk),
    .D(_01319_),
    .Q(\cpuregs[30] [17]),
    .QN(_27869_)
  );
  DFF_X1 cpuregs_reg_30__18_  (
    .CK(clk),
    .D(_01320_),
    .Q(\cpuregs[30] [18]),
    .QN(_27868_)
  );
  DFF_X1 cpuregs_reg_30__19_  (
    .CK(clk),
    .D(_01321_),
    .Q(\cpuregs[30] [19]),
    .QN(_27867_)
  );
  DFF_X1 cpuregs_reg_30__1_  (
    .CK(clk),
    .D(_01303_),
    .Q(\cpuregs[30] [1]),
    .QN(_27885_)
  );
  DFF_X1 cpuregs_reg_30__20_  (
    .CK(clk),
    .D(_01322_),
    .Q(\cpuregs[30] [20]),
    .QN(_27866_)
  );
  DFF_X1 cpuregs_reg_30__21_  (
    .CK(clk),
    .D(_01323_),
    .Q(\cpuregs[30] [21]),
    .QN(_27865_)
  );
  DFF_X1 cpuregs_reg_30__22_  (
    .CK(clk),
    .D(_01324_),
    .Q(\cpuregs[30] [22]),
    .QN(_27864_)
  );
  DFF_X1 cpuregs_reg_30__23_  (
    .CK(clk),
    .D(_01325_),
    .Q(\cpuregs[30] [23]),
    .QN(_27863_)
  );
  DFF_X1 cpuregs_reg_30__24_  (
    .CK(clk),
    .D(_01326_),
    .Q(\cpuregs[30] [24]),
    .QN(_27862_)
  );
  DFF_X1 cpuregs_reg_30__25_  (
    .CK(clk),
    .D(_01327_),
    .Q(\cpuregs[30] [25]),
    .QN(_27861_)
  );
  DFF_X1 cpuregs_reg_30__26_  (
    .CK(clk),
    .D(_01328_),
    .Q(\cpuregs[30] [26]),
    .QN(_27860_)
  );
  DFF_X1 cpuregs_reg_30__27_  (
    .CK(clk),
    .D(_01329_),
    .Q(\cpuregs[30] [27]),
    .QN(_27859_)
  );
  DFF_X1 cpuregs_reg_30__28_  (
    .CK(clk),
    .D(_01330_),
    .Q(\cpuregs[30] [28]),
    .QN(_27858_)
  );
  DFF_X1 cpuregs_reg_30__29_  (
    .CK(clk),
    .D(_01331_),
    .Q(\cpuregs[30] [29]),
    .QN(_27857_)
  );
  DFF_X1 cpuregs_reg_30__2_  (
    .CK(clk),
    .D(_01304_),
    .Q(\cpuregs[30] [2]),
    .QN(_27884_)
  );
  DFF_X1 cpuregs_reg_30__30_  (
    .CK(clk),
    .D(_01332_),
    .Q(\cpuregs[30] [30]),
    .QN(_27856_)
  );
  DFF_X1 cpuregs_reg_30__31_  (
    .CK(clk),
    .D(_00503_),
    .Q(\cpuregs[30] [31]),
    .QN(_28685_)
  );
  DFF_X1 cpuregs_reg_30__3_  (
    .CK(clk),
    .D(_01305_),
    .Q(\cpuregs[30] [3]),
    .QN(_27883_)
  );
  DFF_X1 cpuregs_reg_30__4_  (
    .CK(clk),
    .D(_01306_),
    .Q(\cpuregs[30] [4]),
    .QN(_27882_)
  );
  DFF_X1 cpuregs_reg_30__5_  (
    .CK(clk),
    .D(_01307_),
    .Q(\cpuregs[30] [5]),
    .QN(_27881_)
  );
  DFF_X1 cpuregs_reg_30__6_  (
    .CK(clk),
    .D(_01308_),
    .Q(\cpuregs[30] [6]),
    .QN(_27880_)
  );
  DFF_X1 cpuregs_reg_30__7_  (
    .CK(clk),
    .D(_01309_),
    .Q(\cpuregs[30] [7]),
    .QN(_27879_)
  );
  DFF_X1 cpuregs_reg_30__8_  (
    .CK(clk),
    .D(_01310_),
    .Q(\cpuregs[30] [8]),
    .QN(_27878_)
  );
  DFF_X1 cpuregs_reg_30__9_  (
    .CK(clk),
    .D(_01311_),
    .Q(\cpuregs[30] [9]),
    .QN(_27877_)
  );
  DFF_X1 cpuregs_reg_31__0_  (
    .CK(clk),
    .D(_01457_),
    .Q(\cpuregs[31] [0]),
    .QN(_27731_)
  );
  DFF_X1 cpuregs_reg_31__10_  (
    .CK(clk),
    .D(_01467_),
    .Q(\cpuregs[31] [10]),
    .QN(_27721_)
  );
  DFF_X1 cpuregs_reg_31__11_  (
    .CK(clk),
    .D(_01468_),
    .Q(\cpuregs[31] [11]),
    .QN(_27720_)
  );
  DFF_X1 cpuregs_reg_31__12_  (
    .CK(clk),
    .D(_01469_),
    .Q(\cpuregs[31] [12]),
    .QN(_27719_)
  );
  DFF_X1 cpuregs_reg_31__13_  (
    .CK(clk),
    .D(_01470_),
    .Q(\cpuregs[31] [13]),
    .QN(_27718_)
  );
  DFF_X1 cpuregs_reg_31__14_  (
    .CK(clk),
    .D(_01471_),
    .Q(\cpuregs[31] [14]),
    .QN(_27717_)
  );
  DFF_X1 cpuregs_reg_31__15_  (
    .CK(clk),
    .D(_01472_),
    .Q(\cpuregs[31] [15]),
    .QN(_27716_)
  );
  DFF_X1 cpuregs_reg_31__16_  (
    .CK(clk),
    .D(_01473_),
    .Q(\cpuregs[31] [16]),
    .QN(_27715_)
  );
  DFF_X1 cpuregs_reg_31__17_  (
    .CK(clk),
    .D(_01474_),
    .Q(\cpuregs[31] [17]),
    .QN(_27714_)
  );
  DFF_X1 cpuregs_reg_31__18_  (
    .CK(clk),
    .D(_01475_),
    .Q(\cpuregs[31] [18]),
    .QN(_27713_)
  );
  DFF_X1 cpuregs_reg_31__19_  (
    .CK(clk),
    .D(_01476_),
    .Q(\cpuregs[31] [19]),
    .QN(_27712_)
  );
  DFF_X1 cpuregs_reg_31__1_  (
    .CK(clk),
    .D(_01458_),
    .Q(\cpuregs[31] [1]),
    .QN(_27730_)
  );
  DFF_X1 cpuregs_reg_31__20_  (
    .CK(clk),
    .D(_01477_),
    .Q(\cpuregs[31] [20]),
    .QN(_27711_)
  );
  DFF_X1 cpuregs_reg_31__21_  (
    .CK(clk),
    .D(_01478_),
    .Q(\cpuregs[31] [21]),
    .QN(_27710_)
  );
  DFF_X1 cpuregs_reg_31__22_  (
    .CK(clk),
    .D(_01479_),
    .Q(\cpuregs[31] [22]),
    .QN(_27709_)
  );
  DFF_X1 cpuregs_reg_31__23_  (
    .CK(clk),
    .D(_01480_),
    .Q(\cpuregs[31] [23]),
    .QN(_27708_)
  );
  DFF_X1 cpuregs_reg_31__24_  (
    .CK(clk),
    .D(_01481_),
    .Q(\cpuregs[31] [24]),
    .QN(_27707_)
  );
  DFF_X1 cpuregs_reg_31__25_  (
    .CK(clk),
    .D(_01482_),
    .Q(\cpuregs[31] [25]),
    .QN(_27706_)
  );
  DFF_X1 cpuregs_reg_31__26_  (
    .CK(clk),
    .D(_01483_),
    .Q(\cpuregs[31] [26]),
    .QN(_27705_)
  );
  DFF_X1 cpuregs_reg_31__27_  (
    .CK(clk),
    .D(_01484_),
    .Q(\cpuregs[31] [27]),
    .QN(_27704_)
  );
  DFF_X1 cpuregs_reg_31__28_  (
    .CK(clk),
    .D(_01485_),
    .Q(\cpuregs[31] [28]),
    .QN(_27703_)
  );
  DFF_X1 cpuregs_reg_31__29_  (
    .CK(clk),
    .D(_01486_),
    .Q(\cpuregs[31] [29]),
    .QN(_27702_)
  );
  DFF_X1 cpuregs_reg_31__2_  (
    .CK(clk),
    .D(_01459_),
    .Q(\cpuregs[31] [2]),
    .QN(_27729_)
  );
  DFF_X1 cpuregs_reg_31__30_  (
    .CK(clk),
    .D(_01487_),
    .Q(\cpuregs[31] [30]),
    .QN(_27701_)
  );
  DFF_X1 cpuregs_reg_31__31_  (
    .CK(clk),
    .D(_00502_),
    .Q(\cpuregs[31] [31]),
    .QN(_28686_)
  );
  DFF_X1 cpuregs_reg_31__3_  (
    .CK(clk),
    .D(_01460_),
    .Q(\cpuregs[31] [3]),
    .QN(_27728_)
  );
  DFF_X1 cpuregs_reg_31__4_  (
    .CK(clk),
    .D(_01461_),
    .Q(\cpuregs[31] [4]),
    .QN(_27727_)
  );
  DFF_X1 cpuregs_reg_31__5_  (
    .CK(clk),
    .D(_01462_),
    .Q(\cpuregs[31] [5]),
    .QN(_27726_)
  );
  DFF_X1 cpuregs_reg_31__6_  (
    .CK(clk),
    .D(_01463_),
    .Q(\cpuregs[31] [6]),
    .QN(_27725_)
  );
  DFF_X1 cpuregs_reg_31__7_  (
    .CK(clk),
    .D(_01464_),
    .Q(\cpuregs[31] [7]),
    .QN(_27724_)
  );
  DFF_X1 cpuregs_reg_31__8_  (
    .CK(clk),
    .D(_01465_),
    .Q(\cpuregs[31] [8]),
    .QN(_27723_)
  );
  DFF_X1 cpuregs_reg_31__9_  (
    .CK(clk),
    .D(_01466_),
    .Q(\cpuregs[31] [9]),
    .QN(_27722_)
  );
  DFF_X1 cpuregs_reg_3__0_  (
    .CK(clk),
    .D(_00744_),
    .Q(\cpuregs[3] [0]),
    .QN(_28444_)
  );
  DFF_X1 cpuregs_reg_3__10_  (
    .CK(clk),
    .D(_00754_),
    .Q(\cpuregs[3] [10]),
    .QN(_28434_)
  );
  DFF_X1 cpuregs_reg_3__11_  (
    .CK(clk),
    .D(_00755_),
    .Q(\cpuregs[3] [11]),
    .QN(_28433_)
  );
  DFF_X1 cpuregs_reg_3__12_  (
    .CK(clk),
    .D(_00756_),
    .Q(\cpuregs[3] [12]),
    .QN(_28432_)
  );
  DFF_X1 cpuregs_reg_3__13_  (
    .CK(clk),
    .D(_00757_),
    .Q(\cpuregs[3] [13]),
    .QN(_28431_)
  );
  DFF_X1 cpuregs_reg_3__14_  (
    .CK(clk),
    .D(_00758_),
    .Q(\cpuregs[3] [14]),
    .QN(_28430_)
  );
  DFF_X1 cpuregs_reg_3__15_  (
    .CK(clk),
    .D(_00759_),
    .Q(\cpuregs[3] [15]),
    .QN(_28429_)
  );
  DFF_X1 cpuregs_reg_3__16_  (
    .CK(clk),
    .D(_00760_),
    .Q(\cpuregs[3] [16]),
    .QN(_28428_)
  );
  DFF_X1 cpuregs_reg_3__17_  (
    .CK(clk),
    .D(_00761_),
    .Q(\cpuregs[3] [17]),
    .QN(_28427_)
  );
  DFF_X1 cpuregs_reg_3__18_  (
    .CK(clk),
    .D(_00762_),
    .Q(\cpuregs[3] [18]),
    .QN(_28426_)
  );
  DFF_X1 cpuregs_reg_3__19_  (
    .CK(clk),
    .D(_00763_),
    .Q(\cpuregs[3] [19]),
    .QN(_28425_)
  );
  DFF_X1 cpuregs_reg_3__1_  (
    .CK(clk),
    .D(_00745_),
    .Q(\cpuregs[3] [1]),
    .QN(_28443_)
  );
  DFF_X1 cpuregs_reg_3__20_  (
    .CK(clk),
    .D(_00764_),
    .Q(\cpuregs[3] [20]),
    .QN(_28424_)
  );
  DFF_X1 cpuregs_reg_3__21_  (
    .CK(clk),
    .D(_00765_),
    .Q(\cpuregs[3] [21]),
    .QN(_28423_)
  );
  DFF_X1 cpuregs_reg_3__22_  (
    .CK(clk),
    .D(_00766_),
    .Q(\cpuregs[3] [22]),
    .QN(_28422_)
  );
  DFF_X1 cpuregs_reg_3__23_  (
    .CK(clk),
    .D(_00767_),
    .Q(\cpuregs[3] [23]),
    .QN(_28421_)
  );
  DFF_X1 cpuregs_reg_3__24_  (
    .CK(clk),
    .D(_00768_),
    .Q(\cpuregs[3] [24]),
    .QN(_28420_)
  );
  DFF_X1 cpuregs_reg_3__25_  (
    .CK(clk),
    .D(_00769_),
    .Q(\cpuregs[3] [25]),
    .QN(_28419_)
  );
  DFF_X1 cpuregs_reg_3__26_  (
    .CK(clk),
    .D(_00770_),
    .Q(\cpuregs[3] [26]),
    .QN(_28418_)
  );
  DFF_X1 cpuregs_reg_3__27_  (
    .CK(clk),
    .D(_00771_),
    .Q(\cpuregs[3] [27]),
    .QN(_28417_)
  );
  DFF_X1 cpuregs_reg_3__28_  (
    .CK(clk),
    .D(_00772_),
    .Q(\cpuregs[3] [28]),
    .QN(_28416_)
  );
  DFF_X1 cpuregs_reg_3__29_  (
    .CK(clk),
    .D(_00773_),
    .Q(\cpuregs[3] [29]),
    .QN(_28415_)
  );
  DFF_X1 cpuregs_reg_3__2_  (
    .CK(clk),
    .D(_00746_),
    .Q(\cpuregs[3] [2]),
    .QN(_28442_)
  );
  DFF_X1 cpuregs_reg_3__30_  (
    .CK(clk),
    .D(_00774_),
    .Q(\cpuregs[3] [30]),
    .QN(_28414_)
  );
  DFF_X1 cpuregs_reg_3__31_  (
    .CK(clk),
    .D(_00501_),
    .Q(\cpuregs[3] [31]),
    .QN(_28687_)
  );
  DFF_X1 cpuregs_reg_3__3_  (
    .CK(clk),
    .D(_00747_),
    .Q(\cpuregs[3] [3]),
    .QN(_28441_)
  );
  DFF_X1 cpuregs_reg_3__4_  (
    .CK(clk),
    .D(_00748_),
    .Q(\cpuregs[3] [4]),
    .QN(_28440_)
  );
  DFF_X1 cpuregs_reg_3__5_  (
    .CK(clk),
    .D(_00749_),
    .Q(\cpuregs[3] [5]),
    .QN(_28439_)
  );
  DFF_X1 cpuregs_reg_3__6_  (
    .CK(clk),
    .D(_00750_),
    .Q(\cpuregs[3] [6]),
    .QN(_28438_)
  );
  DFF_X1 cpuregs_reg_3__7_  (
    .CK(clk),
    .D(_00751_),
    .Q(\cpuregs[3] [7]),
    .QN(_28437_)
  );
  DFF_X1 cpuregs_reg_3__8_  (
    .CK(clk),
    .D(_00752_),
    .Q(\cpuregs[3] [8]),
    .QN(_28436_)
  );
  DFF_X1 cpuregs_reg_3__9_  (
    .CK(clk),
    .D(_00753_),
    .Q(\cpuregs[3] [9]),
    .QN(_28435_)
  );
  DFF_X1 cpuregs_reg_4__0_  (
    .CK(clk),
    .D(_01023_),
    .Q(\cpuregs[4] [0]),
    .QN(_28165_)
  );
  DFF_X1 cpuregs_reg_4__10_  (
    .CK(clk),
    .D(_01033_),
    .Q(\cpuregs[4] [10]),
    .QN(_28155_)
  );
  DFF_X1 cpuregs_reg_4__11_  (
    .CK(clk),
    .D(_01034_),
    .Q(\cpuregs[4] [11]),
    .QN(_28154_)
  );
  DFF_X1 cpuregs_reg_4__12_  (
    .CK(clk),
    .D(_01035_),
    .Q(\cpuregs[4] [12]),
    .QN(_28153_)
  );
  DFF_X1 cpuregs_reg_4__13_  (
    .CK(clk),
    .D(_01036_),
    .Q(\cpuregs[4] [13]),
    .QN(_28152_)
  );
  DFF_X1 cpuregs_reg_4__14_  (
    .CK(clk),
    .D(_01037_),
    .Q(\cpuregs[4] [14]),
    .QN(_28151_)
  );
  DFF_X1 cpuregs_reg_4__15_  (
    .CK(clk),
    .D(_01038_),
    .Q(\cpuregs[4] [15]),
    .QN(_28150_)
  );
  DFF_X1 cpuregs_reg_4__16_  (
    .CK(clk),
    .D(_01039_),
    .Q(\cpuregs[4] [16]),
    .QN(_28149_)
  );
  DFF_X1 cpuregs_reg_4__17_  (
    .CK(clk),
    .D(_01040_),
    .Q(\cpuregs[4] [17]),
    .QN(_28148_)
  );
  DFF_X1 cpuregs_reg_4__18_  (
    .CK(clk),
    .D(_01041_),
    .Q(\cpuregs[4] [18]),
    .QN(_28147_)
  );
  DFF_X1 cpuregs_reg_4__19_  (
    .CK(clk),
    .D(_01042_),
    .Q(\cpuregs[4] [19]),
    .QN(_28146_)
  );
  DFF_X1 cpuregs_reg_4__1_  (
    .CK(clk),
    .D(_01024_),
    .Q(\cpuregs[4] [1]),
    .QN(_28164_)
  );
  DFF_X1 cpuregs_reg_4__20_  (
    .CK(clk),
    .D(_01043_),
    .Q(\cpuregs[4] [20]),
    .QN(_28145_)
  );
  DFF_X1 cpuregs_reg_4__21_  (
    .CK(clk),
    .D(_01044_),
    .Q(\cpuregs[4] [21]),
    .QN(_28144_)
  );
  DFF_X1 cpuregs_reg_4__22_  (
    .CK(clk),
    .D(_01045_),
    .Q(\cpuregs[4] [22]),
    .QN(_28143_)
  );
  DFF_X1 cpuregs_reg_4__23_  (
    .CK(clk),
    .D(_01046_),
    .Q(\cpuregs[4] [23]),
    .QN(_28142_)
  );
  DFF_X1 cpuregs_reg_4__24_  (
    .CK(clk),
    .D(_01047_),
    .Q(\cpuregs[4] [24]),
    .QN(_28141_)
  );
  DFF_X1 cpuregs_reg_4__25_  (
    .CK(clk),
    .D(_01048_),
    .Q(\cpuregs[4] [25]),
    .QN(_28140_)
  );
  DFF_X1 cpuregs_reg_4__26_  (
    .CK(clk),
    .D(_01049_),
    .Q(\cpuregs[4] [26]),
    .QN(_28139_)
  );
  DFF_X1 cpuregs_reg_4__27_  (
    .CK(clk),
    .D(_01050_),
    .Q(\cpuregs[4] [27]),
    .QN(_28138_)
  );
  DFF_X1 cpuregs_reg_4__28_  (
    .CK(clk),
    .D(_01051_),
    .Q(\cpuregs[4] [28]),
    .QN(_28137_)
  );
  DFF_X1 cpuregs_reg_4__29_  (
    .CK(clk),
    .D(_01052_),
    .Q(\cpuregs[4] [29]),
    .QN(_28136_)
  );
  DFF_X1 cpuregs_reg_4__2_  (
    .CK(clk),
    .D(_01025_),
    .Q(\cpuregs[4] [2]),
    .QN(_28163_)
  );
  DFF_X1 cpuregs_reg_4__30_  (
    .CK(clk),
    .D(_01053_),
    .Q(\cpuregs[4] [30]),
    .QN(_28135_)
  );
  DFF_X1 cpuregs_reg_4__31_  (
    .CK(clk),
    .D(_00500_),
    .Q(\cpuregs[4] [31]),
    .QN(_28688_)
  );
  DFF_X1 cpuregs_reg_4__3_  (
    .CK(clk),
    .D(_01026_),
    .Q(\cpuregs[4] [3]),
    .QN(_28162_)
  );
  DFF_X1 cpuregs_reg_4__4_  (
    .CK(clk),
    .D(_01027_),
    .Q(\cpuregs[4] [4]),
    .QN(_28161_)
  );
  DFF_X1 cpuregs_reg_4__5_  (
    .CK(clk),
    .D(_01028_),
    .Q(\cpuregs[4] [5]),
    .QN(_28160_)
  );
  DFF_X1 cpuregs_reg_4__6_  (
    .CK(clk),
    .D(_01029_),
    .Q(\cpuregs[4] [6]),
    .QN(_28159_)
  );
  DFF_X1 cpuregs_reg_4__7_  (
    .CK(clk),
    .D(_01030_),
    .Q(\cpuregs[4] [7]),
    .QN(_28158_)
  );
  DFF_X1 cpuregs_reg_4__8_  (
    .CK(clk),
    .D(_01031_),
    .Q(\cpuregs[4] [8]),
    .QN(_28157_)
  );
  DFF_X1 cpuregs_reg_4__9_  (
    .CK(clk),
    .D(_01032_),
    .Q(\cpuregs[4] [9]),
    .QN(_28156_)
  );
  DFF_X1 cpuregs_reg_5__0_  (
    .CK(clk),
    .D(_01147_),
    .Q(\cpuregs[5] [0]),
    .QN(_28041_)
  );
  DFF_X1 cpuregs_reg_5__10_  (
    .CK(clk),
    .D(_01157_),
    .Q(\cpuregs[5] [10]),
    .QN(_28031_)
  );
  DFF_X1 cpuregs_reg_5__11_  (
    .CK(clk),
    .D(_01158_),
    .Q(\cpuregs[5] [11]),
    .QN(_28030_)
  );
  DFF_X1 cpuregs_reg_5__12_  (
    .CK(clk),
    .D(_01159_),
    .Q(\cpuregs[5] [12]),
    .QN(_28029_)
  );
  DFF_X1 cpuregs_reg_5__13_  (
    .CK(clk),
    .D(_01160_),
    .Q(\cpuregs[5] [13]),
    .QN(_28028_)
  );
  DFF_X1 cpuregs_reg_5__14_  (
    .CK(clk),
    .D(_01161_),
    .Q(\cpuregs[5] [14]),
    .QN(_28027_)
  );
  DFF_X1 cpuregs_reg_5__15_  (
    .CK(clk),
    .D(_01162_),
    .Q(\cpuregs[5] [15]),
    .QN(_28026_)
  );
  DFF_X1 cpuregs_reg_5__16_  (
    .CK(clk),
    .D(_01163_),
    .Q(\cpuregs[5] [16]),
    .QN(_28025_)
  );
  DFF_X1 cpuregs_reg_5__17_  (
    .CK(clk),
    .D(_01164_),
    .Q(\cpuregs[5] [17]),
    .QN(_28024_)
  );
  DFF_X1 cpuregs_reg_5__18_  (
    .CK(clk),
    .D(_01165_),
    .Q(\cpuregs[5] [18]),
    .QN(_28023_)
  );
  DFF_X1 cpuregs_reg_5__19_  (
    .CK(clk),
    .D(_01166_),
    .Q(\cpuregs[5] [19]),
    .QN(_28022_)
  );
  DFF_X1 cpuregs_reg_5__1_  (
    .CK(clk),
    .D(_01148_),
    .Q(\cpuregs[5] [1]),
    .QN(_28040_)
  );
  DFF_X1 cpuregs_reg_5__20_  (
    .CK(clk),
    .D(_01167_),
    .Q(\cpuregs[5] [20]),
    .QN(_28021_)
  );
  DFF_X1 cpuregs_reg_5__21_  (
    .CK(clk),
    .D(_01168_),
    .Q(\cpuregs[5] [21]),
    .QN(_28020_)
  );
  DFF_X1 cpuregs_reg_5__22_  (
    .CK(clk),
    .D(_01169_),
    .Q(\cpuregs[5] [22]),
    .QN(_28019_)
  );
  DFF_X1 cpuregs_reg_5__23_  (
    .CK(clk),
    .D(_01170_),
    .Q(\cpuregs[5] [23]),
    .QN(_28018_)
  );
  DFF_X1 cpuregs_reg_5__24_  (
    .CK(clk),
    .D(_01171_),
    .Q(\cpuregs[5] [24]),
    .QN(_28017_)
  );
  DFF_X1 cpuregs_reg_5__25_  (
    .CK(clk),
    .D(_01172_),
    .Q(\cpuregs[5] [25]),
    .QN(_28016_)
  );
  DFF_X1 cpuregs_reg_5__26_  (
    .CK(clk),
    .D(_01173_),
    .Q(\cpuregs[5] [26]),
    .QN(_28015_)
  );
  DFF_X1 cpuregs_reg_5__27_  (
    .CK(clk),
    .D(_01174_),
    .Q(\cpuregs[5] [27]),
    .QN(_28014_)
  );
  DFF_X1 cpuregs_reg_5__28_  (
    .CK(clk),
    .D(_01175_),
    .Q(\cpuregs[5] [28]),
    .QN(_28013_)
  );
  DFF_X1 cpuregs_reg_5__29_  (
    .CK(clk),
    .D(_01176_),
    .Q(\cpuregs[5] [29]),
    .QN(_28012_)
  );
  DFF_X1 cpuregs_reg_5__2_  (
    .CK(clk),
    .D(_01149_),
    .Q(\cpuregs[5] [2]),
    .QN(_28039_)
  );
  DFF_X1 cpuregs_reg_5__30_  (
    .CK(clk),
    .D(_01177_),
    .Q(\cpuregs[5] [30]),
    .QN(_28011_)
  );
  DFF_X1 cpuregs_reg_5__31_  (
    .CK(clk),
    .D(_00499_),
    .Q(\cpuregs[5] [31]),
    .QN(_28689_)
  );
  DFF_X1 cpuregs_reg_5__3_  (
    .CK(clk),
    .D(_01150_),
    .Q(\cpuregs[5] [3]),
    .QN(_28038_)
  );
  DFF_X1 cpuregs_reg_5__4_  (
    .CK(clk),
    .D(_01151_),
    .Q(\cpuregs[5] [4]),
    .QN(_28037_)
  );
  DFF_X1 cpuregs_reg_5__5_  (
    .CK(clk),
    .D(_01152_),
    .Q(\cpuregs[5] [5]),
    .QN(_28036_)
  );
  DFF_X1 cpuregs_reg_5__6_  (
    .CK(clk),
    .D(_01153_),
    .Q(\cpuregs[5] [6]),
    .QN(_28035_)
  );
  DFF_X1 cpuregs_reg_5__7_  (
    .CK(clk),
    .D(_01154_),
    .Q(\cpuregs[5] [7]),
    .QN(_28034_)
  );
  DFF_X1 cpuregs_reg_5__8_  (
    .CK(clk),
    .D(_01155_),
    .Q(\cpuregs[5] [8]),
    .QN(_28033_)
  );
  DFF_X1 cpuregs_reg_5__9_  (
    .CK(clk),
    .D(_01156_),
    .Q(\cpuregs[5] [9]),
    .QN(_28032_)
  );
  DFF_X1 cpuregs_reg_6__0_  (
    .CK(clk),
    .D(_01240_),
    .Q(\cpuregs[6] [0]),
    .QN(_27948_)
  );
  DFF_X1 cpuregs_reg_6__10_  (
    .CK(clk),
    .D(_01250_),
    .Q(\cpuregs[6] [10]),
    .QN(_27938_)
  );
  DFF_X1 cpuregs_reg_6__11_  (
    .CK(clk),
    .D(_01251_),
    .Q(\cpuregs[6] [11]),
    .QN(_27937_)
  );
  DFF_X1 cpuregs_reg_6__12_  (
    .CK(clk),
    .D(_01252_),
    .Q(\cpuregs[6] [12]),
    .QN(_27936_)
  );
  DFF_X1 cpuregs_reg_6__13_  (
    .CK(clk),
    .D(_01253_),
    .Q(\cpuregs[6] [13]),
    .QN(_27935_)
  );
  DFF_X1 cpuregs_reg_6__14_  (
    .CK(clk),
    .D(_01254_),
    .Q(\cpuregs[6] [14]),
    .QN(_27934_)
  );
  DFF_X1 cpuregs_reg_6__15_  (
    .CK(clk),
    .D(_01255_),
    .Q(\cpuregs[6] [15]),
    .QN(_27933_)
  );
  DFF_X1 cpuregs_reg_6__16_  (
    .CK(clk),
    .D(_01256_),
    .Q(\cpuregs[6] [16]),
    .QN(_27932_)
  );
  DFF_X1 cpuregs_reg_6__17_  (
    .CK(clk),
    .D(_01257_),
    .Q(\cpuregs[6] [17]),
    .QN(_27931_)
  );
  DFF_X1 cpuregs_reg_6__18_  (
    .CK(clk),
    .D(_01258_),
    .Q(\cpuregs[6] [18]),
    .QN(_27930_)
  );
  DFF_X1 cpuregs_reg_6__19_  (
    .CK(clk),
    .D(_01259_),
    .Q(\cpuregs[6] [19]),
    .QN(_27929_)
  );
  DFF_X1 cpuregs_reg_6__1_  (
    .CK(clk),
    .D(_01241_),
    .Q(\cpuregs[6] [1]),
    .QN(_27947_)
  );
  DFF_X1 cpuregs_reg_6__20_  (
    .CK(clk),
    .D(_01260_),
    .Q(\cpuregs[6] [20]),
    .QN(_27928_)
  );
  DFF_X1 cpuregs_reg_6__21_  (
    .CK(clk),
    .D(_01261_),
    .Q(\cpuregs[6] [21]),
    .QN(_27927_)
  );
  DFF_X1 cpuregs_reg_6__22_  (
    .CK(clk),
    .D(_01262_),
    .Q(\cpuregs[6] [22]),
    .QN(_27926_)
  );
  DFF_X1 cpuregs_reg_6__23_  (
    .CK(clk),
    .D(_01263_),
    .Q(\cpuregs[6] [23]),
    .QN(_27925_)
  );
  DFF_X1 cpuregs_reg_6__24_  (
    .CK(clk),
    .D(_01264_),
    .Q(\cpuregs[6] [24]),
    .QN(_27924_)
  );
  DFF_X1 cpuregs_reg_6__25_  (
    .CK(clk),
    .D(_01265_),
    .Q(\cpuregs[6] [25]),
    .QN(_27923_)
  );
  DFF_X1 cpuregs_reg_6__26_  (
    .CK(clk),
    .D(_01266_),
    .Q(\cpuregs[6] [26]),
    .QN(_27922_)
  );
  DFF_X1 cpuregs_reg_6__27_  (
    .CK(clk),
    .D(_01267_),
    .Q(\cpuregs[6] [27]),
    .QN(_27921_)
  );
  DFF_X1 cpuregs_reg_6__28_  (
    .CK(clk),
    .D(_01268_),
    .Q(\cpuregs[6] [28]),
    .QN(_27920_)
  );
  DFF_X1 cpuregs_reg_6__29_  (
    .CK(clk),
    .D(_01269_),
    .Q(\cpuregs[6] [29]),
    .QN(_27919_)
  );
  DFF_X1 cpuregs_reg_6__2_  (
    .CK(clk),
    .D(_01242_),
    .Q(\cpuregs[6] [2]),
    .QN(_27946_)
  );
  DFF_X1 cpuregs_reg_6__30_  (
    .CK(clk),
    .D(_01270_),
    .Q(\cpuregs[6] [30]),
    .QN(_27918_)
  );
  DFF_X1 cpuregs_reg_6__31_  (
    .CK(clk),
    .D(_00498_),
    .Q(\cpuregs[6] [31]),
    .QN(_28690_)
  );
  DFF_X1 cpuregs_reg_6__3_  (
    .CK(clk),
    .D(_01243_),
    .Q(\cpuregs[6] [3]),
    .QN(_27945_)
  );
  DFF_X1 cpuregs_reg_6__4_  (
    .CK(clk),
    .D(_01244_),
    .Q(\cpuregs[6] [4]),
    .QN(_27944_)
  );
  DFF_X1 cpuregs_reg_6__5_  (
    .CK(clk),
    .D(_01245_),
    .Q(\cpuregs[6] [5]),
    .QN(_27943_)
  );
  DFF_X1 cpuregs_reg_6__6_  (
    .CK(clk),
    .D(_01246_),
    .Q(\cpuregs[6] [6]),
    .QN(_27942_)
  );
  DFF_X1 cpuregs_reg_6__7_  (
    .CK(clk),
    .D(_01247_),
    .Q(\cpuregs[6] [7]),
    .QN(_27941_)
  );
  DFF_X1 cpuregs_reg_6__8_  (
    .CK(clk),
    .D(_01248_),
    .Q(\cpuregs[6] [8]),
    .QN(_27940_)
  );
  DFF_X1 cpuregs_reg_6__9_  (
    .CK(clk),
    .D(_01249_),
    .Q(\cpuregs[6] [9]),
    .QN(_27939_)
  );
  DFF_X1 cpuregs_reg_7__0_  (
    .CK(clk),
    .D(_01209_),
    .Q(\cpuregs[7] [0]),
    .QN(_27979_)
  );
  DFF_X1 cpuregs_reg_7__10_  (
    .CK(clk),
    .D(_01219_),
    .Q(\cpuregs[7] [10]),
    .QN(_27969_)
  );
  DFF_X1 cpuregs_reg_7__11_  (
    .CK(clk),
    .D(_01220_),
    .Q(\cpuregs[7] [11]),
    .QN(_27968_)
  );
  DFF_X1 cpuregs_reg_7__12_  (
    .CK(clk),
    .D(_01221_),
    .Q(\cpuregs[7] [12]),
    .QN(_27967_)
  );
  DFF_X1 cpuregs_reg_7__13_  (
    .CK(clk),
    .D(_01222_),
    .Q(\cpuregs[7] [13]),
    .QN(_27966_)
  );
  DFF_X1 cpuregs_reg_7__14_  (
    .CK(clk),
    .D(_01223_),
    .Q(\cpuregs[7] [14]),
    .QN(_27965_)
  );
  DFF_X1 cpuregs_reg_7__15_  (
    .CK(clk),
    .D(_01224_),
    .Q(\cpuregs[7] [15]),
    .QN(_27964_)
  );
  DFF_X1 cpuregs_reg_7__16_  (
    .CK(clk),
    .D(_01225_),
    .Q(\cpuregs[7] [16]),
    .QN(_27963_)
  );
  DFF_X1 cpuregs_reg_7__17_  (
    .CK(clk),
    .D(_01226_),
    .Q(\cpuregs[7] [17]),
    .QN(_27962_)
  );
  DFF_X1 cpuregs_reg_7__18_  (
    .CK(clk),
    .D(_01227_),
    .Q(\cpuregs[7] [18]),
    .QN(_27961_)
  );
  DFF_X1 cpuregs_reg_7__19_  (
    .CK(clk),
    .D(_01228_),
    .Q(\cpuregs[7] [19]),
    .QN(_27960_)
  );
  DFF_X1 cpuregs_reg_7__1_  (
    .CK(clk),
    .D(_01210_),
    .Q(\cpuregs[7] [1]),
    .QN(_27978_)
  );
  DFF_X1 cpuregs_reg_7__20_  (
    .CK(clk),
    .D(_01229_),
    .Q(\cpuregs[7] [20]),
    .QN(_27959_)
  );
  DFF_X1 cpuregs_reg_7__21_  (
    .CK(clk),
    .D(_01230_),
    .Q(\cpuregs[7] [21]),
    .QN(_27958_)
  );
  DFF_X1 cpuregs_reg_7__22_  (
    .CK(clk),
    .D(_01231_),
    .Q(\cpuregs[7] [22]),
    .QN(_27957_)
  );
  DFF_X1 cpuregs_reg_7__23_  (
    .CK(clk),
    .D(_01232_),
    .Q(\cpuregs[7] [23]),
    .QN(_27956_)
  );
  DFF_X1 cpuregs_reg_7__24_  (
    .CK(clk),
    .D(_01233_),
    .Q(\cpuregs[7] [24]),
    .QN(_27955_)
  );
  DFF_X1 cpuregs_reg_7__25_  (
    .CK(clk),
    .D(_01234_),
    .Q(\cpuregs[7] [25]),
    .QN(_27954_)
  );
  DFF_X1 cpuregs_reg_7__26_  (
    .CK(clk),
    .D(_01235_),
    .Q(\cpuregs[7] [26]),
    .QN(_27953_)
  );
  DFF_X1 cpuregs_reg_7__27_  (
    .CK(clk),
    .D(_01236_),
    .Q(\cpuregs[7] [27]),
    .QN(_27952_)
  );
  DFF_X1 cpuregs_reg_7__28_  (
    .CK(clk),
    .D(_01237_),
    .Q(\cpuregs[7] [28]),
    .QN(_27951_)
  );
  DFF_X1 cpuregs_reg_7__29_  (
    .CK(clk),
    .D(_01238_),
    .Q(\cpuregs[7] [29]),
    .QN(_27950_)
  );
  DFF_X1 cpuregs_reg_7__2_  (
    .CK(clk),
    .D(_01211_),
    .Q(\cpuregs[7] [2]),
    .QN(_27977_)
  );
  DFF_X1 cpuregs_reg_7__30_  (
    .CK(clk),
    .D(_01239_),
    .Q(\cpuregs[7] [30]),
    .QN(_27949_)
  );
  DFF_X1 cpuregs_reg_7__31_  (
    .CK(clk),
    .D(_00497_),
    .Q(\cpuregs[7] [31]),
    .QN(_28691_)
  );
  DFF_X1 cpuregs_reg_7__3_  (
    .CK(clk),
    .D(_01212_),
    .Q(\cpuregs[7] [3]),
    .QN(_27976_)
  );
  DFF_X1 cpuregs_reg_7__4_  (
    .CK(clk),
    .D(_01213_),
    .Q(\cpuregs[7] [4]),
    .QN(_27975_)
  );
  DFF_X1 cpuregs_reg_7__5_  (
    .CK(clk),
    .D(_01214_),
    .Q(\cpuregs[7] [5]),
    .QN(_27974_)
  );
  DFF_X1 cpuregs_reg_7__6_  (
    .CK(clk),
    .D(_01215_),
    .Q(\cpuregs[7] [6]),
    .QN(_27973_)
  );
  DFF_X1 cpuregs_reg_7__7_  (
    .CK(clk),
    .D(_01216_),
    .Q(\cpuregs[7] [7]),
    .QN(_27972_)
  );
  DFF_X1 cpuregs_reg_7__8_  (
    .CK(clk),
    .D(_01217_),
    .Q(\cpuregs[7] [8]),
    .QN(_27971_)
  );
  DFF_X1 cpuregs_reg_7__9_  (
    .CK(clk),
    .D(_01218_),
    .Q(\cpuregs[7] [9]),
    .QN(_27970_)
  );
  DFF_X1 cpuregs_reg_8__0_  (
    .CK(clk),
    .D(_01116_),
    .Q(\cpuregs[8] [0]),
    .QN(_28072_)
  );
  DFF_X1 cpuregs_reg_8__10_  (
    .CK(clk),
    .D(_01126_),
    .Q(\cpuregs[8] [10]),
    .QN(_28062_)
  );
  DFF_X1 cpuregs_reg_8__11_  (
    .CK(clk),
    .D(_01127_),
    .Q(\cpuregs[8] [11]),
    .QN(_28061_)
  );
  DFF_X1 cpuregs_reg_8__12_  (
    .CK(clk),
    .D(_01128_),
    .Q(\cpuregs[8] [12]),
    .QN(_28060_)
  );
  DFF_X1 cpuregs_reg_8__13_  (
    .CK(clk),
    .D(_01129_),
    .Q(\cpuregs[8] [13]),
    .QN(_28059_)
  );
  DFF_X1 cpuregs_reg_8__14_  (
    .CK(clk),
    .D(_01130_),
    .Q(\cpuregs[8] [14]),
    .QN(_28058_)
  );
  DFF_X1 cpuregs_reg_8__15_  (
    .CK(clk),
    .D(_01131_),
    .Q(\cpuregs[8] [15]),
    .QN(_28057_)
  );
  DFF_X1 cpuregs_reg_8__16_  (
    .CK(clk),
    .D(_01132_),
    .Q(\cpuregs[8] [16]),
    .QN(_28056_)
  );
  DFF_X1 cpuregs_reg_8__17_  (
    .CK(clk),
    .D(_01133_),
    .Q(\cpuregs[8] [17]),
    .QN(_28055_)
  );
  DFF_X1 cpuregs_reg_8__18_  (
    .CK(clk),
    .D(_01134_),
    .Q(\cpuregs[8] [18]),
    .QN(_28054_)
  );
  DFF_X1 cpuregs_reg_8__19_  (
    .CK(clk),
    .D(_01135_),
    .Q(\cpuregs[8] [19]),
    .QN(_28053_)
  );
  DFF_X1 cpuregs_reg_8__1_  (
    .CK(clk),
    .D(_01117_),
    .Q(\cpuregs[8] [1]),
    .QN(_28071_)
  );
  DFF_X1 cpuregs_reg_8__20_  (
    .CK(clk),
    .D(_01136_),
    .Q(\cpuregs[8] [20]),
    .QN(_28052_)
  );
  DFF_X1 cpuregs_reg_8__21_  (
    .CK(clk),
    .D(_01137_),
    .Q(\cpuregs[8] [21]),
    .QN(_28051_)
  );
  DFF_X1 cpuregs_reg_8__22_  (
    .CK(clk),
    .D(_01138_),
    .Q(\cpuregs[8] [22]),
    .QN(_28050_)
  );
  DFF_X1 cpuregs_reg_8__23_  (
    .CK(clk),
    .D(_01139_),
    .Q(\cpuregs[8] [23]),
    .QN(_28049_)
  );
  DFF_X1 cpuregs_reg_8__24_  (
    .CK(clk),
    .D(_01140_),
    .Q(\cpuregs[8] [24]),
    .QN(_28048_)
  );
  DFF_X1 cpuregs_reg_8__25_  (
    .CK(clk),
    .D(_01141_),
    .Q(\cpuregs[8] [25]),
    .QN(_28047_)
  );
  DFF_X1 cpuregs_reg_8__26_  (
    .CK(clk),
    .D(_01142_),
    .Q(\cpuregs[8] [26]),
    .QN(_28046_)
  );
  DFF_X1 cpuregs_reg_8__27_  (
    .CK(clk),
    .D(_01143_),
    .Q(\cpuregs[8] [27]),
    .QN(_28045_)
  );
  DFF_X1 cpuregs_reg_8__28_  (
    .CK(clk),
    .D(_01144_),
    .Q(\cpuregs[8] [28]),
    .QN(_28044_)
  );
  DFF_X1 cpuregs_reg_8__29_  (
    .CK(clk),
    .D(_01145_),
    .Q(\cpuregs[8] [29]),
    .QN(_28043_)
  );
  DFF_X1 cpuregs_reg_8__2_  (
    .CK(clk),
    .D(_01118_),
    .Q(\cpuregs[8] [2]),
    .QN(_28070_)
  );
  DFF_X1 cpuregs_reg_8__30_  (
    .CK(clk),
    .D(_01146_),
    .Q(\cpuregs[8] [30]),
    .QN(_28042_)
  );
  DFF_X1 cpuregs_reg_8__31_  (
    .CK(clk),
    .D(_00496_),
    .Q(\cpuregs[8] [31]),
    .QN(_28692_)
  );
  DFF_X1 cpuregs_reg_8__3_  (
    .CK(clk),
    .D(_01119_),
    .Q(\cpuregs[8] [3]),
    .QN(_28069_)
  );
  DFF_X1 cpuregs_reg_8__4_  (
    .CK(clk),
    .D(_01120_),
    .Q(\cpuregs[8] [4]),
    .QN(_28068_)
  );
  DFF_X1 cpuregs_reg_8__5_  (
    .CK(clk),
    .D(_01121_),
    .Q(\cpuregs[8] [5]),
    .QN(_28067_)
  );
  DFF_X1 cpuregs_reg_8__6_  (
    .CK(clk),
    .D(_01122_),
    .Q(\cpuregs[8] [6]),
    .QN(_28066_)
  );
  DFF_X1 cpuregs_reg_8__7_  (
    .CK(clk),
    .D(_01123_),
    .Q(\cpuregs[8] [7]),
    .QN(_28065_)
  );
  DFF_X1 cpuregs_reg_8__8_  (
    .CK(clk),
    .D(_01124_),
    .Q(\cpuregs[8] [8]),
    .QN(_28064_)
  );
  DFF_X1 cpuregs_reg_8__9_  (
    .CK(clk),
    .D(_01125_),
    .Q(\cpuregs[8] [9]),
    .QN(_28063_)
  );
  DFF_X1 cpuregs_reg_9__0_  (
    .CK(clk),
    .D(_01085_),
    .Q(\cpuregs[9] [0]),
    .QN(_28103_)
  );
  DFF_X1 cpuregs_reg_9__10_  (
    .CK(clk),
    .D(_01095_),
    .Q(\cpuregs[9] [10]),
    .QN(_28093_)
  );
  DFF_X1 cpuregs_reg_9__11_  (
    .CK(clk),
    .D(_01096_),
    .Q(\cpuregs[9] [11]),
    .QN(_28092_)
  );
  DFF_X1 cpuregs_reg_9__12_  (
    .CK(clk),
    .D(_01097_),
    .Q(\cpuregs[9] [12]),
    .QN(_28091_)
  );
  DFF_X1 cpuregs_reg_9__13_  (
    .CK(clk),
    .D(_01098_),
    .Q(\cpuregs[9] [13]),
    .QN(_28090_)
  );
  DFF_X1 cpuregs_reg_9__14_  (
    .CK(clk),
    .D(_01099_),
    .Q(\cpuregs[9] [14]),
    .QN(_28089_)
  );
  DFF_X1 cpuregs_reg_9__15_  (
    .CK(clk),
    .D(_01100_),
    .Q(\cpuregs[9] [15]),
    .QN(_28088_)
  );
  DFF_X1 cpuregs_reg_9__16_  (
    .CK(clk),
    .D(_01101_),
    .Q(\cpuregs[9] [16]),
    .QN(_28087_)
  );
  DFF_X1 cpuregs_reg_9__17_  (
    .CK(clk),
    .D(_01102_),
    .Q(\cpuregs[9] [17]),
    .QN(_28086_)
  );
  DFF_X1 cpuregs_reg_9__18_  (
    .CK(clk),
    .D(_01103_),
    .Q(\cpuregs[9] [18]),
    .QN(_28085_)
  );
  DFF_X1 cpuregs_reg_9__19_  (
    .CK(clk),
    .D(_01104_),
    .Q(\cpuregs[9] [19]),
    .QN(_28084_)
  );
  DFF_X1 cpuregs_reg_9__1_  (
    .CK(clk),
    .D(_01086_),
    .Q(\cpuregs[9] [1]),
    .QN(_28102_)
  );
  DFF_X1 cpuregs_reg_9__20_  (
    .CK(clk),
    .D(_01105_),
    .Q(\cpuregs[9] [20]),
    .QN(_28083_)
  );
  DFF_X1 cpuregs_reg_9__21_  (
    .CK(clk),
    .D(_01106_),
    .Q(\cpuregs[9] [21]),
    .QN(_28082_)
  );
  DFF_X1 cpuregs_reg_9__22_  (
    .CK(clk),
    .D(_01107_),
    .Q(\cpuregs[9] [22]),
    .QN(_28081_)
  );
  DFF_X1 cpuregs_reg_9__23_  (
    .CK(clk),
    .D(_01108_),
    .Q(\cpuregs[9] [23]),
    .QN(_28080_)
  );
  DFF_X1 cpuregs_reg_9__24_  (
    .CK(clk),
    .D(_01109_),
    .Q(\cpuregs[9] [24]),
    .QN(_28079_)
  );
  DFF_X1 cpuregs_reg_9__25_  (
    .CK(clk),
    .D(_01110_),
    .Q(\cpuregs[9] [25]),
    .QN(_28078_)
  );
  DFF_X1 cpuregs_reg_9__26_  (
    .CK(clk),
    .D(_01111_),
    .Q(\cpuregs[9] [26]),
    .QN(_28077_)
  );
  DFF_X1 cpuregs_reg_9__27_  (
    .CK(clk),
    .D(_01112_),
    .Q(\cpuregs[9] [27]),
    .QN(_28076_)
  );
  DFF_X1 cpuregs_reg_9__28_  (
    .CK(clk),
    .D(_01113_),
    .Q(\cpuregs[9] [28]),
    .QN(_28075_)
  );
  DFF_X1 cpuregs_reg_9__29_  (
    .CK(clk),
    .D(_01114_),
    .Q(\cpuregs[9] [29]),
    .QN(_28074_)
  );
  DFF_X1 cpuregs_reg_9__2_  (
    .CK(clk),
    .D(_01087_),
    .Q(\cpuregs[9] [2]),
    .QN(_28101_)
  );
  DFF_X1 cpuregs_reg_9__30_  (
    .CK(clk),
    .D(_01115_),
    .Q(\cpuregs[9] [30]),
    .QN(_28073_)
  );
  DFF_X1 cpuregs_reg_9__31_  (
    .CK(clk),
    .D(_00495_),
    .Q(\cpuregs[9] [31]),
    .QN(_28693_)
  );
  DFF_X1 cpuregs_reg_9__3_  (
    .CK(clk),
    .D(_01088_),
    .Q(\cpuregs[9] [3]),
    .QN(_28100_)
  );
  DFF_X1 cpuregs_reg_9__4_  (
    .CK(clk),
    .D(_01089_),
    .Q(\cpuregs[9] [4]),
    .QN(_28099_)
  );
  DFF_X1 cpuregs_reg_9__5_  (
    .CK(clk),
    .D(_01090_),
    .Q(\cpuregs[9] [5]),
    .QN(_28098_)
  );
  DFF_X1 cpuregs_reg_9__6_  (
    .CK(clk),
    .D(_01091_),
    .Q(\cpuregs[9] [6]),
    .QN(_28097_)
  );
  DFF_X1 cpuregs_reg_9__7_  (
    .CK(clk),
    .D(_01092_),
    .Q(\cpuregs[9] [7]),
    .QN(_28096_)
  );
  DFF_X1 cpuregs_reg_9__8_  (
    .CK(clk),
    .D(_01093_),
    .Q(\cpuregs[9] [8]),
    .QN(_28095_)
  );
  DFF_X1 cpuregs_reg_9__9_  (
    .CK(clk),
    .D(_01094_),
    .Q(\cpuregs[9] [9]),
    .QN(_28094_)
  );
  DFF_X1 decoded_imm_reg_0_  (
    .CK(clk),
    .D(_00406_),
    .Q(decoded_imm[0]),
    .QN(_28772_)
  );
  DFF_X1 decoded_imm_reg_10_  (
    .CK(clk),
    .D(_01540_),
    .Q(decoded_imm[10]),
    .QN(_27648_)
  );
  DFF_X1 decoded_imm_reg_11_  (
    .CK(clk),
    .D(_01539_),
    .Q(decoded_imm[11]),
    .QN(_27649_)
  );
  DFF_X1 decoded_imm_reg_12_  (
    .CK(clk),
    .D(_01538_),
    .Q(decoded_imm[12]),
    .QN(_27650_)
  );
  DFF_X1 decoded_imm_reg_13_  (
    .CK(clk),
    .D(_01537_),
    .Q(decoded_imm[13]),
    .QN(_27651_)
  );
  DFF_X1 decoded_imm_reg_14_  (
    .CK(clk),
    .D(_01536_),
    .Q(decoded_imm[14]),
    .QN(_27652_)
  );
  DFF_X1 decoded_imm_reg_15_  (
    .CK(clk),
    .D(_01535_),
    .Q(decoded_imm[15]),
    .QN(_27653_)
  );
  DFF_X1 decoded_imm_reg_16_  (
    .CK(clk),
    .D(_01534_),
    .Q(decoded_imm[16]),
    .QN(_27654_)
  );
  DFF_X1 decoded_imm_reg_17_  (
    .CK(clk),
    .D(_01533_),
    .Q(decoded_imm[17]),
    .QN(_27655_)
  );
  DFF_X1 decoded_imm_reg_18_  (
    .CK(clk),
    .D(_01532_),
    .Q(decoded_imm[18]),
    .QN(_27656_)
  );
  DFF_X1 decoded_imm_reg_19_  (
    .CK(clk),
    .D(_01531_),
    .Q(decoded_imm[19]),
    .QN(_27657_)
  );
  DFF_X1 decoded_imm_reg_1_  (
    .CK(clk),
    .D(_01549_),
    .Q(decoded_imm[1]),
    .QN(_27639_)
  );
  DFF_X1 decoded_imm_reg_20_  (
    .CK(clk),
    .D(_01530_),
    .Q(decoded_imm[20]),
    .QN(_27658_)
  );
  DFF_X1 decoded_imm_reg_21_  (
    .CK(clk),
    .D(_01529_),
    .Q(decoded_imm[21]),
    .QN(_27659_)
  );
  DFF_X1 decoded_imm_reg_22_  (
    .CK(clk),
    .D(_01528_),
    .Q(decoded_imm[22]),
    .QN(_27660_)
  );
  DFF_X1 decoded_imm_reg_23_  (
    .CK(clk),
    .D(_01527_),
    .Q(decoded_imm[23]),
    .QN(_27661_)
  );
  DFF_X1 decoded_imm_reg_24_  (
    .CK(clk),
    .D(_01526_),
    .Q(decoded_imm[24]),
    .QN(_27662_)
  );
  DFF_X1 decoded_imm_reg_25_  (
    .CK(clk),
    .D(_01525_),
    .Q(decoded_imm[25]),
    .QN(_27663_)
  );
  DFF_X1 decoded_imm_reg_26_  (
    .CK(clk),
    .D(_01524_),
    .Q(decoded_imm[26]),
    .QN(_27664_)
  );
  DFF_X1 decoded_imm_reg_27_  (
    .CK(clk),
    .D(_01523_),
    .Q(decoded_imm[27]),
    .QN(_27665_)
  );
  DFF_X1 decoded_imm_reg_28_  (
    .CK(clk),
    .D(_01522_),
    .Q(decoded_imm[28]),
    .QN(_27666_)
  );
  DFF_X1 decoded_imm_reg_29_  (
    .CK(clk),
    .D(_01521_),
    .Q(decoded_imm[29]),
    .QN(_27667_)
  );
  DFF_X1 decoded_imm_reg_2_  (
    .CK(clk),
    .D(_01548_),
    .Q(decoded_imm[2]),
    .QN(_27640_)
  );
  DFF_X1 decoded_imm_reg_30_  (
    .CK(clk),
    .D(_01520_),
    .Q(decoded_imm[30]),
    .QN(_27668_)
  );
  DFF_X1 decoded_imm_reg_31_  (
    .CK(clk),
    .D(_01519_),
    .Q(decoded_imm[31]),
    .QN(_27669_)
  );
  DFF_X1 decoded_imm_reg_3_  (
    .CK(clk),
    .D(_01547_),
    .Q(decoded_imm[3]),
    .QN(_27641_)
  );
  DFF_X1 decoded_imm_reg_4_  (
    .CK(clk),
    .D(_01546_),
    .Q(decoded_imm[4]),
    .QN(_27642_)
  );
  DFF_X1 decoded_imm_reg_5_  (
    .CK(clk),
    .D(_01545_),
    .Q(decoded_imm[5]),
    .QN(_27643_)
  );
  DFF_X1 decoded_imm_reg_6_  (
    .CK(clk),
    .D(_01544_),
    .Q(decoded_imm[6]),
    .QN(_27644_)
  );
  DFF_X1 decoded_imm_reg_7_  (
    .CK(clk),
    .D(_01543_),
    .Q(decoded_imm[7]),
    .QN(_27645_)
  );
  DFF_X1 decoded_imm_reg_8_  (
    .CK(clk),
    .D(_01542_),
    .Q(decoded_imm[8]),
    .QN(_27646_)
  );
  DFF_X1 decoded_imm_reg_9_  (
    .CK(clk),
    .D(_01541_),
    .Q(decoded_imm[9]),
    .QN(_27647_)
  );
  DFF_X1 decoded_imm_j_reg_10_  (
    .CK(clk),
    .D(_00407_),
    .Q(decoded_imm_j[10]),
    .QN(_29143_)
  );
  DFF_X1 decoded_imm_j_reg_12_  (
    .CK(clk),
    .D(_01559_),
    .Q(decoded_imm_j[12]),
    .QN(_27630_)
  );
  DFF_X1 decoded_imm_j_reg_13_  (
    .CK(clk),
    .D(_01560_),
    .Q(decoded_imm_j[13]),
    .QN(_27629_)
  );
  DFF_X1 decoded_imm_j_reg_14_  (
    .CK(clk),
    .D(_01561_),
    .Q(decoded_imm_j[14]),
    .QN(_27628_)
  );
  DFF_X1 decoded_imm_j_reg_18_  (
    .CK(clk),
    .D(_01562_),
    .Q(decoded_imm_j[18]),
    .QN(_27627_)
  );
  DFF_X1 decoded_imm_j_reg_19_  (
    .CK(clk),
    .D(_01563_),
    .Q(decoded_imm_j[19]),
    .QN(_27626_)
  );
  DFF_X1 decoded_imm_j_reg_30_  (
    .CK(clk),
    .D(_01557_),
    .Q(decoded_imm_j[30]),
    .QN(_27632_)
  );
  DFF_X1 decoded_imm_j_reg_4_  (
    .CK(clk),
    .D(_01558_),
    .Q(decoded_imm_j[4]),
    .QN(_27631_)
  );
  DFF_X1 decoded_imm_j_reg_5_  (
    .CK(clk),
    .D(_01554_),
    .Q(decoded_imm_j[5]),
    .QN(_27635_)
  );
  DFF_X1 decoded_imm_j_reg_6_  (
    .CK(clk),
    .D(_01553_),
    .Q(decoded_imm_j[6]),
    .QN(_27636_)
  );
  DFF_X1 decoded_imm_j_reg_7_  (
    .CK(clk),
    .D(_01552_),
    .Q(decoded_imm_j[7]),
    .QN(_27637_)
  );
  DFF_X1 decoded_imm_j_reg_8_  (
    .CK(clk),
    .D(_01555_),
    .Q(decoded_imm_j[8]),
    .QN(_27634_)
  );
  DFF_X1 decoded_imm_j_reg_9_  (
    .CK(clk),
    .D(_01556_),
    .Q(decoded_imm_j[9]),
    .QN(_27633_)
  );
  DFF_X1 decoded_rd_reg_0_  (
    .CK(clk),
    .D(_00397_),
    .Q(decoded_rd[0]),
    .QN(_28781_)
  );
  DFF_X1 decoded_rd_reg_1_  (
    .CK(clk),
    .D(_00398_),
    .Q(decoded_rd[1]),
    .QN(_28780_)
  );
  DFF_X1 decoded_rd_reg_2_  (
    .CK(clk),
    .D(_00399_),
    .Q(decoded_rd[2]),
    .QN(_28779_)
  );
  DFF_X1 decoded_rd_reg_3_  (
    .CK(clk),
    .D(_00400_),
    .Q(decoded_rd[3]),
    .QN(_28778_)
  );
  DFF_X1 decoded_rd_reg_4_  (
    .CK(clk),
    .D(_00401_),
    .Q(decoded_rd[4]),
    .QN(_28777_)
  );
  DFF_X1 decoded_rs1_reg_0_  (
    .CK(clk),
    .D(_01564_),
    .Q(decoded_rs1[0]),
    .QN(_27625_)
  );
  DFF_X1 decoded_rs1_reg_1_  (
    .CK(clk),
    .D(_01565_),
    .Q(decoded_rs1[1]),
    .QN(_27624_)
  );
  DFF_X1 decoded_rs1_reg_2_  (
    .CK(clk),
    .D(_01566_),
    .Q(decoded_rs1[2]),
    .QN(_27623_)
  );
  DFF_X1 decoded_rs2_reg_0_  (
    .CK(clk),
    .D(_00402_),
    .Q(decoded_rs2[0]),
    .QN(_28776_)
  );
  DFF_X1 decoded_rs2_reg_1_  (
    .CK(clk),
    .D(_00403_),
    .Q(decoded_rs2[1]),
    .QN(_28775_)
  );
  DFF_X1 decoded_rs2_reg_2_  (
    .CK(clk),
    .D(_00404_),
    .Q(decoded_rs2[2]),
    .QN(_28774_)
  );
  DFF_X1 decoded_rs2_reg_3_  (
    .CK(clk),
    .D(_00405_),
    .Q(decoded_rs2[3]),
    .QN(_28773_)
  );
  DFF_X1 decoder_pseudo_trigger_reg  (
    .CK(clk),
    .D(_01550_),
    .Q(decoder_pseudo_trigger),
    .QN(_00017_)
  );
  DFF_X1 decoder_trigger_reg  (
    .CK(clk),
    .D(_00000_),
    .Q(decoder_trigger),
    .QN(_00033_)
  );
  DFF_X1 eoi_reg_30_  (
    .CK(clk),
    .D(_00152_),
    .Q(eoi[30]),
    .QN(_28975_)
  );
  DFF_X1 instr_add_reg  (
    .CK(clk),
    .D(_00381_),
    .Q(instr_add),
    .QN(_28797_)
  );
  DFF_X1 instr_addi_reg  (
    .CK(clk),
    .D(_00372_),
    .Q(instr_addi),
    .QN(_28806_)
  );
  DFF_X1 instr_and_reg  (
    .CK(clk),
    .D(_00390_),
    .Q(instr_and),
    .QN(_28788_)
  );
  DFF_X1 instr_andi_reg  (
    .CK(clk),
    .D(_00377_),
    .Q(instr_andi),
    .QN(_28801_)
  );
  DFF_X1 instr_auipc_reg  (
    .CK(clk),
    .D(_00356_),
    .Q(instr_auipc),
    .QN(_28820_)
  );
  DFF_X1 instr_beq_reg  (
    .CK(clk),
    .D(_00358_),
    .Q(instr_beq),
    .QN(_28819_)
  );
  DFF_X1 instr_bge_reg  (
    .CK(clk),
    .D(_00361_),
    .Q(instr_bge),
    .QN(_28816_)
  );
  DFF_X1 instr_bgeu_reg  (
    .CK(clk),
    .D(_00363_),
    .Q(instr_bgeu),
    .QN(_28814_)
  );
  DFF_X1 instr_blt_reg  (
    .CK(clk),
    .D(_00360_),
    .Q(instr_blt),
    .QN(_28817_)
  );
  DFF_X1 instr_bltu_reg  (
    .CK(clk),
    .D(_00362_),
    .Q(instr_bltu),
    .QN(_28815_)
  );
  DFF_X1 instr_bne_reg  (
    .CK(clk),
    .D(_00359_),
    .Q(instr_bne),
    .QN(_28818_)
  );
  DFF_X1 instr_fence_reg  (
    .CK(clk),
    .D(_00396_),
    .Q(instr_fence),
    .QN(_28782_)
  );
  DFF_X1 instr_jal_reg  (
    .CK(clk),
    .D(_00357_),
    .Q(instr_jal),
    .QN(_00029_)
  );
  DFF_X1 instr_jalr_reg  (
    .CK(clk),
    .D(_00364_),
    .Q(instr_jalr),
    .QN(_00028_)
  );
  DFF_X1 instr_lb_reg  (
    .CK(clk),
    .D(_00365_),
    .Q(instr_lb),
    .QN(_28813_)
  );
  DFF_X1 instr_lbu_reg  (
    .CK(clk),
    .D(_00368_),
    .Q(instr_lbu),
    .QN(_28810_)
  );
  DFF_X1 instr_lh_reg  (
    .CK(clk),
    .D(_00366_),
    .Q(instr_lh),
    .QN(_28812_)
  );
  DFF_X1 instr_lhu_reg  (
    .CK(clk),
    .D(_00369_),
    .Q(instr_lhu),
    .QN(_28809_)
  );
  DFF_X1 instr_lui_reg  (
    .CK(clk),
    .D(_00355_),
    .Q(instr_lui),
    .QN(_28821_)
  );
  DFF_X1 instr_lw_reg  (
    .CK(clk),
    .D(_00367_),
    .Q(instr_lw),
    .QN(_28811_)
  );
  DFF_X1 instr_or_reg  (
    .CK(clk),
    .D(_00389_),
    .Q(instr_or),
    .QN(_28789_)
  );
  DFF_X1 instr_ori_reg  (
    .CK(clk),
    .D(_00376_),
    .Q(instr_ori),
    .QN(_28802_)
  );
  DFF_X1 instr_rdcycle_reg  (
    .CK(clk),
    .D(_00392_),
    .Q(instr_rdcycle),
    .QN(_28786_)
  );
  DFF_X1 instr_rdcycleh_reg  (
    .CK(clk),
    .D(_00393_),
    .Q(instr_rdcycleh),
    .QN(_28785_)
  );
  DFF_X1 instr_rdinstr_reg  (
    .CK(clk),
    .D(_00394_),
    .Q(instr_rdinstr),
    .QN(_28784_)
  );
  DFF_X1 instr_rdinstrh_reg  (
    .CK(clk),
    .D(_00395_),
    .Q(instr_rdinstrh),
    .QN(_28783_)
  );
  DFF_X1 instr_sb_reg  (
    .CK(clk),
    .D(_00378_),
    .Q(instr_sb),
    .QN(_28800_)
  );
  DFF_X1 instr_sh_reg  (
    .CK(clk),
    .D(_00371_),
    .Q(instr_sh),
    .QN(_28807_)
  );
  DFF_X1 instr_sll_reg  (
    .CK(clk),
    .D(_00383_),
    .Q(instr_sll),
    .QN(_28795_)
  );
  DFF_X1 instr_slli_reg  (
    .CK(clk),
    .D(_00379_),
    .Q(instr_slli),
    .QN(_28799_)
  );
  DFF_X1 instr_slt_reg  (
    .CK(clk),
    .D(_00384_),
    .Q(instr_slt),
    .QN(_28794_)
  );
  DFF_X1 instr_slti_reg  (
    .CK(clk),
    .D(_00373_),
    .Q(instr_slti),
    .QN(_28805_)
  );
  DFF_X1 instr_sltiu_reg  (
    .CK(clk),
    .D(_00374_),
    .Q(instr_sltiu),
    .QN(_28804_)
  );
  DFF_X1 instr_sltu_reg  (
    .CK(clk),
    .D(_00385_),
    .Q(instr_sltu),
    .QN(_28793_)
  );
  DFF_X1 instr_sra_reg  (
    .CK(clk),
    .D(_00388_),
    .Q(instr_sra),
    .QN(_28790_)
  );
  DFF_X1 instr_srai_reg  (
    .CK(clk),
    .D(_00391_),
    .Q(instr_srai),
    .QN(_28787_)
  );
  DFF_X1 instr_srl_reg  (
    .CK(clk),
    .D(_00387_),
    .Q(instr_srl),
    .QN(_28791_)
  );
  DFF_X1 instr_srli_reg  (
    .CK(clk),
    .D(_00380_),
    .Q(instr_srli),
    .QN(_28798_)
  );
  DFF_X1 instr_sub_reg  (
    .CK(clk),
    .D(_00382_),
    .Q(instr_sub),
    .QN(_28796_)
  );
  DFF_X1 instr_sw_reg  (
    .CK(clk),
    .D(_00153_),
    .Q(instr_sw),
    .QN(_28974_)
  );
  DFF_X1 instr_xor_reg  (
    .CK(clk),
    .D(_00386_),
    .Q(instr_xor),
    .QN(_28792_)
  );
  DFF_X1 instr_xori_reg  (
    .CK(clk),
    .D(_00375_),
    .Q(instr_xori),
    .QN(_28803_)
  );
  DFF_X1 is_alu_reg_imm_reg  (
    .CK(clk),
    .D(_00414_),
    .Q(is_alu_reg_imm),
    .QN(_28765_)
  );
  DFF_X1 is_alu_reg_reg_reg  (
    .CK(clk),
    .D(_00417_),
    .Q(is_alu_reg_reg),
    .QN(_28762_)
  );
  DFF_X1 is_beq_bne_blt_bge_bltu_bgeu_reg  (
    .CK(clk),
    .D(_00412_),
    .Q(is_beq_bne_blt_bge_bltu_bgeu),
    .QN(_00047_)
  );
  DFF_X1 is_compare_reg  (
    .CK(clk),
    .D(_00416_),
    .Q(is_compare),
    .QN(_28763_)
  );
  DFF_X1 is_jalr_addi_slti_sltiu_xori_ori_andi_reg  (
    .CK(clk),
    .D(_00415_),
    .Q(is_jalr_addi_slti_sltiu_xori_ori_andi),
    .QN(_28764_)
  );
  DFF_X1 is_lb_lh_lw_lbu_lhu_reg  (
    .CK(clk),
    .D(_00408_),
    .Q(is_lb_lh_lw_lbu_lhu),
    .QN(_28770_)
  );
  DFF_X1 is_lbu_lhu_lw_reg  (
    .CK(clk),
    .D(_00001_),
    .Q(is_lbu_lhu_lw),
    .QN(_28767_)
  );
  DFF_X1 is_lui_auipc_jal_reg  (
    .CK(clk),
    .D(_00002_),
    .Q(is_lui_auipc_jal),
    .QN(_28771_)
  );
  DFF_X1 is_lui_auipc_jal_jalr_addi_add_sub_reg  (
    .CK(clk),
    .D(_00413_),
    .Q(is_lui_auipc_jal_jalr_addi_add_sub),
    .QN(_28766_)
  );
  DFF_X1 is_sb_sh_sw_reg  (
    .CK(clk),
    .D(_00410_),
    .Q(is_sb_sh_sw),
    .QN(_28769_)
  );
  DFF_X1 is_sll_srl_sra_reg  (
    .CK(clk),
    .D(_00411_),
    .Q(is_sll_srl_sra),
    .QN(_00046_)
  );
  DFF_X1 is_slli_srli_srai_reg  (
    .CK(clk),
    .D(_00409_),
    .Q(is_slli_srli_srai),
    .QN(_00027_)
  );
  DFF_X1 is_slti_blt_slt_reg  (
    .CK(clk),
    .D(_00003_),
    .Q(is_slti_blt_slt),
    .QN(_29144_)
  );
  DFF_X1 is_sltiu_bltu_sltu_reg  (
    .CK(clk),
    .D(_00004_),
    .Q(is_sltiu_bltu_sltu),
    .QN(_28768_)
  );
  DFF_X1 latched_branch_reg  (
    .CK(clk),
    .D(_00346_),
    .Q(latched_branch),
    .QN(_00030_)
  );
  DFF_X1 latched_is_lb_reg  (
    .CK(clk),
    .D(_00349_),
    .Q(latched_is_lb),
    .QN(_28827_)
  );
  DFF_X1 latched_is_lh_reg  (
    .CK(clk),
    .D(_00348_),
    .Q(latched_is_lh),
    .QN(_28828_)
  );
  DFF_X1 latched_is_lu_reg  (
    .CK(clk),
    .D(_00347_),
    .Q(latched_is_lu),
    .QN(_28829_)
  );
  DFF_X1 latched_rd_reg_0_  (
    .CK(clk),
    .D(_00350_),
    .Q(latched_rd[0]),
    .QN(_28826_)
  );
  DFF_X1 latched_rd_reg_1_  (
    .CK(clk),
    .D(_00351_),
    .Q(latched_rd[1]),
    .QN(_28825_)
  );
  DFF_X1 latched_rd_reg_2_  (
    .CK(clk),
    .D(_00352_),
    .Q(latched_rd[2]),
    .QN(_28824_)
  );
  DFF_X1 latched_rd_reg_3_  (
    .CK(clk),
    .D(_00353_),
    .Q(latched_rd[3]),
    .QN(_28823_)
  );
  DFF_X1 latched_rd_reg_4_  (
    .CK(clk),
    .D(_00354_),
    .Q(latched_rd[4]),
    .QN(_29111_)
  );
  DFF_X1 latched_stalu_reg  (
    .CK(clk),
    .D(_00345_),
    .Q(latched_stalu),
    .QN(_28830_)
  );
  DFF_X1 latched_store_reg  (
    .CK(clk),
    .D(_00344_),
    .Q(latched_store),
    .QN(_28831_)
  );
  DFF_X1 mem_addr_reg_10_  (
    .CK(clk),
    .D(_00428_),
    .Q(mem_addr[10]),
    .QN(_28751_)
  );
  DFF_X1 mem_addr_reg_11_  (
    .CK(clk),
    .D(_00429_),
    .Q(mem_addr[11]),
    .QN(_28750_)
  );
  DFF_X1 mem_addr_reg_12_  (
    .CK(clk),
    .D(_00430_),
    .Q(mem_addr[12]),
    .QN(_28749_)
  );
  DFF_X1 mem_addr_reg_13_  (
    .CK(clk),
    .D(_00431_),
    .Q(mem_addr[13]),
    .QN(_28748_)
  );
  DFF_X1 mem_addr_reg_14_  (
    .CK(clk),
    .D(_00432_),
    .Q(mem_addr[14]),
    .QN(_28747_)
  );
  DFF_X1 mem_addr_reg_15_  (
    .CK(clk),
    .D(_00433_),
    .Q(mem_addr[15]),
    .QN(_28746_)
  );
  DFF_X1 mem_addr_reg_16_  (
    .CK(clk),
    .D(_00434_),
    .Q(mem_addr[16]),
    .QN(_28745_)
  );
  DFF_X1 mem_addr_reg_17_  (
    .CK(clk),
    .D(_00435_),
    .Q(mem_addr[17]),
    .QN(_28744_)
  );
  DFF_X1 mem_addr_reg_18_  (
    .CK(clk),
    .D(_00436_),
    .Q(mem_addr[18]),
    .QN(_28743_)
  );
  DFF_X1 mem_addr_reg_19_  (
    .CK(clk),
    .D(_00437_),
    .Q(mem_addr[19]),
    .QN(_28742_)
  );
  DFF_X1 mem_addr_reg_20_  (
    .CK(clk),
    .D(_00438_),
    .Q(mem_addr[20]),
    .QN(_28741_)
  );
  DFF_X1 mem_addr_reg_21_  (
    .CK(clk),
    .D(_00439_),
    .Q(mem_addr[21]),
    .QN(_28740_)
  );
  DFF_X1 mem_addr_reg_22_  (
    .CK(clk),
    .D(_00440_),
    .Q(mem_addr[22]),
    .QN(_28739_)
  );
  DFF_X1 mem_addr_reg_23_  (
    .CK(clk),
    .D(_00441_),
    .Q(mem_addr[23]),
    .QN(_28738_)
  );
  DFF_X1 mem_addr_reg_24_  (
    .CK(clk),
    .D(_00442_),
    .Q(mem_addr[24]),
    .QN(_28737_)
  );
  DFF_X1 mem_addr_reg_25_  (
    .CK(clk),
    .D(_00443_),
    .Q(mem_addr[25]),
    .QN(_28736_)
  );
  DFF_X1 mem_addr_reg_26_  (
    .CK(clk),
    .D(_00444_),
    .Q(mem_addr[26]),
    .QN(_28735_)
  );
  DFF_X1 mem_addr_reg_27_  (
    .CK(clk),
    .D(_00445_),
    .Q(mem_addr[27]),
    .QN(_28734_)
  );
  DFF_X1 mem_addr_reg_28_  (
    .CK(clk),
    .D(_00446_),
    .Q(mem_addr[28]),
    .QN(_28733_)
  );
  DFF_X1 mem_addr_reg_29_  (
    .CK(clk),
    .D(_00447_),
    .Q(mem_addr[29]),
    .QN(_28732_)
  );
  DFF_X1 mem_addr_reg_2_  (
    .CK(clk),
    .D(_00420_),
    .Q(mem_addr[2]),
    .QN(_28759_)
  );
  DFF_X1 mem_addr_reg_30_  (
    .CK(clk),
    .D(_00448_),
    .Q(mem_addr[30]),
    .QN(_28731_)
  );
  DFF_X1 mem_addr_reg_31_  (
    .CK(clk),
    .D(_00449_),
    .Q(mem_addr[31]),
    .QN(_28730_)
  );
  DFF_X1 mem_addr_reg_3_  (
    .CK(clk),
    .D(_00421_),
    .Q(mem_addr[3]),
    .QN(_28758_)
  );
  DFF_X1 mem_addr_reg_4_  (
    .CK(clk),
    .D(_00422_),
    .Q(mem_addr[4]),
    .QN(_28757_)
  );
  DFF_X1 mem_addr_reg_5_  (
    .CK(clk),
    .D(_00423_),
    .Q(mem_addr[5]),
    .QN(_28756_)
  );
  DFF_X1 mem_addr_reg_6_  (
    .CK(clk),
    .D(_00424_),
    .Q(mem_addr[6]),
    .QN(_28755_)
  );
  DFF_X1 mem_addr_reg_7_  (
    .CK(clk),
    .D(_00425_),
    .Q(mem_addr[7]),
    .QN(_28754_)
  );
  DFF_X1 mem_addr_reg_8_  (
    .CK(clk),
    .D(_00426_),
    .Q(mem_addr[8]),
    .QN(_28753_)
  );
  DFF_X1 mem_addr_reg_9_  (
    .CK(clk),
    .D(_00427_),
    .Q(mem_addr[9]),
    .QN(_28752_)
  );
  DFF_X1 mem_do_prefetch_reg  (
    .CK(clk),
    .D(_00338_),
    .Q(mem_do_prefetch),
    .QN(_00035_)
  );
  DFF_X1 mem_do_rdata_reg  (
    .CK(clk),
    .D(_00340_),
    .Q(mem_do_rdata),
    .QN(_00034_)
  );
  DFF_X1 mem_do_rinst_reg  (
    .CK(clk),
    .D(_00339_),
    .Q(mem_do_rinst),
    .QN(_28832_)
  );
  DFF_X1 mem_do_wdata_reg  (
    .CK(clk),
    .D(_00341_),
    .Q(mem_do_wdata),
    .QN(_00045_)
  );
  DFF_X1 mem_instr_reg  (
    .CK(clk),
    .D(_00418_),
    .Q(mem_instr),
    .QN(_28761_)
  );
  DFF_X1 mem_rdata_q_reg_0_  (
    .CK(clk),
    .D(_00488_),
    .Q(mem_rdata_q[0]),
    .QN(_00024_)
  );
  DFF_X1 mem_rdata_q_reg_10_  (
    .CK(clk),
    .D(_00316_),
    .Q(mem_rdata_q[10]),
    .QN(_28846_)
  );
  DFF_X1 mem_rdata_q_reg_11_  (
    .CK(clk),
    .D(_00317_),
    .Q(mem_rdata_q[11]),
    .QN(_28845_)
  );
  DFF_X1 mem_rdata_q_reg_12_  (
    .CK(clk),
    .D(_00318_),
    .Q(mem_rdata_q[12]),
    .QN(_00043_)
  );
  DFF_X1 mem_rdata_q_reg_13_  (
    .CK(clk),
    .D(_00319_),
    .Q(mem_rdata_q[13]),
    .QN(_00042_)
  );
  DFF_X1 mem_rdata_q_reg_14_  (
    .CK(clk),
    .D(_00320_),
    .Q(mem_rdata_q[14]),
    .QN(_00041_)
  );
  DFF_X1 mem_rdata_q_reg_15_  (
    .CK(clk),
    .D(_00321_),
    .Q(mem_rdata_q[15]),
    .QN(_28844_)
  );
  DFF_X1 mem_rdata_q_reg_16_  (
    .CK(clk),
    .D(_00322_),
    .Q(mem_rdata_q[16]),
    .QN(_28843_)
  );
  DFF_X1 mem_rdata_q_reg_17_  (
    .CK(clk),
    .D(_00323_),
    .Q(mem_rdata_q[17]),
    .QN(_28842_)
  );
  DFF_X1 mem_rdata_q_reg_18_  (
    .CK(clk),
    .D(_00324_),
    .Q(mem_rdata_q[18]),
    .QN(_28841_)
  );
  DFF_X1 mem_rdata_q_reg_19_  (
    .CK(clk),
    .D(_00325_),
    .Q(mem_rdata_q[19]),
    .QN(_28840_)
  );
  DFF_X1 mem_rdata_q_reg_1_  (
    .CK(clk),
    .D(_00489_),
    .Q(mem_rdata_q[1]),
    .QN(_00023_)
  );
  DFF_X1 mem_rdata_q_reg_20_  (
    .CK(clk),
    .D(_00326_),
    .Q(mem_rdata_q[20]),
    .QN(_00040_)
  );
  DFF_X1 mem_rdata_q_reg_21_  (
    .CK(clk),
    .D(_00327_),
    .Q(mem_rdata_q[21]),
    .QN(_00039_)
  );
  DFF_X1 mem_rdata_q_reg_22_  (
    .CK(clk),
    .D(_00328_),
    .Q(mem_rdata_q[22]),
    .QN(_28839_)
  );
  DFF_X1 mem_rdata_q_reg_23_  (
    .CK(clk),
    .D(_00329_),
    .Q(mem_rdata_q[23]),
    .QN(_28838_)
  );
  DFF_X1 mem_rdata_q_reg_24_  (
    .CK(clk),
    .D(_00330_),
    .Q(mem_rdata_q[24]),
    .QN(_28837_)
  );
  DFF_X1 mem_rdata_q_reg_25_  (
    .CK(clk),
    .D(_00331_),
    .Q(mem_rdata_q[25]),
    .QN(_28836_)
  );
  DFF_X1 mem_rdata_q_reg_26_  (
    .CK(clk),
    .D(_00332_),
    .Q(mem_rdata_q[26]),
    .QN(_28835_)
  );
  DFF_X1 mem_rdata_q_reg_27_  (
    .CK(clk),
    .D(_00333_),
    .Q(mem_rdata_q[27]),
    .QN(_00038_)
  );
  DFF_X1 mem_rdata_q_reg_28_  (
    .CK(clk),
    .D(_00334_),
    .Q(mem_rdata_q[28]),
    .QN(_28834_)
  );
  DFF_X1 mem_rdata_q_reg_29_  (
    .CK(clk),
    .D(_00335_),
    .Q(mem_rdata_q[29]),
    .QN(_28833_)
  );
  DFF_X1 mem_rdata_q_reg_2_  (
    .CK(clk),
    .D(_00490_),
    .Q(mem_rdata_q[2]),
    .QN(_00022_)
  );
  DFF_X1 mem_rdata_q_reg_30_  (
    .CK(clk),
    .D(_00336_),
    .Q(mem_rdata_q[30]),
    .QN(_00037_)
  );
  DFF_X1 mem_rdata_q_reg_31_  (
    .CK(clk),
    .D(_00337_),
    .Q(mem_rdata_q[31]),
    .QN(_00036_)
  );
  DFF_X1 mem_rdata_q_reg_3_  (
    .CK(clk),
    .D(_00491_),
    .Q(mem_rdata_q[3]),
    .QN(_00021_)
  );
  DFF_X1 mem_rdata_q_reg_4_  (
    .CK(clk),
    .D(_00492_),
    .Q(mem_rdata_q[4]),
    .QN(_00020_)
  );
  DFF_X1 mem_rdata_q_reg_5_  (
    .CK(clk),
    .D(_00493_),
    .Q(mem_rdata_q[5]),
    .QN(_00019_)
  );
  DFF_X1 mem_rdata_q_reg_6_  (
    .CK(clk),
    .D(_00494_),
    .Q(mem_rdata_q[6]),
    .QN(_00018_)
  );
  DFF_X1 mem_rdata_q_reg_7_  (
    .CK(clk),
    .D(_00313_),
    .Q(mem_rdata_q[7]),
    .QN(_28849_)
  );
  DFF_X1 mem_rdata_q_reg_8_  (
    .CK(clk),
    .D(_00314_),
    .Q(mem_rdata_q[8]),
    .QN(_28848_)
  );
  DFF_X1 mem_rdata_q_reg_9_  (
    .CK(clk),
    .D(_00315_),
    .Q(mem_rdata_q[9]),
    .QN(_28847_)
  );
  DFF_X1 mem_state_reg_0_  (
    .CK(clk),
    .D(_00486_),
    .Q(mem_state[0]),
    .QN(_00026_)
  );
  DFF_X1 mem_state_reg_1_  (
    .CK(clk),
    .D(_00487_),
    .Q(mem_state[1]),
    .QN(_00025_)
  );
  DFF_X1 mem_valid_reg  (
    .CK(clk),
    .D(_00419_),
    .Q(mem_valid),
    .QN(_28760_)
  );
  DFF_X1 mem_wdata_reg_0_  (
    .CK(clk),
    .D(_00450_),
    .Q(mem_wdata[0]),
    .QN(_28729_)
  );
  DFF_X1 mem_wdata_reg_10_  (
    .CK(clk),
    .D(_00460_),
    .Q(mem_wdata[10]),
    .QN(_28719_)
  );
  DFF_X1 mem_wdata_reg_11_  (
    .CK(clk),
    .D(_00461_),
    .Q(mem_wdata[11]),
    .QN(_28718_)
  );
  DFF_X1 mem_wdata_reg_12_  (
    .CK(clk),
    .D(_00462_),
    .Q(mem_wdata[12]),
    .QN(_28717_)
  );
  DFF_X1 mem_wdata_reg_13_  (
    .CK(clk),
    .D(_00463_),
    .Q(mem_wdata[13]),
    .QN(_28716_)
  );
  DFF_X1 mem_wdata_reg_14_  (
    .CK(clk),
    .D(_00464_),
    .Q(mem_wdata[14]),
    .QN(_28715_)
  );
  DFF_X1 mem_wdata_reg_15_  (
    .CK(clk),
    .D(_00465_),
    .Q(mem_wdata[15]),
    .QN(_28714_)
  );
  DFF_X1 mem_wdata_reg_16_  (
    .CK(clk),
    .D(_00466_),
    .Q(mem_wdata[16]),
    .QN(_28713_)
  );
  DFF_X1 mem_wdata_reg_17_  (
    .CK(clk),
    .D(_00467_),
    .Q(mem_wdata[17]),
    .QN(_28712_)
  );
  DFF_X1 mem_wdata_reg_18_  (
    .CK(clk),
    .D(_00468_),
    .Q(mem_wdata[18]),
    .QN(_28711_)
  );
  DFF_X1 mem_wdata_reg_19_  (
    .CK(clk),
    .D(_00469_),
    .Q(mem_wdata[19]),
    .QN(_28710_)
  );
  DFF_X1 mem_wdata_reg_1_  (
    .CK(clk),
    .D(_00451_),
    .Q(mem_wdata[1]),
    .QN(_28728_)
  );
  DFF_X1 mem_wdata_reg_20_  (
    .CK(clk),
    .D(_00470_),
    .Q(mem_wdata[20]),
    .QN(_28709_)
  );
  DFF_X1 mem_wdata_reg_21_  (
    .CK(clk),
    .D(_00471_),
    .Q(mem_wdata[21]),
    .QN(_28708_)
  );
  DFF_X1 mem_wdata_reg_22_  (
    .CK(clk),
    .D(_00472_),
    .Q(mem_wdata[22]),
    .QN(_28707_)
  );
  DFF_X1 mem_wdata_reg_23_  (
    .CK(clk),
    .D(_00473_),
    .Q(mem_wdata[23]),
    .QN(_28706_)
  );
  DFF_X1 mem_wdata_reg_24_  (
    .CK(clk),
    .D(_00474_),
    .Q(mem_wdata[24]),
    .QN(_28705_)
  );
  DFF_X1 mem_wdata_reg_25_  (
    .CK(clk),
    .D(_00475_),
    .Q(mem_wdata[25]),
    .QN(_28704_)
  );
  DFF_X1 mem_wdata_reg_26_  (
    .CK(clk),
    .D(_00476_),
    .Q(mem_wdata[26]),
    .QN(_28703_)
  );
  DFF_X1 mem_wdata_reg_27_  (
    .CK(clk),
    .D(_00477_),
    .Q(mem_wdata[27]),
    .QN(_28702_)
  );
  DFF_X1 mem_wdata_reg_28_  (
    .CK(clk),
    .D(_00478_),
    .Q(mem_wdata[28]),
    .QN(_28701_)
  );
  DFF_X1 mem_wdata_reg_29_  (
    .CK(clk),
    .D(_00479_),
    .Q(mem_wdata[29]),
    .QN(_28700_)
  );
  DFF_X1 mem_wdata_reg_2_  (
    .CK(clk),
    .D(_00452_),
    .Q(mem_wdata[2]),
    .QN(_28727_)
  );
  DFF_X1 mem_wdata_reg_30_  (
    .CK(clk),
    .D(_00480_),
    .Q(mem_wdata[30]),
    .QN(_28699_)
  );
  DFF_X1 mem_wdata_reg_31_  (
    .CK(clk),
    .D(_00481_),
    .Q(mem_wdata[31]),
    .QN(_28698_)
  );
  DFF_X1 mem_wdata_reg_3_  (
    .CK(clk),
    .D(_00453_),
    .Q(mem_wdata[3]),
    .QN(_28726_)
  );
  DFF_X1 mem_wdata_reg_4_  (
    .CK(clk),
    .D(_00454_),
    .Q(mem_wdata[4]),
    .QN(_28725_)
  );
  DFF_X1 mem_wdata_reg_5_  (
    .CK(clk),
    .D(_00455_),
    .Q(mem_wdata[5]),
    .QN(_28724_)
  );
  DFF_X1 mem_wdata_reg_6_  (
    .CK(clk),
    .D(_00456_),
    .Q(mem_wdata[6]),
    .QN(_28723_)
  );
  DFF_X1 mem_wdata_reg_7_  (
    .CK(clk),
    .D(_00457_),
    .Q(mem_wdata[7]),
    .QN(_28722_)
  );
  DFF_X1 mem_wdata_reg_8_  (
    .CK(clk),
    .D(_00458_),
    .Q(mem_wdata[8]),
    .QN(_28721_)
  );
  DFF_X1 mem_wdata_reg_9_  (
    .CK(clk),
    .D(_00459_),
    .Q(mem_wdata[9]),
    .QN(_28720_)
  );
  DFF_X1 mem_wordsize_reg_0_  (
    .CK(clk),
    .D(_00342_),
    .Q(mem_wordsize[0]),
    .QN(_00032_)
  );
  DFF_X1 mem_wordsize_reg_1_  (
    .CK(clk),
    .D(_00343_),
    .Q(mem_wordsize[1]),
    .QN(_00031_)
  );
  DFF_X1 mem_wstrb_reg_0_  (
    .CK(clk),
    .D(_00482_),
    .Q(mem_wstrb[0]),
    .QN(_28697_)
  );
  DFF_X1 mem_wstrb_reg_1_  (
    .CK(clk),
    .D(_00483_),
    .Q(mem_wstrb[1]),
    .QN(_28696_)
  );
  DFF_X1 mem_wstrb_reg_2_  (
    .CK(clk),
    .D(_00484_),
    .Q(mem_wstrb[2]),
    .QN(_28695_)
  );
  DFF_X1 mem_wstrb_reg_3_  (
    .CK(clk),
    .D(_00485_),
    .Q(mem_wstrb[3]),
    .QN(_28694_)
  );
  DFF_X1 reg_next_pc_reg_0_  (
    .CK(clk),
    .D(_01551_),
    .Q(reg_next_pc[0]),
    .QN(_27638_)
  );
  DFF_X1 reg_next_pc_reg_10_  (
    .CK(clk),
    .D(_00194_),
    .Q(reg_next_pc[10]),
    .QN(_28934_)
  );
  DFF_X1 reg_next_pc_reg_11_  (
    .CK(clk),
    .D(_00195_),
    .Q(reg_next_pc[11]),
    .QN(_28933_)
  );
  DFF_X1 reg_next_pc_reg_12_  (
    .CK(clk),
    .D(_00196_),
    .Q(reg_next_pc[12]),
    .QN(_28932_)
  );
  DFF_X1 reg_next_pc_reg_13_  (
    .CK(clk),
    .D(_00197_),
    .Q(reg_next_pc[13]),
    .QN(_28931_)
  );
  DFF_X1 reg_next_pc_reg_14_  (
    .CK(clk),
    .D(_00198_),
    .Q(reg_next_pc[14]),
    .QN(_28930_)
  );
  DFF_X1 reg_next_pc_reg_15_  (
    .CK(clk),
    .D(_00199_),
    .Q(reg_next_pc[15]),
    .QN(_28929_)
  );
  DFF_X1 reg_next_pc_reg_16_  (
    .CK(clk),
    .D(_00200_),
    .Q(reg_next_pc[16]),
    .QN(_28928_)
  );
  DFF_X1 reg_next_pc_reg_17_  (
    .CK(clk),
    .D(_00201_),
    .Q(reg_next_pc[17]),
    .QN(_28927_)
  );
  DFF_X1 reg_next_pc_reg_18_  (
    .CK(clk),
    .D(_00202_),
    .Q(reg_next_pc[18]),
    .QN(_28926_)
  );
  DFF_X1 reg_next_pc_reg_19_  (
    .CK(clk),
    .D(_00203_),
    .Q(reg_next_pc[19]),
    .QN(_28925_)
  );
  DFF_X1 reg_next_pc_reg_1_  (
    .CK(clk),
    .D(_00185_),
    .Q(reg_next_pc[1]),
    .QN(_28943_)
  );
  DFF_X1 reg_next_pc_reg_20_  (
    .CK(clk),
    .D(_00204_),
    .Q(reg_next_pc[20]),
    .QN(_28924_)
  );
  DFF_X1 reg_next_pc_reg_21_  (
    .CK(clk),
    .D(_00205_),
    .Q(reg_next_pc[21]),
    .QN(_28923_)
  );
  DFF_X1 reg_next_pc_reg_22_  (
    .CK(clk),
    .D(_00206_),
    .Q(reg_next_pc[22]),
    .QN(_28922_)
  );
  DFF_X1 reg_next_pc_reg_23_  (
    .CK(clk),
    .D(_00207_),
    .Q(reg_next_pc[23]),
    .QN(_28921_)
  );
  DFF_X1 reg_next_pc_reg_24_  (
    .CK(clk),
    .D(_00208_),
    .Q(reg_next_pc[24]),
    .QN(_28920_)
  );
  DFF_X1 reg_next_pc_reg_25_  (
    .CK(clk),
    .D(_00209_),
    .Q(reg_next_pc[25]),
    .QN(_28919_)
  );
  DFF_X1 reg_next_pc_reg_26_  (
    .CK(clk),
    .D(_00210_),
    .Q(reg_next_pc[26]),
    .QN(_28918_)
  );
  DFF_X1 reg_next_pc_reg_27_  (
    .CK(clk),
    .D(_00211_),
    .Q(reg_next_pc[27]),
    .QN(_28917_)
  );
  DFF_X1 reg_next_pc_reg_28_  (
    .CK(clk),
    .D(_00212_),
    .Q(reg_next_pc[28]),
    .QN(_28916_)
  );
  DFF_X1 reg_next_pc_reg_29_  (
    .CK(clk),
    .D(_00213_),
    .Q(reg_next_pc[29]),
    .QN(_28915_)
  );
  DFF_X1 reg_next_pc_reg_2_  (
    .CK(clk),
    .D(_00186_),
    .Q(reg_next_pc[2]),
    .QN(_28942_)
  );
  DFF_X1 reg_next_pc_reg_30_  (
    .CK(clk),
    .D(_00214_),
    .Q(reg_next_pc[30]),
    .QN(_28914_)
  );
  DFF_X1 reg_next_pc_reg_31_  (
    .CK(clk),
    .D(_00215_),
    .Q(reg_next_pc[31]),
    .QN(_28913_)
  );
  DFF_X1 reg_next_pc_reg_3_  (
    .CK(clk),
    .D(_00187_),
    .Q(reg_next_pc[3]),
    .QN(_28941_)
  );
  DFF_X1 reg_next_pc_reg_4_  (
    .CK(clk),
    .D(_00188_),
    .Q(reg_next_pc[4]),
    .QN(_28940_)
  );
  DFF_X1 reg_next_pc_reg_5_  (
    .CK(clk),
    .D(_00189_),
    .Q(reg_next_pc[5]),
    .QN(_28939_)
  );
  DFF_X1 reg_next_pc_reg_6_  (
    .CK(clk),
    .D(_00190_),
    .Q(reg_next_pc[6]),
    .QN(_28938_)
  );
  DFF_X1 reg_next_pc_reg_7_  (
    .CK(clk),
    .D(_00191_),
    .Q(reg_next_pc[7]),
    .QN(_28937_)
  );
  DFF_X1 reg_next_pc_reg_8_  (
    .CK(clk),
    .D(_00192_),
    .Q(reg_next_pc[8]),
    .QN(_28936_)
  );
  DFF_X1 reg_next_pc_reg_9_  (
    .CK(clk),
    .D(_00193_),
    .Q(reg_next_pc[9]),
    .QN(_28935_)
  );
  DFF_X1 reg_op1_reg_0_  (
    .CK(clk),
    .D(_00058_),
    .Q(reg_op1[0]),
    .QN(_00044_)
  );
  DFF_X1 reg_op1_reg_10_  (
    .CK(clk),
    .D(_00067_),
    .Q(reg_op1[10]),
    .QN(_29059_)
  );
  DFF_X1 reg_op1_reg_11_  (
    .CK(clk),
    .D(_00068_),
    .Q(reg_op1[11]),
    .QN(_29058_)
  );
  DFF_X1 reg_op1_reg_12_  (
    .CK(clk),
    .D(_00069_),
    .Q(reg_op1[12]),
    .QN(_29057_)
  );
  DFF_X1 reg_op1_reg_13_  (
    .CK(clk),
    .D(_00070_),
    .Q(reg_op1[13]),
    .QN(_29056_)
  );
  DFF_X1 reg_op1_reg_14_  (
    .CK(clk),
    .D(_00071_),
    .Q(reg_op1[14]),
    .QN(_29055_)
  );
  DFF_X1 reg_op1_reg_15_  (
    .CK(clk),
    .D(_00072_),
    .Q(reg_op1[15]),
    .QN(_29054_)
  );
  DFF_X1 reg_op1_reg_16_  (
    .CK(clk),
    .D(_00073_),
    .Q(reg_op1[16]),
    .QN(_29053_)
  );
  DFF_X1 reg_op1_reg_17_  (
    .CK(clk),
    .D(_00074_),
    .Q(reg_op1[17]),
    .QN(_29052_)
  );
  DFF_X1 reg_op1_reg_18_  (
    .CK(clk),
    .D(_00075_),
    .Q(reg_op1[18]),
    .QN(_29051_)
  );
  DFF_X1 reg_op1_reg_19_  (
    .CK(clk),
    .D(_00076_),
    .Q(reg_op1[19]),
    .QN(_29050_)
  );
  DFF_X1 reg_op1_reg_1_  (
    .CK(clk),
    .D(_01575_),
    .Q(reg_op1[1]),
    .QN(_29146_[1])
  );
  DFF_X1 reg_op1_reg_20_  (
    .CK(clk),
    .D(_00077_),
    .Q(reg_op1[20]),
    .QN(_29049_)
  );
  DFF_X1 reg_op1_reg_21_  (
    .CK(clk),
    .D(_00078_),
    .Q(reg_op1[21]),
    .QN(_29048_)
  );
  DFF_X1 reg_op1_reg_22_  (
    .CK(clk),
    .D(_00079_),
    .Q(reg_op1[22]),
    .QN(_29047_)
  );
  DFF_X1 reg_op1_reg_23_  (
    .CK(clk),
    .D(_00080_),
    .Q(reg_op1[23]),
    .QN(_29046_)
  );
  DFF_X1 reg_op1_reg_24_  (
    .CK(clk),
    .D(_00081_),
    .Q(reg_op1[24]),
    .QN(_29045_)
  );
  DFF_X1 reg_op1_reg_25_  (
    .CK(clk),
    .D(_00082_),
    .Q(reg_op1[25]),
    .QN(_29044_)
  );
  DFF_X1 reg_op1_reg_26_  (
    .CK(clk),
    .D(_00083_),
    .Q(reg_op1[26]),
    .QN(_29043_)
  );
  DFF_X1 reg_op1_reg_27_  (
    .CK(clk),
    .D(_00084_),
    .Q(reg_op1[27]),
    .QN(_29042_)
  );
  DFF_X1 reg_op1_reg_28_  (
    .CK(clk),
    .D(_00085_),
    .Q(reg_op1[28]),
    .QN(_29041_)
  );
  DFF_X1 reg_op1_reg_29_  (
    .CK(clk),
    .D(_00086_),
    .Q(reg_op1[29]),
    .QN(_29040_)
  );
  DFF_X1 reg_op1_reg_2_  (
    .CK(clk),
    .D(_00059_),
    .Q(reg_op1[2]),
    .QN(_29067_)
  );
  DFF_X1 reg_op1_reg_30_  (
    .CK(clk),
    .D(_00087_),
    .Q(reg_op1[30]),
    .QN(_29068_)
  );
  DFF_X1 reg_op1_reg_31_  (
    .CK(clk),
    .D(_00280_),
    .Q(reg_op1[31]),
    .QN(_29078_)
  );
  DFF_X1 reg_op1_reg_3_  (
    .CK(clk),
    .D(_00060_),
    .Q(reg_op1[3]),
    .QN(_29066_)
  );
  DFF_X1 reg_op1_reg_4_  (
    .CK(clk),
    .D(_00061_),
    .Q(reg_op1[4]),
    .QN(_29065_)
  );
  DFF_X1 reg_op1_reg_5_  (
    .CK(clk),
    .D(_00062_),
    .Q(reg_op1[5]),
    .QN(_29064_)
  );
  DFF_X1 reg_op1_reg_6_  (
    .CK(clk),
    .D(_00063_),
    .Q(reg_op1[6]),
    .QN(_29063_)
  );
  DFF_X1 reg_op1_reg_7_  (
    .CK(clk),
    .D(_00064_),
    .Q(reg_op1[7]),
    .QN(_29062_)
  );
  DFF_X1 reg_op1_reg_8_  (
    .CK(clk),
    .D(_00065_),
    .Q(reg_op1[8]),
    .QN(_29061_)
  );
  DFF_X1 reg_op1_reg_9_  (
    .CK(clk),
    .D(_00066_),
    .Q(reg_op1[9]),
    .QN(_29060_)
  );
  DFF_X1 reg_op2_reg_0_  (
    .CK(clk),
    .D(_00281_),
    .Q(reg_op2[0]),
    .QN(_29151_[0])
  );
  DFF_X1 reg_op2_reg_10_  (
    .CK(clk),
    .D(_00291_),
    .Q(reg_op2[10]),
    .QN(_29151_[10])
  );
  DFF_X1 reg_op2_reg_11_  (
    .CK(clk),
    .D(_00292_),
    .Q(reg_op2[11]),
    .QN(_29151_[11])
  );
  DFF_X1 reg_op2_reg_12_  (
    .CK(clk),
    .D(_00293_),
    .Q(reg_op2[12]),
    .QN(_29151_[12])
  );
  DFF_X1 reg_op2_reg_13_  (
    .CK(clk),
    .D(_00294_),
    .Q(reg_op2[13]),
    .QN(_29151_[13])
  );
  DFF_X1 reg_op2_reg_14_  (
    .CK(clk),
    .D(_00295_),
    .Q(reg_op2[14]),
    .QN(_29151_[14])
  );
  DFF_X1 reg_op2_reg_15_  (
    .CK(clk),
    .D(_00296_),
    .Q(reg_op2[15]),
    .QN(_29151_[15])
  );
  DFF_X1 reg_op2_reg_16_  (
    .CK(clk),
    .D(_00297_),
    .Q(reg_op2[16]),
    .QN(_29151_[16])
  );
  DFF_X1 reg_op2_reg_17_  (
    .CK(clk),
    .D(_00298_),
    .Q(reg_op2[17]),
    .QN(_29151_[17])
  );
  DFF_X1 reg_op2_reg_18_  (
    .CK(clk),
    .D(_00299_),
    .Q(reg_op2[18]),
    .QN(_29151_[18])
  );
  DFF_X1 reg_op2_reg_19_  (
    .CK(clk),
    .D(_00300_),
    .Q(reg_op2[19]),
    .QN(_29151_[19])
  );
  DFF_X1 reg_op2_reg_1_  (
    .CK(clk),
    .D(_00282_),
    .Q(reg_op2[1]),
    .QN(_29151_[1])
  );
  DFF_X1 reg_op2_reg_20_  (
    .CK(clk),
    .D(_00301_),
    .Q(reg_op2[20]),
    .QN(_29151_[20])
  );
  DFF_X1 reg_op2_reg_21_  (
    .CK(clk),
    .D(_00302_),
    .Q(reg_op2[21]),
    .QN(_29151_[21])
  );
  DFF_X1 reg_op2_reg_22_  (
    .CK(clk),
    .D(_00303_),
    .Q(reg_op2[22]),
    .QN(_29151_[22])
  );
  DFF_X1 reg_op2_reg_23_  (
    .CK(clk),
    .D(_00304_),
    .Q(reg_op2[23]),
    .QN(_29151_[23])
  );
  DFF_X1 reg_op2_reg_24_  (
    .CK(clk),
    .D(_00305_),
    .Q(reg_op2[24]),
    .QN(_29151_[24])
  );
  DFF_X1 reg_op2_reg_25_  (
    .CK(clk),
    .D(_00306_),
    .Q(reg_op2[25]),
    .QN(_29151_[25])
  );
  DFF_X1 reg_op2_reg_26_  (
    .CK(clk),
    .D(_00307_),
    .Q(reg_op2[26]),
    .QN(_29151_[26])
  );
  DFF_X1 reg_op2_reg_27_  (
    .CK(clk),
    .D(_00308_),
    .Q(reg_op2[27]),
    .QN(_29151_[27])
  );
  DFF_X1 reg_op2_reg_28_  (
    .CK(clk),
    .D(_00309_),
    .Q(reg_op2[28]),
    .QN(_29151_[28])
  );
  DFF_X1 reg_op2_reg_29_  (
    .CK(clk),
    .D(_00310_),
    .Q(reg_op2[29]),
    .QN(_29151_[29])
  );
  DFF_X1 reg_op2_reg_2_  (
    .CK(clk),
    .D(_00283_),
    .Q(reg_op2[2]),
    .QN(_29151_[2])
  );
  DFF_X1 reg_op2_reg_30_  (
    .CK(clk),
    .D(_00311_),
    .Q(reg_op2[30]),
    .QN(_29151_[30])
  );
  DFF_X1 reg_op2_reg_31_  (
    .CK(clk),
    .D(_00312_),
    .Q(reg_op2[31]),
    .QN(_29151_[31])
  );
  DFF_X1 reg_op2_reg_3_  (
    .CK(clk),
    .D(_00284_),
    .Q(reg_op2[3]),
    .QN(_29151_[3])
  );
  DFF_X1 reg_op2_reg_4_  (
    .CK(clk),
    .D(_00285_),
    .Q(reg_op2[4]),
    .QN(_29151_[4])
  );
  DFF_X1 reg_op2_reg_5_  (
    .CK(clk),
    .D(_00286_),
    .Q(reg_op2[5]),
    .QN(_29151_[5])
  );
  DFF_X1 reg_op2_reg_6_  (
    .CK(clk),
    .D(_00287_),
    .Q(reg_op2[6]),
    .QN(_29151_[6])
  );
  DFF_X1 reg_op2_reg_7_  (
    .CK(clk),
    .D(_00288_),
    .Q(reg_op2[7]),
    .QN(_29151_[7])
  );
  DFF_X1 reg_op2_reg_8_  (
    .CK(clk),
    .D(_00289_),
    .Q(reg_op2[8]),
    .QN(_29151_[8])
  );
  DFF_X1 reg_op2_reg_9_  (
    .CK(clk),
    .D(_00290_),
    .Q(reg_op2[9]),
    .QN(_29151_[9])
  );
  DFF_X1 reg_out_reg_0_  (
    .CK(clk),
    .D(_00005_[0]),
    .Q(reg_out[0]),
    .QN(_29079_)
  );
  DFF_X1 reg_out_reg_10_  (
    .CK(clk),
    .D(_00005_[10]),
    .Q(reg_out[10]),
    .QN(_29089_)
  );
  DFF_X1 reg_out_reg_11_  (
    .CK(clk),
    .D(_00005_[11]),
    .Q(reg_out[11]),
    .QN(_29090_)
  );
  DFF_X1 reg_out_reg_12_  (
    .CK(clk),
    .D(_00005_[12]),
    .Q(reg_out[12]),
    .QN(_29091_)
  );
  DFF_X1 reg_out_reg_13_  (
    .CK(clk),
    .D(_00005_[13]),
    .Q(reg_out[13]),
    .QN(_29092_)
  );
  DFF_X1 reg_out_reg_14_  (
    .CK(clk),
    .D(_00005_[14]),
    .Q(reg_out[14]),
    .QN(_29093_)
  );
  DFF_X1 reg_out_reg_15_  (
    .CK(clk),
    .D(_00005_[15]),
    .Q(reg_out[15]),
    .QN(_29094_)
  );
  DFF_X1 reg_out_reg_16_  (
    .CK(clk),
    .D(_00005_[16]),
    .Q(reg_out[16]),
    .QN(_29095_)
  );
  DFF_X1 reg_out_reg_17_  (
    .CK(clk),
    .D(_00005_[17]),
    .Q(reg_out[17]),
    .QN(_29096_)
  );
  DFF_X1 reg_out_reg_18_  (
    .CK(clk),
    .D(_00005_[18]),
    .Q(reg_out[18]),
    .QN(_29097_)
  );
  DFF_X1 reg_out_reg_19_  (
    .CK(clk),
    .D(_00005_[19]),
    .Q(reg_out[19]),
    .QN(_29098_)
  );
  DFF_X1 reg_out_reg_1_  (
    .CK(clk),
    .D(_00005_[1]),
    .Q(reg_out[1]),
    .QN(_29080_)
  );
  DFF_X1 reg_out_reg_20_  (
    .CK(clk),
    .D(_00005_[20]),
    .Q(reg_out[20]),
    .QN(_29099_)
  );
  DFF_X1 reg_out_reg_21_  (
    .CK(clk),
    .D(_00005_[21]),
    .Q(reg_out[21]),
    .QN(_29100_)
  );
  DFF_X1 reg_out_reg_22_  (
    .CK(clk),
    .D(_00005_[22]),
    .Q(reg_out[22]),
    .QN(_29101_)
  );
  DFF_X1 reg_out_reg_23_  (
    .CK(clk),
    .D(_00005_[23]),
    .Q(reg_out[23]),
    .QN(_29102_)
  );
  DFF_X1 reg_out_reg_24_  (
    .CK(clk),
    .D(_00005_[24]),
    .Q(reg_out[24]),
    .QN(_29103_)
  );
  DFF_X1 reg_out_reg_25_  (
    .CK(clk),
    .D(_00005_[25]),
    .Q(reg_out[25]),
    .QN(_29104_)
  );
  DFF_X1 reg_out_reg_26_  (
    .CK(clk),
    .D(_00005_[26]),
    .Q(reg_out[26]),
    .QN(_29105_)
  );
  DFF_X1 reg_out_reg_27_  (
    .CK(clk),
    .D(_00005_[27]),
    .Q(reg_out[27]),
    .QN(_29106_)
  );
  DFF_X1 reg_out_reg_28_  (
    .CK(clk),
    .D(_00005_[28]),
    .Q(reg_out[28]),
    .QN(_29107_)
  );
  DFF_X1 reg_out_reg_29_  (
    .CK(clk),
    .D(_00005_[29]),
    .Q(reg_out[29]),
    .QN(_29108_)
  );
  DFF_X1 reg_out_reg_2_  (
    .CK(clk),
    .D(_00005_[2]),
    .Q(reg_out[2]),
    .QN(_29081_)
  );
  DFF_X1 reg_out_reg_30_  (
    .CK(clk),
    .D(_00005_[30]),
    .Q(reg_out[30]),
    .QN(_29109_)
  );
  DFF_X1 reg_out_reg_31_  (
    .CK(clk),
    .D(_00005_[31]),
    .Q(reg_out[31]),
    .QN(_29110_)
  );
  DFF_X1 reg_out_reg_3_  (
    .CK(clk),
    .D(_00005_[3]),
    .Q(reg_out[3]),
    .QN(_29082_)
  );
  DFF_X1 reg_out_reg_4_  (
    .CK(clk),
    .D(_00005_[4]),
    .Q(reg_out[4]),
    .QN(_29083_)
  );
  DFF_X1 reg_out_reg_5_  (
    .CK(clk),
    .D(_00005_[5]),
    .Q(reg_out[5]),
    .QN(_29084_)
  );
  DFF_X1 reg_out_reg_6_  (
    .CK(clk),
    .D(_00005_[6]),
    .Q(reg_out[6]),
    .QN(_29085_)
  );
  DFF_X1 reg_out_reg_7_  (
    .CK(clk),
    .D(_00005_[7]),
    .Q(reg_out[7]),
    .QN(_29086_)
  );
  DFF_X1 reg_out_reg_8_  (
    .CK(clk),
    .D(_00005_[8]),
    .Q(reg_out[8]),
    .QN(_29087_)
  );
  DFF_X1 reg_out_reg_9_  (
    .CK(clk),
    .D(_00005_[9]),
    .Q(reg_out[9]),
    .QN(_29088_)
  );
  DFF_X1 reg_pc_reg_10_  (
    .CK(clk),
    .D(_00163_),
    .Q(reg_pc[10]),
    .QN(_28965_)
  );
  DFF_X1 reg_pc_reg_11_  (
    .CK(clk),
    .D(_00164_),
    .Q(reg_pc[11]),
    .QN(_28964_)
  );
  DFF_X1 reg_pc_reg_12_  (
    .CK(clk),
    .D(_00165_),
    .Q(reg_pc[12]),
    .QN(_28963_)
  );
  DFF_X1 reg_pc_reg_13_  (
    .CK(clk),
    .D(_00166_),
    .Q(reg_pc[13]),
    .QN(_28962_)
  );
  DFF_X1 reg_pc_reg_14_  (
    .CK(clk),
    .D(_00167_),
    .Q(reg_pc[14]),
    .QN(_28961_)
  );
  DFF_X1 reg_pc_reg_15_  (
    .CK(clk),
    .D(_00168_),
    .Q(reg_pc[15]),
    .QN(_28960_)
  );
  DFF_X1 reg_pc_reg_16_  (
    .CK(clk),
    .D(_00169_),
    .Q(reg_pc[16]),
    .QN(_28959_)
  );
  DFF_X1 reg_pc_reg_17_  (
    .CK(clk),
    .D(_00170_),
    .Q(reg_pc[17]),
    .QN(_28958_)
  );
  DFF_X1 reg_pc_reg_18_  (
    .CK(clk),
    .D(_00171_),
    .Q(reg_pc[18]),
    .QN(_28957_)
  );
  DFF_X1 reg_pc_reg_19_  (
    .CK(clk),
    .D(_00172_),
    .Q(reg_pc[19]),
    .QN(_28956_)
  );
  DFF_X1 reg_pc_reg_1_  (
    .CK(clk),
    .D(_00154_),
    .Q(reg_pc[1]),
    .QN(_28973_)
  );
  DFF_X1 reg_pc_reg_20_  (
    .CK(clk),
    .D(_00173_),
    .Q(reg_pc[20]),
    .QN(_28955_)
  );
  DFF_X1 reg_pc_reg_21_  (
    .CK(clk),
    .D(_00174_),
    .Q(reg_pc[21]),
    .QN(_28954_)
  );
  DFF_X1 reg_pc_reg_22_  (
    .CK(clk),
    .D(_00175_),
    .Q(reg_pc[22]),
    .QN(_28953_)
  );
  DFF_X1 reg_pc_reg_23_  (
    .CK(clk),
    .D(_00176_),
    .Q(reg_pc[23]),
    .QN(_28952_)
  );
  DFF_X1 reg_pc_reg_24_  (
    .CK(clk),
    .D(_00177_),
    .Q(reg_pc[24]),
    .QN(_28951_)
  );
  DFF_X1 reg_pc_reg_25_  (
    .CK(clk),
    .D(_00178_),
    .Q(reg_pc[25]),
    .QN(_28950_)
  );
  DFF_X1 reg_pc_reg_26_  (
    .CK(clk),
    .D(_00179_),
    .Q(reg_pc[26]),
    .QN(_28949_)
  );
  DFF_X1 reg_pc_reg_27_  (
    .CK(clk),
    .D(_00180_),
    .Q(reg_pc[27]),
    .QN(_28948_)
  );
  DFF_X1 reg_pc_reg_28_  (
    .CK(clk),
    .D(_00181_),
    .Q(reg_pc[28]),
    .QN(_28947_)
  );
  DFF_X1 reg_pc_reg_29_  (
    .CK(clk),
    .D(_00182_),
    .Q(reg_pc[29]),
    .QN(_28946_)
  );
  DFF_X1 reg_pc_reg_2_  (
    .CK(clk),
    .D(_00155_),
    .Q(reg_pc[2]),
    .QN(_29145_[98])
  );
  DFF_X1 reg_pc_reg_30_  (
    .CK(clk),
    .D(_00183_),
    .Q(reg_pc[30]),
    .QN(_28945_)
  );
  DFF_X1 reg_pc_reg_31_  (
    .CK(clk),
    .D(_00184_),
    .Q(reg_pc[31]),
    .QN(_28944_)
  );
  DFF_X1 reg_pc_reg_3_  (
    .CK(clk),
    .D(_00156_),
    .Q(reg_pc[3]),
    .QN(_28972_)
  );
  DFF_X1 reg_pc_reg_4_  (
    .CK(clk),
    .D(_00157_),
    .Q(reg_pc[4]),
    .QN(_28971_)
  );
  DFF_X1 reg_pc_reg_5_  (
    .CK(clk),
    .D(_00158_),
    .Q(reg_pc[5]),
    .QN(_28970_)
  );
  DFF_X1 reg_pc_reg_6_  (
    .CK(clk),
    .D(_00159_),
    .Q(reg_pc[6]),
    .QN(_28969_)
  );
  DFF_X1 reg_pc_reg_7_  (
    .CK(clk),
    .D(_00160_),
    .Q(reg_pc[7]),
    .QN(_28968_)
  );
  DFF_X1 reg_pc_reg_8_  (
    .CK(clk),
    .D(_00161_),
    .Q(reg_pc[8]),
    .QN(_28967_)
  );
  DFF_X1 reg_pc_reg_9_  (
    .CK(clk),
    .D(_00162_),
    .Q(reg_pc[9]),
    .QN(_28966_)
  );
  DFF_X1 reg_sh_reg_0_  (
    .CK(clk),
    .D(_00006_[0]),
    .Q(reg_sh[0]),
    .QN(_29149_[0])
  );
  DFF_X1 reg_sh_reg_1_  (
    .CK(clk),
    .D(_00006_[1]),
    .Q(reg_sh[1]),
    .QN(_29149_[1])
  );
  DFF_X1 reg_sh_reg_2_  (
    .CK(clk),
    .D(_00006_[2]),
    .Q(reg_sh[2]),
    .QN(_29150_[2])
  );
  DFF_X1 reg_sh_reg_3_  (
    .CK(clk),
    .D(_00006_[3]),
    .Q(reg_sh[3]),
    .QN(_29149_[3])
  );
  DFF_X1 reg_sh_reg_4_  (
    .CK(clk),
    .D(_00006_[4]),
    .Q(reg_sh[4]),
    .QN(_29149_[4])
  );
  DFF_X1 trap_reg  (
    .CK(clk),
    .D(_00370_),
    .Q(trap),
    .QN(_28808_)
  );
  assign { _29145_[97:96], _29145_[63:0] } = { reg_pc[1], reg_next_pc[0], reg_next_pc, 1'b1 };
  assign _29146_[0] = reg_op1[1];
  assign _29147_[63:1] = count_cycle[63:1];
  assign _29148_[63:1] = count_instr[63:1];
  assign { _29149_[31:5], _29149_[2] } = { 1'b1, reg_sh[2] };
  assign { _29150_[30:5], _29150_[1:0] } = { _29150_[31], _29150_[31], _29150_[31], _29150_[31], _29150_[31], _29150_[31], _29150_[31], _29150_[31], _29150_[31], _29150_[31], _29150_[31], _29150_[31], _29150_[31], _29150_[31], _29150_[31], _29150_[31], _29150_[31], _29150_[31], _29150_[31], _29150_[31], _29150_[31], _29150_[31], _29150_[31], _29150_[31], _29150_[31], _29150_[31], reg_sh[1:0] };
  assign compressed_instr = 1'b1;
  assign current_pc = 1'b1;
  assign dbg_mem_addr = { mem_addr[31:2], 1'b1 };
  assign dbg_mem_instr = mem_instr;
  assign dbg_mem_rdata = mem_rdata;
  assign dbg_mem_ready = mem_ready;
  assign dbg_mem_valid = mem_valid;
  assign dbg_mem_wdata = mem_wdata;
  assign dbg_mem_wstrb = mem_wstrb;
  assign { decoded_imm_j[31], decoded_imm_j[29:20], decoded_imm_j[17:15], decoded_imm_j[11], decoded_imm_j[3:0] } = { decoded_imm_j[30], decoded_imm_j[30], decoded_imm_j[30], decoded_imm_j[30], decoded_imm_j[30], decoded_imm_j[30], decoded_imm_j[30], decoded_imm_j[30], decoded_imm_j[30], decoded_imm_j[30], decoded_imm_j[30], decoded_rs1[2:0], decoded_rs2[0], decoded_rs2[3:1], 1'b1 };
  assign decoded_rs = 1'b1;
  assign decoded_rs1[4:3] = decoded_imm_j[19:18];
  assign decoded_rs2[4] = decoded_imm_j[4];
  assign do_waitirq = 1'b1;
  assign { eoi[31], eoi[29:0] } = { eoi[30], eoi[30], eoi[30], eoi[30], eoi[30], eoi[30], eoi[30], eoi[30], eoi[30], eoi[30], eoi[30], eoi[30], eoi[30], eoi[30], eoi[30], eoi[30], eoi[30], eoi[30], eoi[30], eoi[30], eoi[30], eoi[30], eoi[30], eoi[30], eoi[30], eoi[30], eoi[30], eoi[30], eoi[30], eoi[30], eoi[30] };
  assign instr_getq = 1'b1;
  assign instr_maskirq = 1'b1;
  assign instr_retirq = 1'b1;
  assign instr_setq = 1'b1;
  assign instr_timer = 1'b1;
  assign instr_waitirq = 1'b1;
  assign irq_mask = 32'd4294967295;
  assign { irq_pending[31:3], irq_pending[0] } = 1'b1;
  assign latched_compr = 1'b1;
  assign mem_addr[1:0] = 1'b1;
  assign mem_la_addr[1:0] = 1'b1;
  assign mem_la_firstword = 1'b1;
  assign mem_la_firstword_reg = 1'b1;
  assign mem_la_firstword_xfer = 1'b1;
  assign mem_la_secondword = 1'b1;
  assign mem_la_use_prefetched_high_word = 1'b1;
  assign next_irq_pending = { 1'b1, irq_pending[2:1], 1'b1 };
  assign pcpi_div_rd = 1'b1;
  assign pcpi_div_ready = 1'b1;
  assign pcpi_div_wait = 1'b1;
  assign pcpi_div_wr = 1'b1;
  assign pcpi_insn = 1'b1;
  assign pcpi_int_rd = 1'b1;
  assign pcpi_int_ready = 1'b1;
  assign pcpi_int_wait = 1'b1;
  assign pcpi_int_wr = 1'b1;
  assign pcpi_mul_rd = 1'b1;
  assign pcpi_mul_ready = 1'b1;
  assign pcpi_mul_wait = 1'b1;
  assign pcpi_mul_wr = 1'b1;
  assign pcpi_rs1 = reg_op1;
  assign pcpi_rs2 = reg_op2;
  assign pcpi_timeout = 1'b1;
  assign pcpi_valid = 1'b1;
  assign reg_pc[0] = reg_next_pc[0];
  assign timer = 32'd0;
  assign trace_data = 1'b1;
  assign trace_valid = 1'b1;
endmodule
